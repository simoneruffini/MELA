
module CU ( CLK, RST_AN, INSTR, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .CTRL_WORD({
        \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] , 
        \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] , 
        \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] , 
        \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] , 
        \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }) );
  input [31:0] INSTR;
  input CLK, RST_AN, \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] ;
  wire   INSTR_31, INSTR_30, INSTR_29, INSTR_28, INSTR_27, INSTR_26,
         \execute_sig_d1[R_TYPE_SEL] , \execute_sig_d1[IMM_SEL] ,
         \execute_sig_d1[PC_PLS_4_SEL] , \execute_sig_d1[ALU_FUNC][3] ,
         \execute_sig_d1[ALU_FUNC][2] , \execute_sig_d1[ALU_FUNC][1] ,
         \execute_sig_d1[ALU_FUNC][0] , \memory_sig_d1[DMEM_WEN] ,
         \memory_sig_d1[BRANCH_EN] , \memory_sig_d1[JUMP_EN] ,
         \memory_sig_d1[COMP_0_INVERT] ,
         \writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d1[JAL_EN] ,
         \writeback_sig_d1[RF_WEN] , \memory_sig_d2[DMEM_WEN] ,
         \memory_sig_d2[BRANCH_EN] , \memory_sig_d2[JUMP_EN] ,
         \memory_sig_d2[COMP_0_INVERT] ,
         \writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d2[JAL_EN] ,
         \writeback_sig_d2[RF_WEN] , \writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ,
         \writeback_sig_d3[JAL_EN] , \writeback_sig_d3[RF_WEN] , N213, N214,
         N215, N216, N217, N218, N224, N228, N229, N231, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n1, n2, n4, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n20, n21, n22, n23, n24, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n117,
         n118, n119, n120, n121, n122, n123;
  assign INSTR_31 = INSTR[31];
  assign INSTR_30 = INSTR[30];
  assign INSTR_29 = INSTR[29];
  assign INSTR_28 = INSTR[28];
  assign INSTR_27 = INSTR[27];
  assign INSTR_26 = INSTR[26];

  DFFR_X1 \decode_sig_d1_reg[J_TYPE_IMM_SEL]  ( .D(n37), .CK(CLK), .RN(n29), 
        .Q(\CTRL_WORD[J_TYPE_IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[IMM_SEL]  ( .D(N218), .CK(CLK), .RN(n29), .Q(
        \execute_sig_d1[IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[PC_PLS_4_SEL]  ( .D(N217), .CK(CLK), .RN(n29), 
        .Q(\execute_sig_d1[PC_PLS_4_SEL] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][3]  ( .D(N216), .CK(CLK), .SN(n32), 
        .Q(\execute_sig_d1[ALU_FUNC][3] ) );
  DFFR_X1 \execute_sig_d1_reg[ALU_FUNC][2]  ( .D(N215), .CK(CLK), .RN(n29), 
        .Q(\execute_sig_d1[ALU_FUNC][2] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][1]  ( .D(N214), .CK(CLK), .SN(n32), 
        .Q(\execute_sig_d1[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][0]  ( .D(N213), .CK(CLK), .SN(n32), 
        .Q(\execute_sig_d1[ALU_FUNC][0] ) );
  DFFR_X1 \memory_sig_d1_reg[BRANCH_EN]  ( .D(n38), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d1[BRANCH_EN] ) );
  DFFR_X1 \memory_sig_d1_reg[JUMP_EN]  ( .D(n37), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d1[JUMP_EN] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n35), .CK(CLK), 
        .RN(n29), .Q(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WEN]  ( .D(N224), .CK(CLK), .RN(n29), .Q(
        \writeback_sig_d1[RF_WEN] ) );
  SDFFR_X1 \execute_sig_d2_reg[PC_PLS_4_SEL]  ( .D(1'b0), .SI(n34), .SE(
        \execute_sig_d1[PC_PLS_4_SEL] ), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[PC_PLS_4_SEL] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][3]  ( .D(N231), .CK(CLK), .SN(n31), 
        .Q(\CTRL_WORD[ALU_FUNC][3] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][1]  ( .D(N229), .CK(CLK), .SN(n32), 
        .Q(\CTRL_WORD[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][0]  ( .D(N228), .CK(CLK), .SN(n31), 
        .Q(\CTRL_WORD[ALU_FUNC][0] ) );
  SDFFR_X1 \writeback_sig_d4_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(1'b0), .SI(n41), 
        .SE(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ) );
  NAND3_X1 U118 ( .A1(n68), .A2(n40), .A3(INSTR_31), .ZN(n54) );
  NAND3_X1 U119 ( .A1(INSTR_29), .A2(n53), .A3(n46), .ZN(n71) );
  NAND3_X1 U120 ( .A1(INSTR_26), .A2(n80), .A3(INSTR_29), .ZN(n79) );
  OAI33_X1 U121 ( .A1(n122), .A2(INSTR[5]), .A3(n119), .B1(n123), .B2(INSTR[2]), .B3(n98), .ZN(n97) );
  NAND3_X1 U122 ( .A1(INSTR_26), .A2(n51), .A3(INSTR_27), .ZN(n77) );
  NAND3_X1 U123 ( .A1(INSTR_27), .A2(n45), .A3(INSTR_28), .ZN(n108) );
  NAND3_X1 U124 ( .A1(n96), .A2(n117), .A3(INSTR_30), .ZN(n110) );
  NAND3_X1 U125 ( .A1(n113), .A2(n121), .A3(INSTR[2]), .ZN(n104) );
  NAND3_X1 U126 ( .A1(n113), .A2(n120), .A3(INSTR[3]), .ZN(n98) );
  NAND3_X1 U127 ( .A1(n113), .A2(INSTR[5]), .A3(INSTR[1]), .ZN(n114) );
  NAND3_X1 U128 ( .A1(n39), .A2(INSTR_27), .A3(n116), .ZN(n55) );
  DFFRS_X2 \execute_sig_d2_reg[IMM_SEL]  ( .D(n26), .CK(CLK), .RN(RST_AN), 
        .SN(1'b1), .Q(\CTRL_WORD[IMM_SEL] ) );
  SDFFR_X2 \writeback_sig_d4_reg[JAL_EN]  ( .D(1'b0), .SI(n41), .SE(
        \writeback_sig_d3[JAL_EN] ), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[JAL_EN] ) );
  DFFR_X1 \writeback_sig_d3_reg[RF_WEN]  ( .D(n24), .CK(CLK), .RN(RST_AN), .Q(
        \writeback_sig_d3[RF_WEN] ) );
  DFFR_X1 \writeback_sig_d3_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n23), .CK(CLK), 
        .RN(n31), .Q(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d3_reg[JAL_EN]  ( .D(n22), .CK(CLK), .RN(n31), .Q(
        \writeback_sig_d3[JAL_EN] ) );
  DFFR_X1 \memory_sig_d3_reg[JUMP_EN]  ( .D(n21), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[JUMP_EN] ) );
  DFFR_X1 \memory_sig_d3_reg[DMEM_WEN]  ( .D(n20), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d3_reg[COMP_0_INVERT]  ( .D(n18), .CK(CLK), .RN(n31), 
        .Q(\CTRL_WORD[COMP_0_INVERT] ) );
  DFFR_X1 \memory_sig_d3_reg[BRANCH_EN]  ( .D(n17), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[BRANCH_EN] ) );
  DFFR_X1 \execute_sig_d1_reg[R_TYPE_SEL]  ( .D(n16), .CK(CLK), .RN(n30), .Q(
        \execute_sig_d1[R_TYPE_SEL] ) );
  DFFR_X1 \writeback_sig_d2_reg[RF_WEN]  ( .D(n15), .CK(CLK), .RN(n31), .Q(
        \writeback_sig_d2[RF_WEN] ) );
  DFFR_X1 \writeback_sig_d2_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n14), .CK(CLK), 
        .RN(n30), .Q(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d2_reg[JAL_EN]  ( .D(n13), .CK(CLK), .RN(n31), .Q(
        \writeback_sig_d2[JAL_EN] ) );
  DFFR_X1 \memory_sig_d2_reg[JUMP_EN]  ( .D(n12), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d2[JUMP_EN] ) );
  DFFR_X1 \memory_sig_d2_reg[DMEM_WEN]  ( .D(n11), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d2[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d2_reg[COMP_0_INVERT]  ( .D(n10), .CK(CLK), .RN(n30), 
        .Q(\memory_sig_d2[COMP_0_INVERT] ) );
  DFFR_X1 \memory_sig_d2_reg[BRANCH_EN]  ( .D(n9), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d2[BRANCH_EN] ) );
  DFFR_X1 \execute_sig_d2_reg[R_TYPE_SEL]  ( .D(n8), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[R_TYPE_SEL] ) );
  DFFR_X1 \execute_sig_d2_reg[ALU_FUNC][2]  ( .D(n7), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[ALU_FUNC][2] ) );
  DFFR_X1 \memory_sig_d1_reg[DMEM_WEN]  ( .D(n6), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d1[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d1_reg[COMP_0_INVERT]  ( .D(n4), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d1[COMP_0_INVERT] ) );
  DFFR_X1 \writeback_sig_d1_reg[JAL_EN]  ( .D(n2), .CK(CLK), .RN(n29), .Q(
        \writeback_sig_d1[JAL_EN] ) );
  DFFR_X1 \writeback_sig_d4_reg[RF_WEN]  ( .D(n1), .CK(CLK), .RN(n29), .Q(
        \CTRL_WORD[RF_WEN] ) );
  AND2_X1 U3 ( .A1(\writeback_sig_d3[RF_WEN] ), .A2(n41), .ZN(n1) );
  AND2_X1 U4 ( .A1(INSTR_26), .A2(n37), .ZN(n2) );
  AND2_X1 U6 ( .A1(INSTR_26), .A2(n38), .ZN(n4) );
  AND2_X1 U8 ( .A1(INSTR_29), .A2(n35), .ZN(n6) );
  AND2_X1 U9 ( .A1(\execute_sig_d1[ALU_FUNC][2] ), .A2(n34), .ZN(n7) );
  AND2_X1 U10 ( .A1(\execute_sig_d1[R_TYPE_SEL] ), .A2(n34), .ZN(n8) );
  AND2_X1 U11 ( .A1(\memory_sig_d1[BRANCH_EN] ), .A2(n34), .ZN(n9) );
  AND2_X1 U12 ( .A1(\memory_sig_d1[COMP_0_INVERT] ), .A2(n34), .ZN(n10) );
  AND2_X1 U13 ( .A1(\memory_sig_d1[DMEM_WEN] ), .A2(n34), .ZN(n11) );
  AND2_X1 U14 ( .A1(\memory_sig_d1[JUMP_EN] ), .A2(n34), .ZN(n12) );
  AND2_X1 U15 ( .A1(\writeback_sig_d1[JAL_EN] ), .A2(n34), .ZN(n13) );
  AND2_X1 U16 ( .A1(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ), .A2(n34), .ZN(
        n14) );
  AND2_X1 U17 ( .A1(\writeback_sig_d1[RF_WEN] ), .A2(n34), .ZN(n15) );
  AND2_X1 U18 ( .A1(n43), .A2(n40), .ZN(n16) );
  AND2_X1 U19 ( .A1(\memory_sig_d2[BRANCH_EN] ), .A2(n33), .ZN(n17) );
  AND2_X1 U20 ( .A1(\memory_sig_d2[COMP_0_INVERT] ), .A2(n33), .ZN(n18) );
  AND2_X1 U22 ( .A1(\memory_sig_d2[DMEM_WEN] ), .A2(n33), .ZN(n20) );
  AND2_X1 U23 ( .A1(\memory_sig_d2[JUMP_EN] ), .A2(n33), .ZN(n21) );
  AND2_X1 U24 ( .A1(\writeback_sig_d2[JAL_EN] ), .A2(n33), .ZN(n22) );
  AND2_X1 U25 ( .A1(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ), .A2(n33), .ZN(
        n23) );
  AND2_X1 U26 ( .A1(\writeback_sig_d2[RF_WEN] ), .A2(n33), .ZN(n24) );
  INV_X1 U27 ( .A(n67), .ZN(n39) );
  INV_X1 U28 ( .A(n64), .ZN(n38) );
  INV_X1 U29 ( .A(\HZRD_SIG[FLUSH_FD] ), .ZN(n40) );
  INV_X1 U30 ( .A(\HZRD_SIG[FLUSH_DE] ), .ZN(n34) );
  INV_X1 U31 ( .A(\HZRD_SIG[FLUSH_EM] ), .ZN(n33) );
  AOI21_X1 U32 ( .B1(n56), .B2(n57), .A(\HZRD_SIG[FLUSH_FD] ), .ZN(N224) );
  OAI21_X1 U33 ( .B1(n60), .B2(n61), .A(n42), .ZN(n56) );
  OAI211_X1 U34 ( .C1(n58), .C2(n59), .A(n51), .B(n45), .ZN(n57) );
  OAI22_X1 U35 ( .A1(n51), .A2(n48), .B1(n50), .B2(n62), .ZN(n61) );
  NAND2_X1 U36 ( .A1(n40), .A2(n42), .ZN(n67) );
  NAND4_X1 U37 ( .A1(n49), .A2(n39), .A3(n53), .A4(n45), .ZN(n64) );
  OAI211_X1 U38 ( .C1(n99), .C2(n74), .A(n100), .B(n36), .ZN(N213) );
  OAI211_X1 U39 ( .C1(n106), .C2(n107), .A(n74), .B(n42), .ZN(n100) );
  NOR3_X1 U40 ( .A1(n112), .A2(n81), .A3(n88), .ZN(n99) );
  OAI211_X1 U41 ( .C1(n109), .C2(n53), .A(n110), .B(n95), .ZN(n106) );
  OAI211_X1 U42 ( .C1(n66), .C2(n67), .A(n55), .B(n54), .ZN(N218) );
  AOI21_X1 U43 ( .B1(n52), .B2(n69), .A(n60), .ZN(n66) );
  INV_X1 U44 ( .A(n55), .ZN(n37) );
  INV_X1 U45 ( .A(n101), .ZN(n36) );
  OAI221_X1 U46 ( .B1(n68), .B2(n42), .C1(n102), .C2(n74), .A(n40), .ZN(n101)
         );
  NOR2_X1 U47 ( .A1(n103), .A2(n89), .ZN(n102) );
  NOR3_X1 U48 ( .A1(n104), .A2(n105), .A3(n123), .ZN(n103) );
  NAND2_X1 U49 ( .A1(n64), .A2(n55), .ZN(N217) );
  INV_X1 U50 ( .A(n54), .ZN(n35) );
  BUF_X1 U51 ( .A(n27), .Z(n29) );
  BUF_X1 U52 ( .A(n28), .Z(n31) );
  INV_X1 U53 ( .A(n74), .ZN(n43) );
  BUF_X1 U54 ( .A(n27), .Z(n30) );
  AOI21_X1 U55 ( .B1(n72), .B2(n85), .A(n53), .ZN(n84) );
  INV_X1 U56 ( .A(n96), .ZN(n49) );
  NAND2_X1 U57 ( .A1(n86), .A2(n117), .ZN(n72) );
  INV_X1 U58 ( .A(n69), .ZN(n46) );
  INV_X1 U59 ( .A(n98), .ZN(n118) );
  INV_X1 U60 ( .A(n62), .ZN(n52) );
  INV_X1 U61 ( .A(n87), .ZN(n119) );
  BUF_X1 U62 ( .A(n28), .Z(n32) );
  INV_X1 U63 ( .A(n105), .ZN(n120) );
  INV_X1 U64 ( .A(n63), .ZN(n48) );
  NOR3_X1 U65 ( .A1(INSTR_28), .A2(INSTR_30), .A3(INSTR_29), .ZN(n116) );
  OAI221_X1 U66 ( .B1(n73), .B2(n74), .C1(n43), .C2(n75), .A(n40), .ZN(N216)
         );
  AOI21_X1 U67 ( .B1(INSTR[0]), .B2(n118), .A(n81), .ZN(n73) );
  AOI221_X1 U68 ( .B1(n76), .B2(n50), .C1(INSTR_31), .C2(n77), .A(n78), .ZN(
        n75) );
  OAI221_X1 U69 ( .B1(INSTR_27), .B2(n69), .C1(n49), .C2(n45), .A(n79), .ZN(
        n78) );
  OAI211_X1 U70 ( .C1(n90), .C2(n74), .A(n91), .B(n36), .ZN(N214) );
  AOI21_X1 U71 ( .B1(n87), .B2(n120), .A(n97), .ZN(n90) );
  OAI211_X1 U72 ( .C1(n92), .C2(n47), .A(n74), .B(n42), .ZN(n91) );
  OR2_X1 U73 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][0] ), 
        .ZN(N228) );
  OR2_X1 U74 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][1] ), 
        .ZN(N229) );
  OR2_X1 U75 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][3] ), 
        .ZN(N231) );
  OAI21_X1 U76 ( .B1(n82), .B2(n65), .A(n83), .ZN(N215) );
  AOI211_X1 U77 ( .C1(INSTR[1]), .C2(n87), .A(n88), .B(n89), .ZN(n82) );
  NAND2_X1 U78 ( .A1(n43), .A2(n40), .ZN(n65) );
  OAI211_X1 U79 ( .C1(n84), .C2(n63), .A(n39), .B(INSTR_28), .ZN(n83) );
  NOR4_X1 U80 ( .A1(n122), .A2(n104), .A3(n123), .A4(INSTR[5]), .ZN(n89) );
  NAND4_X1 U81 ( .A1(n53), .A2(n51), .A3(n117), .A4(n111), .ZN(n74) );
  NOR3_X1 U82 ( .A1(INSTR_29), .A2(INSTR_31), .A3(INSTR_30), .ZN(n111) );
  NOR4_X1 U83 ( .A1(INSTR[6]), .A2(INSTR[4]), .A3(INSTR[10]), .A4(n115), .ZN(
        n113) );
  OR3_X1 U84 ( .A1(INSTR[9]), .A2(INSTR[8]), .A3(INSTR[7]), .ZN(n115) );
  NOR4_X1 U85 ( .A1(n114), .A2(INSTR[0]), .A3(INSTR[3]), .A4(INSTR[2]), .ZN(
        n112) );
  NOR3_X1 U86 ( .A1(INSTR[1]), .A2(INSTR[5]), .A3(n119), .ZN(n88) );
  INV_X1 U87 ( .A(INSTR_27), .ZN(n53) );
  INV_X1 U88 ( .A(INSTR[3]), .ZN(n121) );
  AOI211_X1 U89 ( .C1(INSTR_29), .C2(n42), .A(n53), .B(n117), .ZN(n58) );
  NOR2_X1 U90 ( .A1(n104), .A2(INSTR[0]), .ZN(n87) );
  INV_X1 U91 ( .A(INSTR_28), .ZN(n51) );
  NOR2_X1 U92 ( .A1(n50), .A2(INSTR_30), .ZN(n86) );
  OAI22_X1 U93 ( .A1(INSTR_29), .A2(n44), .B1(INSTR_27), .B2(n85), .ZN(n107)
         );
  INV_X1 U94 ( .A(n76), .ZN(n44) );
  OAI211_X1 U95 ( .C1(n45), .C2(n70), .A(n71), .B(n72), .ZN(n60) );
  INV_X1 U96 ( .A(INSTR_31), .ZN(n42) );
  NOR3_X1 U97 ( .A1(INSTR_26), .A2(INSTR_31), .A3(INSTR_27), .ZN(n59) );
  OAI21_X1 U98 ( .B1(INSTR_28), .B2(INSTR_27), .A(n108), .ZN(n76) );
  NOR2_X1 U99 ( .A1(n85), .A2(INSTR_26), .ZN(n63) );
  INV_X1 U100 ( .A(INSTR_29), .ZN(n50) );
  NOR2_X1 U101 ( .A1(n77), .A2(INSTR_30), .ZN(n68) );
  INV_X1 U102 ( .A(INSTR_30), .ZN(n45) );
  AOI21_X1 U103 ( .B1(INSTR_29), .B2(n51), .A(n46), .ZN(n109) );
  OAI211_X1 U104 ( .C1(INSTR_29), .C2(n94), .A(n70), .B(n95), .ZN(n92) );
  AOI21_X1 U105 ( .B1(n53), .B2(n51), .A(n46), .ZN(n94) );
  NAND2_X1 U106 ( .A1(INSTR_30), .A2(n50), .ZN(n85) );
  INV_X1 U107 ( .A(INSTR_26), .ZN(n117) );
  NAND2_X1 U108 ( .A1(INSTR_28), .A2(n53), .ZN(n62) );
  NAND2_X1 U109 ( .A1(INSTR_30), .A2(INSTR_26), .ZN(n69) );
  OAI22_X1 U110 ( .A1(INSTR_31), .A2(INSTR_28), .B1(n53), .B2(n51), .ZN(n80)
         );
  INV_X1 U111 ( .A(INSTR[0]), .ZN(n123) );
  NAND2_X1 U112 ( .A1(n86), .A2(INSTR_26), .ZN(n95) );
  AND3_X1 U113 ( .A1(n118), .A2(n123), .A3(INSTR[2]), .ZN(n81) );
  NAND2_X1 U114 ( .A1(INSTR[5]), .A2(n122), .ZN(n105) );
  NAND2_X1 U115 ( .A1(n49), .A2(INSTR_27), .ZN(n70) );
  INV_X1 U116 ( .A(INSTR[1]), .ZN(n122) );
  NAND2_X1 U117 ( .A1(INSTR_28), .A2(n50), .ZN(n96) );
  INV_X1 U129 ( .A(n93), .ZN(n47) );
  AOI22_X1 U130 ( .A1(n86), .A2(n52), .B1(n62), .B2(INSTR_30), .ZN(n93) );
  BUF_X1 U131 ( .A(RST_AN), .Z(n28) );
  BUF_X1 U132 ( .A(RST_AN), .Z(n27) );
  INV_X1 U133 ( .A(\HZRD_SIG[FLUSH_MWB] ), .ZN(n41) );
  AND2_X1 U135 ( .A1(\execute_sig_d1[IMM_SEL] ), .A2(n34), .ZN(n26) );
endmodule


module REG_PIPO_32_fffffffc_fffffffc ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n19, n20,
         n21;

  DFFS_X1 \reg_mem_reg[31]  ( .D(n96), .CK(CLK), .SN(n21), .Q(DOUT[31]), .QN(
        n64) );
  DFFS_X1 \reg_mem_reg[30]  ( .D(n95), .CK(CLK), .SN(n21), .Q(DOUT[30]) );
  DFFS_X1 \reg_mem_reg[29]  ( .D(n94), .CK(CLK), .SN(n21), .Q(DOUT[29]) );
  DFFS_X1 \reg_mem_reg[28]  ( .D(n93), .CK(CLK), .SN(n21), .Q(DOUT[28]) );
  DFFS_X1 \reg_mem_reg[27]  ( .D(n92), .CK(CLK), .SN(n21), .Q(DOUT[27]) );
  DFFS_X1 \reg_mem_reg[26]  ( .D(n91), .CK(CLK), .SN(n21), .Q(DOUT[26]) );
  DFFS_X1 \reg_mem_reg[25]  ( .D(n90), .CK(CLK), .SN(n20), .Q(DOUT[25]) );
  DFFS_X1 \reg_mem_reg[24]  ( .D(n89), .CK(CLK), .SN(n20), .Q(DOUT[24]) );
  DFFS_X1 \reg_mem_reg[23]  ( .D(n88), .CK(CLK), .SN(n20), .Q(DOUT[23]) );
  DFFS_X1 \reg_mem_reg[22]  ( .D(n87), .CK(CLK), .SN(n20), .Q(DOUT[22]) );
  DFFS_X1 \reg_mem_reg[21]  ( .D(n86), .CK(CLK), .SN(n20), .Q(DOUT[21]) );
  DFFS_X1 \reg_mem_reg[20]  ( .D(n85), .CK(CLK), .SN(n20), .Q(DOUT[20]) );
  DFFS_X1 \reg_mem_reg[19]  ( .D(n84), .CK(CLK), .SN(n20), .Q(DOUT[19]) );
  DFFS_X1 \reg_mem_reg[18]  ( .D(n83), .CK(CLK), .SN(n20), .Q(DOUT[18]) );
  DFFS_X1 \reg_mem_reg[17]  ( .D(n82), .CK(CLK), .SN(n20), .Q(DOUT[17]), .QN(
        n50) );
  DFFS_X1 \reg_mem_reg[16]  ( .D(n81), .CK(CLK), .SN(n20), .Q(DOUT[16]), .QN(
        n49) );
  DFFS_X1 \reg_mem_reg[15]  ( .D(n80), .CK(CLK), .SN(n20), .Q(DOUT[15]), .QN(
        n48) );
  DFFS_X1 \reg_mem_reg[14]  ( .D(n79), .CK(CLK), .SN(n20), .Q(DOUT[14]), .QN(
        n47) );
  DFFS_X1 \reg_mem_reg[13]  ( .D(n78), .CK(CLK), .SN(n20), .Q(DOUT[13]), .QN(
        n46) );
  DFFS_X1 \reg_mem_reg[12]  ( .D(n77), .CK(CLK), .SN(n19), .Q(DOUT[12]), .QN(
        n45) );
  DFFS_X1 \reg_mem_reg[11]  ( .D(n76), .CK(CLK), .SN(n19), .Q(DOUT[11]), .QN(
        n44) );
  DFFS_X1 \reg_mem_reg[10]  ( .D(n75), .CK(CLK), .SN(n19), .Q(DOUT[10]), .QN(
        n43) );
  DFFS_X1 \reg_mem_reg[9]  ( .D(n74), .CK(CLK), .SN(n19), .Q(DOUT[9]), .QN(n42) );
  DFFS_X1 \reg_mem_reg[8]  ( .D(n73), .CK(CLK), .SN(n19), .Q(DOUT[8]), .QN(n41) );
  DFFS_X1 \reg_mem_reg[7]  ( .D(n72), .CK(CLK), .SN(n19), .Q(DOUT[7]), .QN(n40) );
  DFFS_X1 \reg_mem_reg[6]  ( .D(n71), .CK(CLK), .SN(n19), .Q(DOUT[6]), .QN(n39) );
  DFFS_X1 \reg_mem_reg[5]  ( .D(n70), .CK(CLK), .SN(n19), .Q(DOUT[5]), .QN(n38) );
  DFFS_X1 \reg_mem_reg[4]  ( .D(n69), .CK(CLK), .SN(n19), .Q(DOUT[4]), .QN(n37) );
  DFFS_X1 \reg_mem_reg[3]  ( .D(n68), .CK(CLK), .SN(n19), .Q(DOUT[3]), .QN(n36) );
  DFFS_X1 \reg_mem_reg[2]  ( .D(n67), .CK(CLK), .SN(n19), .Q(DOUT[2]), .QN(n35) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n66), .CK(CLK), .RN(n19), .Q(DOUT[1]), .QN(n34) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n65), .CK(CLK), .RN(n19), .Q(DOUT[0]), .QN(n33) );
  BUF_X1 U2 ( .A(RST_AN), .Z(n19) );
  BUF_X1 U3 ( .A(RST_AN), .Z(n20) );
  BUF_X1 U4 ( .A(RST_AN), .Z(n21) );
  OAI21_X1 U5 ( .B1(n47), .B2(EN), .A(n15), .ZN(n79) );
  NAND2_X1 U6 ( .A1(DIN[14]), .A2(EN), .ZN(n15) );
  OAI21_X1 U7 ( .B1(n48), .B2(EN), .A(n16), .ZN(n80) );
  NAND2_X1 U8 ( .A1(DIN[15]), .A2(EN), .ZN(n16) );
  OAI21_X1 U9 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U11 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U13 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U15 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X1 U17 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  OAI21_X1 U19 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  OAI21_X1 U21 ( .B1(n41), .B2(EN), .A(n9), .ZN(n73) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n9) );
  OAI21_X1 U23 ( .B1(n42), .B2(EN), .A(n10), .ZN(n74) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n10) );
  OAI21_X1 U25 ( .B1(n43), .B2(EN), .A(n11), .ZN(n75) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n11) );
  OAI21_X1 U27 ( .B1(n44), .B2(EN), .A(n12), .ZN(n76) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n12) );
  OAI21_X1 U29 ( .B1(n45), .B2(EN), .A(n13), .ZN(n77) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n13) );
  OAI21_X1 U31 ( .B1(n46), .B2(EN), .A(n14), .ZN(n78) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n14) );
  OAI21_X1 U33 ( .B1(n49), .B2(EN), .A(n17), .ZN(n81) );
  NAND2_X1 U34 ( .A1(DIN[16]), .A2(EN), .ZN(n17) );
  OAI21_X1 U35 ( .B1(n50), .B2(EN), .A(n18), .ZN(n82) );
  NAND2_X1 U36 ( .A1(DIN[17]), .A2(EN), .ZN(n18) );
  OAI21_X1 U37 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X1 U38 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U39 ( .B1(n64), .B2(EN), .A(n32), .ZN(n96) );
  NAND2_X1 U40 ( .A1(DIN[31]), .A2(EN), .ZN(n32) );
  OAI21_X1 U41 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X1 U42 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  MUX2_X1 U43 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n83) );
  MUX2_X1 U44 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n84) );
  MUX2_X1 U45 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n85) );
  MUX2_X1 U46 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n86) );
  MUX2_X1 U47 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n87) );
  MUX2_X1 U48 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n88) );
  MUX2_X1 U49 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n89) );
  MUX2_X1 U50 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n90) );
  MUX2_X1 U51 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n91) );
  MUX2_X1 U52 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n92) );
  MUX2_X1 U53 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n93) );
  MUX2_X1 U54 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n94) );
  MUX2_X1 U55 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n95) );
endmodule


module REG_PIPO_32_00000000_00000000_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n99,
         n100, n101, n102;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n98), .CK(CLK), .RN(n4), .Q(DOUT[31]), .QN(
        n66) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n97), .CK(CLK), .RN(n4), .Q(DOUT[30]), .QN(
        n65) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n96), .CK(CLK), .RN(n4), .Q(DOUT[29]), .QN(
        n64) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n95), .CK(CLK), .RN(n4), .Q(DOUT[28]), .QN(
        n63) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n94), .CK(CLK), .RN(n4), .Q(DOUT[27]), .QN(
        n62) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n93), .CK(CLK), .RN(n4), .Q(DOUT[26]), .QN(
        n61) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n92), .CK(CLK), .RN(n4), .Q(DOUT[25]), .QN(
        n60) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n91), .CK(CLK), .RN(n4), .Q(DOUT[24]), .QN(
        n59) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n90), .CK(CLK), .RN(n4), .Q(DOUT[23]), .QN(
        n58) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n89), .CK(CLK), .RN(n4), .Q(DOUT[22]), .QN(
        n57) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n88), .CK(CLK), .RN(n3), .Q(DOUT[21]), .QN(
        n56) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n87), .CK(CLK), .RN(n3), .Q(DOUT[20]), .QN(
        n55) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n86), .CK(CLK), .RN(n3), .Q(DOUT[19]), .QN(
        n54) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n85), .CK(CLK), .RN(n3), .Q(DOUT[18]), .QN(
        n53) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n84), .CK(CLK), .RN(n3), .Q(DOUT[17]), .QN(
        n52) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n83), .CK(CLK), .RN(n3), .Q(DOUT[16]), .QN(
        n51) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n82), .CK(CLK), .RN(n3), .Q(DOUT[15]), .QN(
        n50) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n81), .CK(CLK), .RN(n3), .Q(DOUT[14]), .QN(
        n49) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n80), .CK(CLK), .RN(n3), .Q(DOUT[13]), .QN(
        n48) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n79), .CK(CLK), .RN(n3), .Q(DOUT[12]), .QN(
        n47) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n78), .CK(CLK), .RN(n3), .Q(DOUT[11]), .QN(
        n46) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n77), .CK(CLK), .RN(n2), .Q(DOUT[10]), .QN(
        n45) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n76), .CK(CLK), .RN(n2), .Q(DOUT[9]), .QN(n44)
         );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n75), .CK(CLK), .RN(n2), .Q(DOUT[8]), .QN(n43)
         );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n74), .CK(CLK), .RN(n2), .Q(DOUT[7]), .QN(n42)
         );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n73), .CK(CLK), .RN(n2), .Q(DOUT[6]), .QN(n41)
         );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n72), .CK(CLK), .RN(n2), .Q(DOUT[5]), .QN(n40)
         );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n71), .CK(CLK), .RN(n2), .Q(DOUT[4]), .QN(n39)
         );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n70), .CK(CLK), .RN(n2), .Q(DOUT[3]), .QN(n38)
         );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n69), .CK(CLK), .RN(n2), .Q(DOUT[2]), .QN(n37)
         );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n68), .CK(CLK), .RN(n2), .Q(DOUT[1]), .QN(n36)
         );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n67), .CK(CLK), .RN(n2), .Q(DOUT[0]), .QN(n35)
         );
  BUF_X1 U2 ( .A(RST_AN), .Z(n2) );
  BUF_X1 U3 ( .A(RST_AN), .Z(n3) );
  BUF_X1 U4 ( .A(RST_AN), .Z(n4) );
  OAI22_X1 U5 ( .A1(n35), .A2(EN), .B1(n1), .B2(n101), .ZN(n67) );
  INV_X1 U6 ( .A(DIN[0]), .ZN(n101) );
  OAI22_X1 U7 ( .A1(n36), .A2(EN), .B1(n1), .B2(n100), .ZN(n68) );
  INV_X1 U8 ( .A(DIN[1]), .ZN(n100) );
  OAI22_X1 U9 ( .A1(n37), .A2(EN), .B1(n1), .B2(n99), .ZN(n69) );
  INV_X1 U10 ( .A(DIN[2]), .ZN(n99) );
  OAI22_X1 U11 ( .A1(n38), .A2(EN), .B1(n1), .B2(n34), .ZN(n70) );
  INV_X1 U12 ( .A(DIN[3]), .ZN(n34) );
  OAI22_X1 U13 ( .A1(n39), .A2(EN), .B1(n1), .B2(n33), .ZN(n71) );
  INV_X1 U14 ( .A(DIN[4]), .ZN(n33) );
  OAI22_X1 U15 ( .A1(n40), .A2(EN), .B1(n1), .B2(n32), .ZN(n72) );
  INV_X1 U16 ( .A(DIN[5]), .ZN(n32) );
  OAI22_X1 U17 ( .A1(n41), .A2(EN), .B1(n1), .B2(n31), .ZN(n73) );
  INV_X1 U18 ( .A(DIN[6]), .ZN(n31) );
  OAI22_X1 U19 ( .A1(n42), .A2(EN), .B1(n1), .B2(n30), .ZN(n74) );
  INV_X1 U20 ( .A(DIN[7]), .ZN(n30) );
  OAI22_X1 U21 ( .A1(n43), .A2(EN), .B1(n1), .B2(n29), .ZN(n75) );
  INV_X1 U22 ( .A(DIN[8]), .ZN(n29) );
  OAI22_X1 U23 ( .A1(n44), .A2(EN), .B1(n1), .B2(n28), .ZN(n76) );
  INV_X1 U24 ( .A(DIN[9]), .ZN(n28) );
  OAI22_X1 U25 ( .A1(n45), .A2(EN), .B1(n1), .B2(n27), .ZN(n77) );
  INV_X1 U26 ( .A(DIN[10]), .ZN(n27) );
  OAI22_X1 U27 ( .A1(n46), .A2(EN), .B1(n1), .B2(n26), .ZN(n78) );
  INV_X1 U28 ( .A(DIN[11]), .ZN(n26) );
  OAI22_X1 U29 ( .A1(n47), .A2(EN), .B1(n1), .B2(n25), .ZN(n79) );
  INV_X1 U30 ( .A(DIN[12]), .ZN(n25) );
  OAI22_X1 U31 ( .A1(n48), .A2(EN), .B1(n1), .B2(n24), .ZN(n80) );
  INV_X1 U32 ( .A(DIN[13]), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n49), .A2(EN), .B1(n1), .B2(n23), .ZN(n81) );
  INV_X1 U34 ( .A(DIN[14]), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n50), .A2(EN), .B1(n1), .B2(n22), .ZN(n82) );
  INV_X1 U36 ( .A(DIN[15]), .ZN(n22) );
  OAI22_X1 U37 ( .A1(n51), .A2(EN), .B1(n1), .B2(n21), .ZN(n83) );
  INV_X1 U38 ( .A(DIN[16]), .ZN(n21) );
  OAI22_X1 U39 ( .A1(n52), .A2(EN), .B1(n1), .B2(n20), .ZN(n84) );
  INV_X1 U40 ( .A(DIN[17]), .ZN(n20) );
  OAI22_X1 U41 ( .A1(n66), .A2(EN), .B1(n1), .B2(n102), .ZN(n98) );
  INV_X1 U42 ( .A(DIN[31]), .ZN(n102) );
  INV_X1 U43 ( .A(EN), .ZN(n5) );
  OR2_X1 U44 ( .A1(INIT), .A2(n5), .ZN(n1) );
  INV_X1 U45 ( .A(n1), .ZN(n18) );
  NAND2_X1 U46 ( .A1(DIN[18]), .A2(n18), .ZN(n6) );
  OAI21_X1 U47 ( .B1(n53), .B2(EN), .A(n6), .ZN(n85) );
  NAND2_X1 U48 ( .A1(DIN[19]), .A2(n18), .ZN(n7) );
  OAI21_X1 U49 ( .B1(n54), .B2(EN), .A(n7), .ZN(n86) );
  NAND2_X1 U50 ( .A1(DIN[20]), .A2(n18), .ZN(n8) );
  OAI21_X1 U51 ( .B1(n55), .B2(EN), .A(n8), .ZN(n87) );
  NAND2_X1 U52 ( .A1(DIN[21]), .A2(n18), .ZN(n9) );
  OAI21_X1 U53 ( .B1(n56), .B2(EN), .A(n9), .ZN(n88) );
  NAND2_X1 U54 ( .A1(DIN[22]), .A2(n18), .ZN(n10) );
  OAI21_X1 U55 ( .B1(n57), .B2(EN), .A(n10), .ZN(n89) );
  NAND2_X1 U56 ( .A1(DIN[23]), .A2(n18), .ZN(n11) );
  OAI21_X1 U57 ( .B1(n58), .B2(EN), .A(n11), .ZN(n90) );
  NAND2_X1 U58 ( .A1(DIN[24]), .A2(n18), .ZN(n12) );
  OAI21_X1 U59 ( .B1(n59), .B2(EN), .A(n12), .ZN(n91) );
  NAND2_X1 U60 ( .A1(DIN[25]), .A2(n18), .ZN(n13) );
  OAI21_X1 U61 ( .B1(n60), .B2(EN), .A(n13), .ZN(n92) );
  NAND2_X1 U62 ( .A1(DIN[26]), .A2(n18), .ZN(n14) );
  OAI21_X1 U63 ( .B1(n61), .B2(EN), .A(n14), .ZN(n93) );
  NAND2_X1 U64 ( .A1(DIN[27]), .A2(n18), .ZN(n15) );
  OAI21_X1 U65 ( .B1(n62), .B2(EN), .A(n15), .ZN(n94) );
  NAND2_X1 U66 ( .A1(DIN[28]), .A2(n18), .ZN(n16) );
  OAI21_X1 U67 ( .B1(n63), .B2(EN), .A(n16), .ZN(n95) );
  NAND2_X1 U68 ( .A1(DIN[29]), .A2(n18), .ZN(n17) );
  OAI21_X1 U69 ( .B1(n64), .B2(EN), .A(n17), .ZN(n96) );
  NAND2_X1 U70 ( .A1(DIN[30]), .A2(n18), .ZN(n19) );
  OAI21_X1 U71 ( .B1(n65), .B2(EN), .A(n19), .ZN(n97) );
endmodule


module REG_PIPO_32_00000000_00000000_11 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module RF_ADDR_W5_DATA_W32 ( CLK, RST_AN, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST_AN, ENABLE, RD1, RD2, WR;
  wire   \registers[1][31] , \registers[1][30] , \registers[1][29] ,
         \registers[1][28] , \registers[1][27] , \registers[1][26] ,
         \registers[1][25] , \registers[1][24] , \registers[1][23] ,
         \registers[1][22] , \registers[1][21] , \registers[1][20] ,
         \registers[1][19] , \registers[1][18] , \registers[1][17] ,
         \registers[1][16] , \registers[1][15] , \registers[1][14] ,
         \registers[1][13] , \registers[1][12] , \registers[1][11] ,
         \registers[1][10] , \registers[1][9] , \registers[1][8] ,
         \registers[1][7] , \registers[1][6] , \registers[1][5] ,
         \registers[1][4] , \registers[1][3] , \registers[1][2] ,
         \registers[1][1] , \registers[1][0] , \registers[6][31] ,
         \registers[6][30] , \registers[6][29] , \registers[6][28] ,
         \registers[6][27] , \registers[6][26] , \registers[6][25] ,
         \registers[6][24] , \registers[6][23] , \registers[6][22] ,
         \registers[6][21] , \registers[6][20] , \registers[6][19] ,
         \registers[6][18] , \registers[6][17] , \registers[6][16] ,
         \registers[6][15] , \registers[6][14] , \registers[6][13] ,
         \registers[6][12] , \registers[6][11] , \registers[6][10] ,
         \registers[6][9] , \registers[6][8] , \registers[6][7] ,
         \registers[6][6] , \registers[6][5] , \registers[6][4] ,
         \registers[6][3] , \registers[6][2] , \registers[6][1] ,
         \registers[6][0] , \registers[7][31] , \registers[7][30] ,
         \registers[7][29] , \registers[7][28] , \registers[7][27] ,
         \registers[7][26] , \registers[7][25] , \registers[7][24] ,
         \registers[7][23] , \registers[7][22] , \registers[7][21] ,
         \registers[7][20] , \registers[7][19] , \registers[7][18] ,
         \registers[7][17] , \registers[7][16] , \registers[7][15] ,
         \registers[7][14] , \registers[7][13] , \registers[7][12] ,
         \registers[7][11] , \registers[7][10] , \registers[7][9] ,
         \registers[7][8] , \registers[7][7] , \registers[7][6] ,
         \registers[7][5] , \registers[7][4] , \registers[7][3] ,
         \registers[7][2] , \registers[7][1] , \registers[7][0] ,
         \registers[8][31] , \registers[8][30] , \registers[8][29] ,
         \registers[8][28] , \registers[8][27] , \registers[8][26] ,
         \registers[8][25] , \registers[8][24] , \registers[8][23] ,
         \registers[8][22] , \registers[8][21] , \registers[8][20] ,
         \registers[8][19] , \registers[8][18] , \registers[8][17] ,
         \registers[8][16] , \registers[8][15] , \registers[8][14] ,
         \registers[8][13] , \registers[8][12] , \registers[8][11] ,
         \registers[8][10] , \registers[8][9] , \registers[8][8] ,
         \registers[8][7] , \registers[8][6] , \registers[8][5] ,
         \registers[8][4] , \registers[8][3] , \registers[8][2] ,
         \registers[8][1] , \registers[8][0] , \registers[9][31] ,
         \registers[9][30] , \registers[9][29] , \registers[9][28] ,
         \registers[9][27] , \registers[9][26] , \registers[9][25] ,
         \registers[9][24] , \registers[9][23] , \registers[9][22] ,
         \registers[9][21] , \registers[9][20] , \registers[9][19] ,
         \registers[9][18] , \registers[9][17] , \registers[9][16] ,
         \registers[9][15] , \registers[9][14] , \registers[9][13] ,
         \registers[9][12] , \registers[9][11] , \registers[9][10] ,
         \registers[9][9] , \registers[9][8] , \registers[9][7] ,
         \registers[9][6] , \registers[9][5] , \registers[9][4] ,
         \registers[9][3] , \registers[9][2] , \registers[9][1] ,
         \registers[9][0] , \registers[12][31] , \registers[12][30] ,
         \registers[12][29] , \registers[12][28] , \registers[12][27] ,
         \registers[12][26] , \registers[12][25] , \registers[12][24] ,
         \registers[12][23] , \registers[12][22] , \registers[12][21] ,
         \registers[12][20] , \registers[12][19] , \registers[12][18] ,
         \registers[12][17] , \registers[12][16] , \registers[12][15] ,
         \registers[12][14] , \registers[12][13] , \registers[12][12] ,
         \registers[12][11] , \registers[12][10] , \registers[12][9] ,
         \registers[12][8] , \registers[12][7] , \registers[12][6] ,
         \registers[12][5] , \registers[12][4] , \registers[12][3] ,
         \registers[12][2] , \registers[12][1] , \registers[12][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[18][31] ,
         \registers[18][30] , \registers[18][29] , \registers[18][28] ,
         \registers[18][27] , \registers[18][26] , \registers[18][25] ,
         \registers[18][24] , \registers[18][23] , \registers[18][22] ,
         \registers[18][21] , \registers[18][20] , \registers[18][19] ,
         \registers[18][18] , \registers[18][17] , \registers[18][16] ,
         \registers[18][15] , \registers[18][14] , \registers[18][13] ,
         \registers[18][12] , \registers[18][11] , \registers[18][10] ,
         \registers[18][9] , \registers[18][8] , \registers[18][7] ,
         \registers[18][6] , \registers[18][5] , \registers[18][4] ,
         \registers[18][3] , \registers[18][2] , \registers[18][1] ,
         \registers[18][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[22][31] , \registers[22][30] , \registers[22][29] ,
         \registers[22][28] , \registers[22][27] , \registers[22][26] ,
         \registers[22][25] , \registers[22][24] , \registers[22][23] ,
         \registers[22][22] , \registers[22][21] , \registers[22][20] ,
         \registers[22][19] , \registers[22][18] , \registers[22][17] ,
         \registers[22][16] , \registers[22][15] , \registers[22][14] ,
         \registers[22][13] , \registers[22][12] , \registers[22][11] ,
         \registers[22][10] , \registers[22][9] , \registers[22][8] ,
         \registers[22][7] , \registers[22][6] , \registers[22][5] ,
         \registers[22][4] , \registers[22][3] , \registers[22][2] ,
         \registers[22][1] , \registers[22][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[24][31] , \registers[24][30] ,
         \registers[24][29] , \registers[24][28] , \registers[24][27] ,
         \registers[24][26] , \registers[24][25] , \registers[24][24] ,
         \registers[24][23] , \registers[24][22] , \registers[24][21] ,
         \registers[24][20] , \registers[24][19] , \registers[24][18] ,
         \registers[24][17] , \registers[24][16] , \registers[24][15] ,
         \registers[24][14] , \registers[24][13] , \registers[24][12] ,
         \registers[24][11] , \registers[24][10] , \registers[24][9] ,
         \registers[24][8] , \registers[24][7] , \registers[24][6] ,
         \registers[24][5] , \registers[24][4] , \registers[24][3] ,
         \registers[24][2] , \registers[24][1] , \registers[24][0] ,
         \registers[25][31] , \registers[25][30] , \registers[25][29] ,
         \registers[25][28] , \registers[25][27] , \registers[25][26] ,
         \registers[25][25] , \registers[25][24] , \registers[25][23] ,
         \registers[25][22] , \registers[25][21] , \registers[25][20] ,
         \registers[25][19] , \registers[25][18] , \registers[25][17] ,
         \registers[25][16] , \registers[25][15] , \registers[25][14] ,
         \registers[25][13] , \registers[25][12] , \registers[25][11] ,
         \registers[25][10] , \registers[25][9] , \registers[25][8] ,
         \registers[25][7] , \registers[25][6] , \registers[25][5] ,
         \registers[25][4] , \registers[25][3] , \registers[25][2] ,
         \registers[25][1] , \registers[25][0] , \registers[28][31] ,
         \registers[28][30] , \registers[28][29] , \registers[28][28] ,
         \registers[28][27] , \registers[28][26] , \registers[28][25] ,
         \registers[28][24] , \registers[28][23] , \registers[28][22] ,
         \registers[28][21] , \registers[28][20] , \registers[28][19] ,
         \registers[28][18] , \registers[28][17] , \registers[28][16] ,
         \registers[28][15] , \registers[28][14] , \registers[28][13] ,
         \registers[28][12] , \registers[28][11] , \registers[28][10] ,
         \registers[28][9] , \registers[28][8] , \registers[28][7] ,
         \registers[28][6] , \registers[28][5] , \registers[28][4] ,
         \registers[28][3] , \registers[28][2] , \registers[28][1] ,
         \registers[28][0] , \registers[29][31] , \registers[29][30] ,
         \registers[29][29] , \registers[29][28] , \registers[29][27] ,
         \registers[29][26] , \registers[29][25] , \registers[29][24] ,
         \registers[29][23] , \registers[29][22] , \registers[29][21] ,
         \registers[29][20] , \registers[29][19] , \registers[29][18] ,
         \registers[29][17] , \registers[29][16] , \registers[29][15] ,
         \registers[29][14] , \registers[29][13] , \registers[29][12] ,
         \registers[29][11] , \registers[29][10] , \registers[29][9] ,
         \registers[29][8] , \registers[29][7] , \registers[29][6] ,
         \registers[29][5] , \registers[29][4] , \registers[29][3] ,
         \registers[29][2] , \registers[29][1] , \registers[29][0] , N83, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n1068, n1069, n1070, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1142, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1249, n1251, n1253, n1255,
         n1256, n1257, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1283, n1284, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1352, n1354, n1355, n1356,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1400,
         n1401, n1402, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1423, n1425, n1426,
         n1428, n1430, n1431, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1071, n1113, n1141, n1143, n1248, n1250,
         n1252, n1254, n1258, n1266, n1280, n1281, n1282, n1285, n1320, n1349,
         n1350, n1351, n1353, n1357, n1367, n1387, n1399, n1403, n1404, n1420,
         n1421, n1422, n1424, n1427, n1429, n1432, n1445, n1555, n1556, n1557,
         n1558, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212;

  DFFR_X1 \registers_reg[1][30]  ( .D(n3857), .CK(n4212), .RN(n3694), .Q(
        \registers[1][30] ) );
  DFFR_X1 \registers_reg[1][29]  ( .D(n3856), .CK(n4212), .RN(n3693), .Q(
        \registers[1][29] ) );
  DFFR_X1 \registers_reg[1][28]  ( .D(n3855), .CK(n4212), .RN(n3693), .Q(
        \registers[1][28] ) );
  DFFR_X1 \registers_reg[1][27]  ( .D(n3854), .CK(n4212), .RN(n3693), .Q(
        \registers[1][27] ) );
  DFFR_X1 \registers_reg[1][26]  ( .D(n3853), .CK(n4212), .RN(n3693), .Q(
        \registers[1][26] ) );
  DFFR_X1 \registers_reg[1][25]  ( .D(n3852), .CK(n4212), .RN(n3693), .Q(
        \registers[1][25] ) );
  DFFR_X1 \registers_reg[1][24]  ( .D(n3851), .CK(n4212), .RN(n3693), .Q(
        \registers[1][24] ) );
  DFFR_X1 \registers_reg[1][21]  ( .D(n3848), .CK(n4212), .RN(n3693), .Q(
        \registers[1][21] ) );
  DFFR_X1 \registers_reg[1][20]  ( .D(n3847), .CK(n4212), .RN(n3693), .Q(
        \registers[1][20] ) );
  DFFR_X1 \registers_reg[1][19]  ( .D(n3846), .CK(n4212), .RN(n3693), .Q(
        \registers[1][19] ) );
  DFFR_X1 \registers_reg[1][17]  ( .D(n3844), .CK(n4212), .RN(n3692), .Q(
        \registers[1][17] ) );
  DFFR_X1 \registers_reg[1][16]  ( .D(n3843), .CK(n4212), .RN(n3692), .Q(
        \registers[1][16] ) );
  DFFR_X1 \registers_reg[1][15]  ( .D(n3842), .CK(n4212), .RN(n3692), .Q(
        \registers[1][15] ) );
  DFFR_X1 \registers_reg[1][14]  ( .D(n3841), .CK(n4212), .RN(n3692), .Q(
        \registers[1][14] ) );
  DFFR_X1 \registers_reg[1][13]  ( .D(n3840), .CK(n4212), .RN(n3692), .Q(
        \registers[1][13] ) );
  DFFR_X1 \registers_reg[1][12]  ( .D(n3839), .CK(n4212), .RN(n3692), .Q(
        \registers[1][12] ) );
  DFFR_X1 \registers_reg[1][11]  ( .D(n3838), .CK(n4212), .RN(n3692), .Q(
        \registers[1][11] ) );
  DFFR_X1 \registers_reg[1][10]  ( .D(n3837), .CK(n4212), .RN(n3692), .Q(
        \registers[1][10] ) );
  DFFR_X1 \registers_reg[1][9]  ( .D(n3836), .CK(n4212), .RN(n3692), .Q(
        \registers[1][9] ) );
  DFFR_X1 \registers_reg[1][5]  ( .D(n3832), .CK(n4212), .RN(n3691), .Q(
        \registers[1][5] ) );
  DFFR_X1 \registers_reg[1][4]  ( .D(n3831), .CK(n4212), .RN(n3691), .Q(
        \registers[1][4] ) );
  DFFR_X1 \registers_reg[1][3]  ( .D(n3830), .CK(n4212), .RN(n3691), .Q(
        \registers[1][3] ) );
  DFFR_X1 \registers_reg[1][1]  ( .D(n3828), .CK(n4212), .RN(n3691), .Q(
        \registers[1][1] ) );
  DFFR_X1 \registers_reg[1][0]  ( .D(n3827), .CK(n4212), .RN(n3691), .Q(
        \registers[1][0] ) );
  DFFR_X1 \registers_reg[2][31]  ( .D(n3285), .CK(n4212), .RN(n3691), .QN(n33)
         );
  DFFR_X1 \registers_reg[2][30]  ( .D(n3284), .CK(n4212), .RN(n3691), .QN(n34)
         );
  DFFR_X1 \registers_reg[2][29]  ( .D(n3283), .CK(n4212), .RN(n3691), .QN(n35)
         );
  DFFR_X1 \registers_reg[2][27]  ( .D(n3281), .CK(n4212), .RN(n3690), .QN(n37)
         );
  DFFR_X1 \registers_reg[2][24]  ( .D(n3278), .CK(n4212), .RN(n3690), .QN(n40)
         );
  DFFR_X1 \registers_reg[2][23]  ( .D(n3277), .CK(n4212), .RN(n3690), .QN(n41)
         );
  DFFR_X1 \registers_reg[2][4]  ( .D(n3258), .CK(n4212), .RN(n3688), .QN(n60)
         );
  DFFR_X1 \registers_reg[2][0]  ( .D(n3254), .CK(n4212), .RN(n3688), .QN(n64)
         );
  DFFR_X1 \registers_reg[3][31]  ( .D(n3253), .CK(n4212), .RN(n3688), .QN(n65)
         );
  DFFR_X1 \registers_reg[3][30]  ( .D(n3252), .CK(n4212), .RN(n3688), .QN(n66)
         );
  DFFR_X1 \registers_reg[3][27]  ( .D(n3249), .CK(n4212), .RN(n3687), .QN(n69)
         );
  DFFR_X1 \registers_reg[3][24]  ( .D(n3246), .CK(n4212), .RN(n3687), .QN(n72)
         );
  DFFR_X1 \registers_reg[3][23]  ( .D(n3245), .CK(n4212), .RN(n3687), .QN(n73)
         );
  DFFR_X1 \registers_reg[3][13]  ( .D(n3235), .CK(n4212), .RN(n3686), .QN(n83)
         );
  DFFR_X1 \registers_reg[3][8]  ( .D(n3230), .CK(n4212), .RN(n3686), .QN(n88)
         );
  DFFR_X1 \registers_reg[3][6]  ( .D(n3228), .CK(n4212), .RN(n3686), .QN(n90)
         );
  DFFR_X1 \registers_reg[3][5]  ( .D(n3227), .CK(n4212), .RN(n3685), .QN(n91)
         );
  DFFR_X1 \registers_reg[3][4]  ( .D(n3226), .CK(n4212), .RN(n3685), .QN(n92)
         );
  DFFR_X1 \registers_reg[4][31]  ( .D(n3221), .CK(n4212), .RN(n3685), .QN(n97)
         );
  DFFR_X1 \registers_reg[4][30]  ( .D(n3220), .CK(n4212), .RN(n3685), .QN(n98)
         );
  DFFR_X1 \registers_reg[4][29]  ( .D(n3219), .CK(n4212), .RN(n3685), .QN(n99)
         );
  DFFR_X1 \registers_reg[4][28]  ( .D(n3218), .CK(n4212), .RN(n3685), .QN(n100) );
  DFFR_X1 \registers_reg[4][27]  ( .D(n3217), .CK(n4212), .RN(n3685), .QN(n101) );
  DFFR_X1 \registers_reg[4][26]  ( .D(n3216), .CK(n4212), .RN(n3684), .QN(n102) );
  DFFR_X1 \registers_reg[4][25]  ( .D(n3215), .CK(n4212), .RN(n3684), .QN(n103) );
  DFFR_X1 \registers_reg[4][24]  ( .D(n3214), .CK(n4212), .RN(n3684), .QN(n104) );
  DFFR_X1 \registers_reg[4][23]  ( .D(n3213), .CK(n4212), .RN(n3684), .QN(n105) );
  DFFR_X1 \registers_reg[4][21]  ( .D(n3211), .CK(n4212), .RN(n3684), .QN(n107) );
  DFFR_X1 \registers_reg[4][20]  ( .D(n3210), .CK(n4212), .RN(n3684), .QN(n108) );
  DFFR_X1 \registers_reg[4][19]  ( .D(n3209), .CK(n4212), .RN(n3684), .QN(n109) );
  DFFR_X1 \registers_reg[4][16]  ( .D(n3206), .CK(n4212), .RN(n3684), .QN(n112) );
  DFFR_X1 \registers_reg[4][13]  ( .D(n3203), .CK(n4212), .RN(n3683), .QN(n115) );
  DFFR_X1 \registers_reg[4][9]  ( .D(n3199), .CK(n4212), .RN(n3683), .QN(n119)
         );
  DFFR_X1 \registers_reg[4][8]  ( .D(n3198), .CK(n4212), .RN(n3683), .QN(n120)
         );
  DFFR_X1 \registers_reg[4][7]  ( .D(n3197), .CK(n4212), .RN(n3683), .QN(n121)
         );
  DFFR_X1 \registers_reg[4][6]  ( .D(n3196), .CK(n4212), .RN(n3683), .QN(n122)
         );
  DFFR_X1 \registers_reg[4][5]  ( .D(n3195), .CK(n4212), .RN(n3683), .QN(n123)
         );
  DFFR_X1 \registers_reg[4][4]  ( .D(n3194), .CK(n4212), .RN(n3682), .QN(n124)
         );
  DFFR_X1 \registers_reg[4][3]  ( .D(n3193), .CK(n4212), .RN(n3682), .QN(n125)
         );
  DFFR_X1 \registers_reg[4][2]  ( .D(n3192), .CK(n4212), .RN(n3682), .QN(n126)
         );
  DFFR_X1 \registers_reg[5][31]  ( .D(n3189), .CK(n4212), .RN(n3682), .QN(n129) );
  DFFR_X1 \registers_reg[5][30]  ( .D(n3188), .CK(n4212), .RN(n3682), .QN(n130) );
  DFFR_X1 \registers_reg[5][29]  ( .D(n3187), .CK(n4212), .RN(n3682), .QN(n131) );
  DFFR_X1 \registers_reg[5][27]  ( .D(n3185), .CK(n4212), .RN(n3682), .QN(n133) );
  DFFR_X1 \registers_reg[5][24]  ( .D(n3182), .CK(n4212), .RN(n3681), .QN(n136) );
  DFFR_X1 \registers_reg[5][23]  ( .D(n3181), .CK(n4212), .RN(n3681), .QN(n137) );
  DFFR_X1 \registers_reg[5][8]  ( .D(n3166), .CK(n4212), .RN(n3680), .QN(n152)
         );
  DFFR_X1 \registers_reg[5][4]  ( .D(n3162), .CK(n4212), .RN(n3680), .QN(n156)
         );
  DFFR_X1 \registers_reg[5][0]  ( .D(n3158), .CK(n4212), .RN(n3679), .QN(n160)
         );
  DFFR_X1 \registers_reg[6][22]  ( .D(n3881), .CK(n4212), .RN(n3678), .Q(
        \registers[6][22] ) );
  DFFR_X1 \registers_reg[6][19]  ( .D(n3878), .CK(n4212), .RN(n3678), .Q(
        \registers[6][19] ) );
  DFFR_X1 \registers_reg[7][31]  ( .D(n3922), .CK(n4212), .RN(n3676), .Q(
        \registers[7][31] ) );
  DFFR_X1 \registers_reg[7][30]  ( .D(n3921), .CK(n4212), .RN(n3676), .Q(
        \registers[7][30] ) );
  DFFR_X1 \registers_reg[7][29]  ( .D(n3920), .CK(n4212), .RN(n3676), .Q(
        \registers[7][29] ) );
  DFFR_X1 \registers_reg[7][28]  ( .D(n3919), .CK(n4212), .RN(n3676), .Q(
        \registers[7][28] ) );
  DFFR_X1 \registers_reg[7][27]  ( .D(n3918), .CK(n4212), .RN(n3676), .Q(
        \registers[7][27] ) );
  DFFR_X1 \registers_reg[7][26]  ( .D(n3917), .CK(n4212), .RN(n3676), .Q(
        \registers[7][26] ) );
  DFFR_X1 \registers_reg[7][25]  ( .D(n3916), .CK(n4212), .RN(n3676), .Q(
        \registers[7][25] ) );
  DFFR_X1 \registers_reg[7][24]  ( .D(n3915), .CK(n4212), .RN(n3676), .Q(
        \registers[7][24] ) );
  DFFR_X1 \registers_reg[7][23]  ( .D(n3914), .CK(n4212), .RN(n3675), .Q(
        \registers[7][23] ) );
  DFFR_X1 \registers_reg[7][22]  ( .D(n3913), .CK(n4212), .RN(n3675), .Q(
        \registers[7][22] ) );
  DFFR_X1 \registers_reg[7][21]  ( .D(n3912), .CK(n4212), .RN(n3675), .Q(
        \registers[7][21] ) );
  DFFR_X1 \registers_reg[7][20]  ( .D(n3911), .CK(n4212), .RN(n3675), .Q(
        \registers[7][20] ) );
  DFFR_X1 \registers_reg[7][19]  ( .D(n3910), .CK(n4212), .RN(n3675), .Q(
        \registers[7][19] ) );
  DFFR_X1 \registers_reg[7][18]  ( .D(n3909), .CK(n4212), .RN(n3675), .Q(
        \registers[7][18] ) );
  DFFR_X1 \registers_reg[7][17]  ( .D(n3908), .CK(n4212), .RN(n3675), .Q(
        \registers[7][17] ) );
  DFFR_X1 \registers_reg[7][16]  ( .D(n3907), .CK(n4212), .RN(n3675), .Q(
        \registers[7][16] ) );
  DFFR_X1 \registers_reg[7][15]  ( .D(n3906), .CK(n4212), .RN(n3675), .Q(
        \registers[7][15] ) );
  DFFR_X1 \registers_reg[7][14]  ( .D(n3905), .CK(n4212), .RN(n3675), .Q(
        \registers[7][14] ) );
  DFFR_X1 \registers_reg[7][13]  ( .D(n3904), .CK(n4212), .RN(n3675), .Q(
        \registers[7][13] ) );
  DFFR_X1 \registers_reg[7][12]  ( .D(n3903), .CK(n4212), .RN(n3674), .Q(
        \registers[7][12] ) );
  DFFR_X1 \registers_reg[7][11]  ( .D(n3902), .CK(n4212), .RN(n3674), .Q(
        \registers[7][11] ) );
  DFFR_X1 \registers_reg[7][10]  ( .D(n3901), .CK(n4212), .RN(n3674), .Q(
        \registers[7][10] ) );
  DFFR_X1 \registers_reg[7][9]  ( .D(n3900), .CK(n4212), .RN(n3674), .Q(
        \registers[7][9] ) );
  DFFR_X1 \registers_reg[7][8]  ( .D(n3899), .CK(n4212), .RN(n3674), .Q(
        \registers[7][8] ) );
  DFFR_X1 \registers_reg[7][7]  ( .D(n3898), .CK(n4212), .RN(n3674), .Q(
        \registers[7][7] ) );
  DFFR_X1 \registers_reg[7][6]  ( .D(n3897), .CK(n4212), .RN(n3674), .Q(
        \registers[7][6] ) );
  DFFR_X1 \registers_reg[7][5]  ( .D(n3896), .CK(n4212), .RN(n3674), .Q(
        \registers[7][5] ) );
  DFFR_X1 \registers_reg[7][4]  ( .D(n3895), .CK(n4212), .RN(n3674), .Q(
        \registers[7][4] ) );
  DFFR_X1 \registers_reg[7][3]  ( .D(n3894), .CK(n4212), .RN(n3674), .Q(
        \registers[7][3] ) );
  DFFR_X1 \registers_reg[7][2]  ( .D(n3893), .CK(n4212), .RN(n3674), .Q(
        \registers[7][2] ) );
  DFFR_X1 \registers_reg[7][1]  ( .D(n3892), .CK(n4212), .RN(n3673), .Q(
        \registers[7][1] ) );
  DFFR_X1 \registers_reg[7][0]  ( .D(n3891), .CK(n4212), .RN(n3673), .Q(
        \registers[7][0] ) );
  DFFR_X1 \registers_reg[8][31]  ( .D(n3742), .CK(n4212), .RN(n3673), .Q(
        \registers[8][31] ) );
  DFFR_X1 \registers_reg[8][30]  ( .D(n3741), .CK(n4212), .RN(n3673), .Q(
        \registers[8][30] ) );
  DFFR_X1 \registers_reg[8][29]  ( .D(n3740), .CK(n4212), .RN(n3673), .Q(
        \registers[8][29] ) );
  DFFR_X1 \registers_reg[8][28]  ( .D(n3739), .CK(n4212), .RN(n3673), .Q(
        \registers[8][28] ) );
  DFFR_X1 \registers_reg[8][27]  ( .D(n3738), .CK(n4212), .RN(n3673), .Q(
        \registers[8][27] ) );
  DFFR_X1 \registers_reg[8][26]  ( .D(n3737), .CK(n4212), .RN(n3673), .Q(
        \registers[8][26] ) );
  DFFR_X1 \registers_reg[8][25]  ( .D(n3736), .CK(n4212), .RN(n3673), .Q(
        \registers[8][25] ) );
  DFFR_X1 \registers_reg[8][24]  ( .D(n3735), .CK(n4212), .RN(n3673), .Q(
        \registers[8][24] ) );
  DFFR_X1 \registers_reg[8][23]  ( .D(n3734), .CK(n4212), .RN(n3673), .Q(
        \registers[8][23] ) );
  DFFR_X1 \registers_reg[8][22]  ( .D(n3733), .CK(n4212), .RN(n3672), .Q(
        \registers[8][22] ) );
  DFFR_X1 \registers_reg[8][21]  ( .D(n3732), .CK(n4212), .RN(n3672), .Q(
        \registers[8][21] ) );
  DFFR_X1 \registers_reg[8][20]  ( .D(n3731), .CK(n4212), .RN(n3672), .Q(
        \registers[8][20] ) );
  DFFR_X1 \registers_reg[8][19]  ( .D(n3730), .CK(n4212), .RN(n3672), .Q(
        \registers[8][19] ) );
  DFFR_X1 \registers_reg[8][18]  ( .D(n3729), .CK(n4212), .RN(n3672), .Q(
        \registers[8][18] ) );
  DFFR_X1 \registers_reg[8][17]  ( .D(n3728), .CK(n4212), .RN(n3672), .Q(
        \registers[8][17] ) );
  DFFR_X1 \registers_reg[8][16]  ( .D(n3727), .CK(n4212), .RN(n3672), .Q(
        \registers[8][16] ) );
  DFFR_X1 \registers_reg[8][15]  ( .D(n3726), .CK(n4212), .RN(n3672), .Q(
        \registers[8][15] ) );
  DFFR_X1 \registers_reg[8][14]  ( .D(n3725), .CK(n4212), .RN(n3672), .Q(
        \registers[8][14] ) );
  DFFR_X1 \registers_reg[8][13]  ( .D(n3724), .CK(n4212), .RN(n3672), .Q(
        \registers[8][13] ) );
  DFFR_X1 \registers_reg[8][12]  ( .D(n3723), .CK(n4212), .RN(n3672), .Q(
        \registers[8][12] ) );
  DFFR_X1 \registers_reg[8][11]  ( .D(n3722), .CK(n4212), .RN(n3671), .Q(
        \registers[8][11] ) );
  DFFR_X1 \registers_reg[8][10]  ( .D(n3721), .CK(n4212), .RN(n3671), .Q(
        \registers[8][10] ) );
  DFFR_X1 \registers_reg[8][9]  ( .D(n3720), .CK(n4212), .RN(n3671), .Q(
        \registers[8][9] ) );
  DFFR_X1 \registers_reg[8][8]  ( .D(n3719), .CK(n4212), .RN(n3671), .Q(
        \registers[8][8] ) );
  DFFR_X1 \registers_reg[8][7]  ( .D(n3718), .CK(n4212), .RN(n3671), .Q(
        \registers[8][7] ) );
  DFFR_X1 \registers_reg[8][6]  ( .D(n3717), .CK(n4212), .RN(n3671), .Q(
        \registers[8][6] ) );
  DFFR_X1 \registers_reg[8][5]  ( .D(n3716), .CK(n4212), .RN(n3671), .Q(
        \registers[8][5] ) );
  DFFR_X1 \registers_reg[8][4]  ( .D(n3715), .CK(n4212), .RN(n3671), .Q(
        \registers[8][4] ) );
  DFFR_X1 \registers_reg[8][3]  ( .D(n3714), .CK(n4212), .RN(n3671), .Q(
        \registers[8][3] ) );
  DFFR_X1 \registers_reg[8][2]  ( .D(n3713), .CK(n4212), .RN(n3671), .Q(
        \registers[8][2] ) );
  DFFR_X1 \registers_reg[8][1]  ( .D(n3712), .CK(n4212), .RN(n3671), .Q(
        \registers[8][1] ) );
  DFFR_X1 \registers_reg[8][0]  ( .D(n3711), .CK(n4212), .RN(n3670), .Q(
        \registers[8][0] ) );
  DFFR_X1 \registers_reg[9][31]  ( .D(n3768), .CK(n4212), .RN(n3670), .Q(
        \registers[9][31] ) );
  DFFR_X1 \registers_reg[9][30]  ( .D(n3767), .CK(n4212), .RN(n3670), .Q(
        \registers[9][30] ) );
  DFFR_X1 \registers_reg[9][27]  ( .D(n3764), .CK(n4212), .RN(n3670), .Q(
        \registers[9][27] ) );
  DFFR_X1 \registers_reg[9][21]  ( .D(n3759), .CK(n4212), .RN(n3669), .Q(
        \registers[9][21] ) );
  DFFR_X1 \registers_reg[9][20]  ( .D(n3758), .CK(n4212), .RN(n3669), .Q(
        \registers[9][20] ) );
  DFFR_X1 \registers_reg[9][19]  ( .D(n3757), .CK(n4212), .RN(n3669), .Q(
        \registers[9][19] ) );
  DFFR_X1 \registers_reg[9][16]  ( .D(n3754), .CK(n4212), .RN(n3669), .Q(
        \registers[9][16] ) );
  DFFR_X1 \registers_reg[9][15]  ( .D(n3753), .CK(n4212), .RN(n3669), .Q(
        \registers[9][15] ) );
  DFFR_X1 \registers_reg[9][14]  ( .D(n3752), .CK(n4212), .RN(n3669), .Q(
        \registers[9][14] ) );
  DFFR_X1 \registers_reg[9][13]  ( .D(n3751), .CK(n4212), .RN(n3669), .Q(
        \registers[9][13] ) );
  DFFR_X1 \registers_reg[9][12]  ( .D(n3750), .CK(n4212), .RN(n3669), .Q(
        \registers[9][12] ) );
  DFFR_X1 \registers_reg[9][11]  ( .D(n3749), .CK(n4212), .RN(n3669), .Q(
        \registers[9][11] ) );
  DFFR_X1 \registers_reg[9][10]  ( .D(n3748), .CK(n4212), .RN(n3668), .Q(
        \registers[9][10] ) );
  DFFR_X1 \registers_reg[9][9]  ( .D(n245), .CK(n4212), .RN(n3668), .Q(
        \registers[9][9] ), .QN(n246) );
  DFFR_X1 \registers_reg[9][8]  ( .D(n3747), .CK(n4212), .RN(n3668), .Q(
        \registers[9][8] ) );
  DFFR_X1 \registers_reg[9][7]  ( .D(n3746), .CK(n4212), .RN(n3668), .Q(
        \registers[9][7] ) );
  DFFR_X1 \registers_reg[9][6]  ( .D(n255), .CK(n4212), .RN(n3668), .Q(
        \registers[9][6] ), .QN(n256) );
  DFFR_X1 \registers_reg[9][5]  ( .D(n3745), .CK(n4212), .RN(n3668), .Q(
        \registers[9][5] ) );
  DFFR_X1 \registers_reg[9][3]  ( .D(n3744), .CK(n4212), .RN(n3668), .Q(
        \registers[9][3] ) );
  DFFR_X1 \registers_reg[9][2]  ( .D(n3743), .CK(n4212), .RN(n3668), .Q(
        \registers[9][2] ) );
  DFFR_X1 \registers_reg[9][0]  ( .D(n260), .CK(n4212), .RN(n3668), .Q(
        \registers[9][0] ), .QN(n261) );
  DFFR_X1 \registers_reg[10][31]  ( .D(n3157), .CK(n4212), .RN(n3667), .QN(
        n289) );
  DFFR_X1 \registers_reg[11][31]  ( .D(n3125), .CK(n4212), .RN(n3665), .QN(
        n321) );
  DFFR_X1 \registers_reg[11][30]  ( .D(n3124), .CK(n4212), .RN(n3664), .QN(
        n322) );
  DFFR_X1 \registers_reg[11][29]  ( .D(n3123), .CK(n4212), .RN(n3664), .QN(
        n323) );
  DFFR_X1 \registers_reg[11][27]  ( .D(n3121), .CK(n4212), .RN(n3664), .QN(
        n325) );
  DFFR_X1 \registers_reg[11][24]  ( .D(n3118), .CK(n4212), .RN(n3664), .QN(
        n328) );
  DFFR_X1 \registers_reg[11][23]  ( .D(n3117), .CK(n4212), .RN(n3664), .QN(
        n329) );
  DFFR_X1 \registers_reg[11][13]  ( .D(n3107), .CK(n4212), .RN(n3663), .QN(
        n339) );
  DFFR_X1 \registers_reg[11][4]  ( .D(n3098), .CK(n4212), .RN(n3662), .QN(n348) );
  DFFR_X1 \registers_reg[12][31]  ( .D(n3796), .CK(n4212), .RN(n3662), .Q(
        \registers[12][31] ) );
  DFFR_X1 \registers_reg[12][30]  ( .D(n3795), .CK(n4212), .RN(n3662), .Q(
        \registers[12][30] ) );
  DFFR_X1 \registers_reg[12][29]  ( .D(n3794), .CK(n4212), .RN(n3661), .Q(
        \registers[12][29] ) );
  DFFR_X1 \registers_reg[12][26]  ( .D(n3791), .CK(n4212), .RN(n3661), .Q(
        \registers[12][26] ) );
  DFFR_X1 \registers_reg[12][25]  ( .D(n3790), .CK(n4212), .RN(n3661), .Q(
        \registers[12][25] ) );
  DFFR_X1 \registers_reg[12][24]  ( .D(n3789), .CK(n4212), .RN(n3661), .Q(
        \registers[12][24] ) );
  DFFR_X1 \registers_reg[12][23]  ( .D(n3788), .CK(n4212), .RN(n3661), .Q(
        \registers[12][23] ) );
  DFFR_X1 \registers_reg[12][22]  ( .D(n3787), .CK(n4212), .RN(n3661), .Q(
        \registers[12][22] ) );
  DFFR_X1 \registers_reg[12][21]  ( .D(n3786), .CK(n4212), .RN(n3661), .Q(
        \registers[12][21] ) );
  DFFR_X1 \registers_reg[12][20]  ( .D(n3785), .CK(n4212), .RN(n3661), .Q(
        \registers[12][20] ) );
  DFFR_X1 \registers_reg[12][19]  ( .D(n3784), .CK(n4212), .RN(n3661), .Q(
        \registers[12][19] ) );
  DFFR_X1 \registers_reg[12][18]  ( .D(n3783), .CK(n4212), .RN(n3660), .Q(
        \registers[12][18] ) );
  DFFR_X1 \registers_reg[12][17]  ( .D(n3782), .CK(n4212), .RN(n3660), .Q(
        \registers[12][17] ) );
  DFFR_X1 \registers_reg[12][16]  ( .D(n209), .CK(n4212), .RN(n3660), .Q(
        \registers[12][16] ), .QN(n210) );
  DFFR_X1 \registers_reg[12][15]  ( .D(n399), .CK(n4212), .RN(n3660), .Q(
        \registers[12][15] ) );
  DFFR_X1 \registers_reg[12][14]  ( .D(n3781), .CK(n4212), .RN(n3660), .Q(
        \registers[12][14] ) );
  DFFR_X1 \registers_reg[12][13]  ( .D(n3780), .CK(n4212), .RN(n3660), .Q(
        \registers[12][13] ) );
  DFFR_X1 \registers_reg[12][12]  ( .D(n3779), .CK(n4212), .RN(n3660), .Q(
        \registers[12][12] ) );
  DFFR_X1 \registers_reg[12][11]  ( .D(n413), .CK(n4212), .RN(n3660), .Q(
        \registers[12][11] ), .QN(n414) );
  DFFR_X1 \registers_reg[12][10]  ( .D(n3778), .CK(n4212), .RN(n3660), .Q(
        \registers[12][10] ) );
  DFFR_X1 \registers_reg[12][9]  ( .D(n3777), .CK(n4212), .RN(n3660), .Q(
        \registers[12][9] ) );
  DFFR_X1 \registers_reg[12][8]  ( .D(n3776), .CK(n4212), .RN(n3660), .Q(
        \registers[12][8] ) );
  DFFR_X1 \registers_reg[12][7]  ( .D(n3775), .CK(n4212), .RN(n3659), .Q(
        \registers[12][7] ) );
  DFFR_X1 \registers_reg[12][5]  ( .D(n3773), .CK(n4212), .RN(n3659), .Q(
        \registers[12][5] ) );
  DFFR_X1 \registers_reg[12][4]  ( .D(n3772), .CK(n4212), .RN(n3659), .Q(
        \registers[12][4] ) );
  DFFR_X1 \registers_reg[12][3]  ( .D(n3771), .CK(n4212), .RN(n3659), .Q(
        \registers[12][3] ) );
  DFFR_X1 \registers_reg[12][2]  ( .D(n3770), .CK(n4212), .RN(n3659), .Q(
        \registers[12][2] ) );
  DFFR_X1 \registers_reg[12][1]  ( .D(n3769), .CK(n4212), .RN(n3659), .Q(
        \registers[12][1] ) );
  DFFR_X1 \registers_reg[13][30]  ( .D(n3825), .CK(n4212), .RN(n3659), .Q(
        \registers[13][30] ) );
  DFFR_X1 \registers_reg[13][29]  ( .D(n3824), .CK(n4212), .RN(n3659), .Q(
        \registers[13][29] ) );
  DFFR_X1 \registers_reg[13][28]  ( .D(n3823), .CK(n4212), .RN(n3658), .Q(
        \registers[13][28] ) );
  DFFR_X1 \registers_reg[13][27]  ( .D(n3822), .CK(n4212), .RN(n3658), .Q(
        \registers[13][27] ) );
  DFFR_X1 \registers_reg[13][26]  ( .D(n3821), .CK(n4212), .RN(n3658), .Q(
        \registers[13][26] ) );
  DFFR_X1 \registers_reg[13][25]  ( .D(n3820), .CK(n4212), .RN(n3658), .Q(
        \registers[13][25] ) );
  DFFR_X1 \registers_reg[13][24]  ( .D(n3819), .CK(n4212), .RN(n3658), .Q(
        \registers[13][24] ) );
  DFFR_X1 \registers_reg[13][23]  ( .D(n3818), .CK(n4212), .RN(n3658), .Q(
        \registers[13][23] ) );
  DFFR_X1 \registers_reg[13][20]  ( .D(n3815), .CK(n4212), .RN(n3658), .Q(
        \registers[13][20] ) );
  DFFR_X1 \registers_reg[13][19]  ( .D(n3814), .CK(n4212), .RN(n3658), .Q(
        \registers[13][19] ) );
  DFFR_X1 \registers_reg[13][17]  ( .D(n3812), .CK(n4212), .RN(n3657), .Q(
        \registers[13][17] ) );
  DFFR_X1 \registers_reg[13][16]  ( .D(n3811), .CK(n4212), .RN(n3657), .Q(
        \registers[13][16] ) );
  DFFR_X1 \registers_reg[13][15]  ( .D(n3810), .CK(n4212), .RN(n3657), .Q(
        \registers[13][15] ) );
  DFFR_X1 \registers_reg[13][13]  ( .D(n3808), .CK(n4212), .RN(n3657), .Q(
        \registers[13][13] ) );
  DFFR_X1 \registers_reg[13][9]  ( .D(n3805), .CK(n4212), .RN(n3657), .Q(
        \registers[13][9] ) );
  DFFR_X1 \registers_reg[13][7]  ( .D(n3803), .CK(n4212), .RN(n3657), .Q(
        \registers[13][7] ) );
  DFFR_X1 \registers_reg[13][6]  ( .D(n3802), .CK(n4212), .RN(n3656), .Q(
        \registers[13][6] ) );
  DFFR_X1 \registers_reg[13][3]  ( .D(n3799), .CK(n4212), .RN(n3656), .Q(
        \registers[13][3] ) );
  DFFR_X1 \registers_reg[13][1]  ( .D(n3798), .CK(n4212), .RN(n3656), .Q(
        \registers[13][1] ) );
  DFFR_X1 \registers_reg[13][0]  ( .D(n3797), .CK(n4212), .RN(n3656), .Q(
        \registers[13][0] ) );
  DFFR_X1 \registers_reg[14][31]  ( .D(n3093), .CK(n4212), .RN(n3656), .QN(
        n417) );
  DFFR_X1 \registers_reg[14][30]  ( .D(n3092), .CK(n4212), .RN(n3656), .QN(
        n418) );
  DFFR_X1 \registers_reg[14][29]  ( .D(n3091), .CK(n4212), .RN(n3656), .QN(
        n419) );
  DFFR_X1 \registers_reg[14][28]  ( .D(n3090), .CK(n4212), .RN(n3656), .QN(
        n420) );
  DFFR_X1 \registers_reg[14][27]  ( .D(n3089), .CK(n4212), .RN(n3655), .QN(
        n421) );
  DFFR_X1 \registers_reg[14][26]  ( .D(n3088), .CK(n4212), .RN(n3655), .QN(
        n422) );
  DFFR_X1 \registers_reg[14][25]  ( .D(n3087), .CK(n4212), .RN(n3655), .QN(
        n423) );
  DFFR_X1 \registers_reg[14][24]  ( .D(n3086), .CK(n4212), .RN(n3655), .QN(
        n424) );
  DFFR_X1 \registers_reg[14][23]  ( .D(n3085), .CK(n4212), .RN(n3655), .QN(
        n425) );
  DFFR_X1 \registers_reg[14][21]  ( .D(n3083), .CK(n4212), .RN(n3655), .QN(
        n427) );
  DFFR_X1 \registers_reg[14][20]  ( .D(n3082), .CK(n4212), .RN(n3655), .QN(
        n428) );
  DFFR_X1 \registers_reg[14][19]  ( .D(n3081), .CK(n4212), .RN(n3655), .QN(
        n429) );
  DFFR_X1 \registers_reg[14][16]  ( .D(n3078), .CK(n4212), .RN(n3654), .QN(
        n432) );
  DFFR_X1 \registers_reg[14][13]  ( .D(n3075), .CK(n4212), .RN(n3654), .QN(
        n435) );
  DFFR_X1 \registers_reg[14][9]  ( .D(n3071), .CK(n4212), .RN(n3654), .QN(n439) );
  DFFR_X1 \registers_reg[14][8]  ( .D(n3070), .CK(n4212), .RN(n3654), .QN(n440) );
  DFFR_X1 \registers_reg[14][7]  ( .D(n3069), .CK(n4212), .RN(n3654), .QN(n441) );
  DFFR_X1 \registers_reg[14][6]  ( .D(n3068), .CK(n4212), .RN(n3654), .QN(n442) );
  DFFR_X1 \registers_reg[14][5]  ( .D(n3067), .CK(n4212), .RN(n3653), .QN(n443) );
  DFFR_X1 \registers_reg[14][4]  ( .D(n3066), .CK(n4212), .RN(n3653), .QN(n444) );
  DFFR_X1 \registers_reg[14][3]  ( .D(n3065), .CK(n4212), .RN(n3653), .QN(n445) );
  DFFR_X1 \registers_reg[14][2]  ( .D(n3064), .CK(n4212), .RN(n3653), .QN(n446) );
  DFFR_X1 \registers_reg[15][31]  ( .D(n3061), .CK(n4212), .RN(n3653), .QN(
        n449) );
  DFFR_X1 \registers_reg[15][30]  ( .D(n3060), .CK(n4212), .RN(n3653), .QN(
        n450) );
  DFFR_X1 \registers_reg[15][28]  ( .D(n3058), .CK(n4212), .RN(n3653), .QN(
        n452) );
  DFFR_X1 \registers_reg[15][26]  ( .D(n3056), .CK(n4212), .RN(n3652), .QN(
        n454) );
  DFFR_X1 \registers_reg[15][25]  ( .D(n3055), .CK(n4212), .RN(n3652), .QN(
        n455) );
  DFFR_X1 \registers_reg[15][22]  ( .D(n3052), .CK(n4212), .RN(n3652), .QN(
        n458) );
  DFFR_X1 \registers_reg[15][18]  ( .D(n3048), .CK(n4212), .RN(n3652), .QN(
        n462) );
  DFFR_X1 \registers_reg[15][12]  ( .D(n3042), .CK(n4212), .RN(n3651), .QN(
        n468) );
  DFFR_X1 \registers_reg[15][11]  ( .D(n3041), .CK(n4212), .RN(n3651), .QN(
        n469) );
  DFFR_X1 \registers_reg[15][10]  ( .D(n3040), .CK(n4212), .RN(n3651), .QN(
        n470) );
  DFFR_X1 \registers_reg[15][5]  ( .D(n3035), .CK(n4212), .RN(n3651), .QN(n475) );
  DFFR_X1 \registers_reg[15][4]  ( .D(n3034), .CK(n4212), .RN(n3650), .QN(n476) );
  DFFR_X1 \registers_reg[15][1]  ( .D(n3031), .CK(n4212), .RN(n3650), .QN(n479) );
  DFFR_X1 \registers_reg[15][0]  ( .D(n3030), .CK(n4212), .RN(n3650), .QN(n480) );
  DFFR_X1 \registers_reg[16][31]  ( .D(n3029), .CK(n4212), .RN(n3650), .QN(
        n481) );
  DFFR_X1 \registers_reg[16][29]  ( .D(n3027), .CK(n4212), .RN(n3650), .QN(
        n483) );
  DFFR_X1 \registers_reg[16][28]  ( .D(n3026), .CK(n4212), .RN(n3650), .QN(
        n484) );
  DFFR_X1 \registers_reg[16][27]  ( .D(n3025), .CK(n4212), .RN(n3650), .QN(
        n485) );
  DFFR_X1 \registers_reg[16][26]  ( .D(n3024), .CK(n4212), .RN(n3650), .QN(
        n486) );
  DFFR_X1 \registers_reg[16][25]  ( .D(n3023), .CK(n4212), .RN(n3649), .QN(
        n487) );
  DFFR_X1 \registers_reg[16][24]  ( .D(n3022), .CK(n4212), .RN(n3649), .QN(
        n488) );
  DFFR_X1 \registers_reg[16][23]  ( .D(n3021), .CK(n4212), .RN(n3649), .QN(
        n489) );
  DFFR_X1 \registers_reg[16][21]  ( .D(n3019), .CK(n4212), .RN(n3649), .QN(
        n491) );
  DFFR_X1 \registers_reg[16][20]  ( .D(n3018), .CK(n4212), .RN(n3649), .QN(
        n492) );
  DFFR_X1 \registers_reg[16][19]  ( .D(n3017), .CK(n4212), .RN(n3649), .QN(
        n493) );
  DFFR_X1 \registers_reg[16][18]  ( .D(n3016), .CK(n4212), .RN(n3649), .QN(
        n494) );
  DFFR_X1 \registers_reg[16][17]  ( .D(n3015), .CK(n4212), .RN(n3649), .QN(
        n495) );
  DFFR_X1 \registers_reg[16][16]  ( .D(n3014), .CK(n4212), .RN(n3649), .QN(
        n496) );
  DFFR_X1 \registers_reg[16][15]  ( .D(n3013), .CK(n4212), .RN(n3649), .QN(
        n497) );
  DFFR_X1 \registers_reg[16][14]  ( .D(n3012), .CK(n4212), .RN(n3648), .QN(
        n498) );
  DFFR_X1 \registers_reg[16][12]  ( .D(n3010), .CK(n4212), .RN(n3648), .QN(
        n500) );
  DFFR_X1 \registers_reg[16][11]  ( .D(n3009), .CK(n4212), .RN(n3648), .QN(
        n501) );
  DFFR_X1 \registers_reg[16][10]  ( .D(n3008), .CK(n4212), .RN(n3648), .QN(
        n502) );
  DFFR_X1 \registers_reg[16][9]  ( .D(n3007), .CK(n4212), .RN(n3648), .QN(n503) );
  DFFR_X1 \registers_reg[16][7]  ( .D(n3005), .CK(n4212), .RN(n3648), .QN(n505) );
  DFFR_X1 \registers_reg[16][6]  ( .D(n3004), .CK(n4212), .RN(n3648), .QN(n506) );
  DFFR_X1 \registers_reg[16][5]  ( .D(n3003), .CK(n4212), .RN(n3648), .QN(n507) );
  DFFR_X1 \registers_reg[16][3]  ( .D(n3001), .CK(n4212), .RN(n3647), .QN(n509) );
  DFFR_X1 \registers_reg[16][2]  ( .D(n3000), .CK(n4212), .RN(n3647), .QN(n510) );
  DFFR_X1 \registers_reg[16][0]  ( .D(n2998), .CK(n4212), .RN(n3647), .QN(n512) );
  DFFR_X1 \registers_reg[18][31]  ( .D(n3954), .CK(n4212), .RN(n3644), .Q(
        \registers[18][31] ) );
  DFFR_X1 \registers_reg[18][30]  ( .D(n3953), .CK(n4212), .RN(n3644), .Q(
        \registers[18][30] ) );
  DFFR_X1 \registers_reg[18][19]  ( .D(n3942), .CK(n4212), .RN(n3643), .Q(
        \registers[18][19] ) );
  DFFR_X1 \registers_reg[18][3]  ( .D(n580), .CK(n4212), .RN(n3642), .Q(
        \registers[18][3] ), .QN(n581) );
  DFFR_X1 \registers_reg[19][31]  ( .D(n3985), .CK(n4212), .RN(n3641), .Q(
        \registers[19][31] ) );
  DFFR_X1 \registers_reg[19][28]  ( .D(n3982), .CK(n4212), .RN(n3641), .Q(
        \registers[19][28] ) );
  DFFR_X1 \registers_reg[19][27]  ( .D(n3981), .CK(n4212), .RN(n3641), .Q(
        \registers[19][27] ) );
  DFFR_X1 \registers_reg[19][26]  ( .D(n3980), .CK(n4212), .RN(n3641), .Q(
        \registers[19][26] ) );
  DFFR_X1 \registers_reg[19][24]  ( .D(n3978), .CK(n4212), .RN(n3641), .Q(
        \registers[19][24] ) );
  DFFR_X1 \registers_reg[19][22]  ( .D(n3976), .CK(n4212), .RN(n3640), .Q(
        \registers[19][22] ) );
  DFFR_X1 \registers_reg[19][21]  ( .D(n3975), .CK(n4212), .RN(n3640), .Q(
        \registers[19][21] ) );
  DFFR_X1 \registers_reg[19][20]  ( .D(n3974), .CK(n4212), .RN(n3640), .Q(
        \registers[19][20] ) );
  DFFR_X1 \registers_reg[19][19]  ( .D(n3973), .CK(n4212), .RN(n3640), .Q(
        \registers[19][19] ) );
  DFFR_X1 \registers_reg[19][17]  ( .D(n3971), .CK(n4212), .RN(n3640), .Q(
        \registers[19][17] ) );
  DFFR_X1 \registers_reg[19][16]  ( .D(n3970), .CK(n4212), .RN(n3640), .Q(
        \registers[19][16] ) );
  DFFR_X1 \registers_reg[19][15]  ( .D(n3969), .CK(n4212), .RN(n3640), .Q(
        \registers[19][15] ) );
  DFFR_X1 \registers_reg[19][11]  ( .D(n3965), .CK(n4212), .RN(n3639), .Q(
        \registers[19][11] ) );
  DFFR_X1 \registers_reg[19][10]  ( .D(n3964), .CK(n4212), .RN(n3639), .Q(
        \registers[19][10] ) );
  DFFR_X1 \registers_reg[19][9]  ( .D(n3963), .CK(n4212), .RN(n3639), .Q(
        \registers[19][9] ) );
  DFFR_X1 \registers_reg[19][7]  ( .D(n3961), .CK(n4212), .RN(n3639), .Q(
        \registers[19][7] ) );
  DFFR_X1 \registers_reg[19][5]  ( .D(n3959), .CK(n4212), .RN(n3639), .Q(
        \registers[19][5] ) );
  DFFR_X1 \registers_reg[19][4]  ( .D(n3958), .CK(n4212), .RN(n3639), .Q(
        \registers[19][4] ) );
  DFFR_X1 \registers_reg[19][3]  ( .D(n3957), .CK(n4212), .RN(n3639), .Q(
        \registers[19][3] ) );
  DFFR_X1 \registers_reg[19][2]  ( .D(n3956), .CK(n4212), .RN(n3639), .Q(
        \registers[19][2] ) );
  DFFR_X1 \registers_reg[19][1]  ( .D(n582), .CK(n4212), .RN(n3639), .Q(
        \registers[19][1] ), .QN(n583) );
  DFFR_X1 \registers_reg[19][0]  ( .D(n3955), .CK(n4212), .RN(n3638), .Q(
        \registers[19][0] ) );
  DFFR_X1 \registers_reg[20][31]  ( .D(n2965), .CK(n4212), .RN(n3638), .QN(
        n609) );
  DFFR_X1 \registers_reg[20][30]  ( .D(n2964), .CK(n4212), .RN(n3638), .QN(
        n610) );
  DFFR_X1 \registers_reg[20][29]  ( .D(n2963), .CK(n4212), .RN(n3638), .QN(
        n611) );
  DFFR_X1 \registers_reg[20][28]  ( .D(n2962), .CK(n4212), .RN(n3638), .QN(
        n612) );
  DFFR_X1 \registers_reg[20][27]  ( .D(n2961), .CK(n4212), .RN(n3638), .QN(
        n613) );
  DFFR_X1 \registers_reg[20][23]  ( .D(n2957), .CK(n4212), .RN(n3638), .QN(
        n617) );
  DFFR_X1 \registers_reg[20][22]  ( .D(n2956), .CK(n4212), .RN(n3638), .QN(
        n618) );
  DFFR_X1 \registers_reg[20][20]  ( .D(n2954), .CK(n4212), .RN(n3637), .QN(
        n620) );
  DFFR_X1 \registers_reg[20][19]  ( .D(n2953), .CK(n4212), .RN(n3637), .QN(
        n621) );
  DFFR_X1 \registers_reg[20][18]  ( .D(n2952), .CK(n4212), .RN(n3637), .QN(
        n622) );
  DFFR_X1 \registers_reg[20][17]  ( .D(n2951), .CK(n4212), .RN(n3637), .QN(
        n623) );
  DFFR_X1 \registers_reg[20][13]  ( .D(n2947), .CK(n4212), .RN(n3637), .QN(
        n627) );
  DFFR_X1 \registers_reg[20][12]  ( .D(n2946), .CK(n4212), .RN(n3637), .QN(
        n628) );
  DFFR_X1 \registers_reg[20][11]  ( .D(n2945), .CK(n4212), .RN(n3637), .QN(
        n629) );
  DFFR_X1 \registers_reg[20][4]  ( .D(n2938), .CK(n4212), .RN(n3636), .QN(n636) );
  DFFR_X1 \registers_reg[20][3]  ( .D(n2937), .CK(n4212), .RN(n3636), .QN(n637) );
  DFFR_X1 \registers_reg[20][0]  ( .D(n2934), .CK(n4212), .RN(n3636), .QN(n640) );
  DFFR_X1 \registers_reg[21][31]  ( .D(n2933), .CK(n4212), .RN(n3635), .QN(
        n641) );
  DFFR_X1 \registers_reg[21][30]  ( .D(n2932), .CK(n4212), .RN(n3635), .QN(
        n642) );
  DFFR_X1 \registers_reg[21][29]  ( .D(n2931), .CK(n4212), .RN(n3635), .QN(
        n643) );
  DFFR_X1 \registers_reg[21][27]  ( .D(n2929), .CK(n4212), .RN(n3635), .QN(
        n645) );
  DFFR_X1 \registers_reg[21][24]  ( .D(n2926), .CK(n4212), .RN(n3635), .QN(
        n648) );
  DFFR_X1 \registers_reg[21][23]  ( .D(n2925), .CK(n4212), .RN(n3635), .QN(
        n649) );
  DFFR_X1 \registers_reg[21][14]  ( .D(n2916), .CK(n4212), .RN(n3634), .QN(
        n658) );
  DFFR_X1 \registers_reg[21][13]  ( .D(n2915), .CK(n4212), .RN(n3634), .QN(
        n659) );
  DFFR_X1 \registers_reg[21][8]  ( .D(n2910), .CK(n4212), .RN(n3633), .QN(n664) );
  DFFR_X1 \registers_reg[21][6]  ( .D(n2908), .CK(n4212), .RN(n3633), .QN(n666) );
  DFFR_X1 \registers_reg[21][4]  ( .D(n2906), .CK(n4212), .RN(n3633), .QN(n668) );
  DFFR_X1 \registers_reg[21][0]  ( .D(n2902), .CK(n4212), .RN(n3633), .QN(n672) );
  DFFR_X1 \registers_reg[22][31]  ( .D(n232), .CK(n4212), .RN(n3633), .Q(
        \registers[22][31] ), .QN(n233) );
  DFFR_X1 \registers_reg[22][30]  ( .D(n4010), .CK(n4212), .RN(n3632), .Q(
        \registers[22][30] ) );
  DFFR_X1 \registers_reg[22][29]  ( .D(n4009), .CK(n4212), .RN(n3632), .Q(
        \registers[22][29] ) );
  DFFR_X1 \registers_reg[22][28]  ( .D(n4008), .CK(n4212), .RN(n3632), .Q(
        \registers[22][28] ) );
  DFFR_X1 \registers_reg[22][27]  ( .D(n4007), .CK(n4212), .RN(n3632), .Q(
        \registers[22][27] ) );
  DFFR_X1 \registers_reg[22][26]  ( .D(n4006), .CK(n4212), .RN(n3632), .Q(
        \registers[22][26] ) );
  DFFR_X1 \registers_reg[22][25]  ( .D(n4005), .CK(n4212), .RN(n3632), .Q(
        \registers[22][25] ) );
  DFFR_X1 \registers_reg[22][24]  ( .D(n4004), .CK(n4212), .RN(n3632), .Q(
        \registers[22][24] ) );
  DFFR_X1 \registers_reg[22][23]  ( .D(n4003), .CK(n4212), .RN(n3632), .Q(
        \registers[22][23] ) );
  DFFR_X1 \registers_reg[22][22]  ( .D(n4002), .CK(n4212), .RN(n3632), .Q(
        \registers[22][22] ) );
  DFFR_X1 \registers_reg[22][21]  ( .D(n4001), .CK(n4212), .RN(n3632), .Q(
        \registers[22][21] ) );
  DFFR_X1 \registers_reg[22][20]  ( .D(n4000), .CK(n4212), .RN(n3632), .Q(
        \registers[22][20] ) );
  DFFR_X1 \registers_reg[22][19]  ( .D(n3999), .CK(n4212), .RN(n3631), .Q(
        \registers[22][19] ) );
  DFFR_X1 \registers_reg[22][18]  ( .D(n3998), .CK(n4212), .RN(n3631), .Q(
        \registers[22][18] ) );
  DFFR_X1 \registers_reg[22][16]  ( .D(n3997), .CK(n4212), .RN(n3631), .Q(
        \registers[22][16] ) );
  DFFR_X1 \registers_reg[22][15]  ( .D(n3996), .CK(n4212), .RN(n3631), .Q(
        \registers[22][15] ) );
  DFFR_X1 \registers_reg[22][14]  ( .D(n3995), .CK(n4212), .RN(n3631), .Q(
        \registers[22][14] ) );
  DFFR_X1 \registers_reg[22][13]  ( .D(n3994), .CK(n4212), .RN(n3631), .Q(
        \registers[22][13] ) );
  DFFR_X1 \registers_reg[22][12]  ( .D(n3993), .CK(n4212), .RN(n3631), .Q(
        \registers[22][12] ) );
  DFFR_X1 \registers_reg[22][11]  ( .D(n3992), .CK(n4212), .RN(n3631), .Q(
        \registers[22][11] ) );
  DFFR_X1 \registers_reg[22][10]  ( .D(n3991), .CK(n4212), .RN(n3631), .Q(
        \registers[22][10] ) );
  DFFR_X1 \registers_reg[22][8]  ( .D(n3990), .CK(n4212), .RN(n3630), .Q(
        \registers[22][8] ) );
  DFFR_X1 \registers_reg[22][7]  ( .D(n3989), .CK(n4212), .RN(n3630), .Q(
        \registers[22][7] ) );
  DFFR_X1 \registers_reg[22][6]  ( .D(n3988), .CK(n4212), .RN(n3630), .Q(
        \registers[22][6] ) );
  DFFR_X1 \registers_reg[22][4]  ( .D(n3987), .CK(n4212), .RN(n3630), .Q(
        \registers[22][4] ) );
  DFFR_X1 \registers_reg[22][3]  ( .D(n415), .CK(n4212), .RN(n3630), .Q(
        \registers[22][3] ), .QN(n416) );
  DFFR_X1 \registers_reg[22][2]  ( .D(n3986), .CK(n4212), .RN(n3630), .Q(
        \registers[22][2] ) );
  DFFR_X1 \registers_reg[22][0]  ( .D(n26), .CK(n4212), .RN(n3630), .Q(
        \registers[22][0] ), .QN(n27) );
  DFFR_X1 \registers_reg[23][31]  ( .D(n4042), .CK(n4212), .RN(n3630), .Q(
        \registers[23][31] ) );
  DFFR_X1 \registers_reg[23][30]  ( .D(n4041), .CK(n4212), .RN(n3630), .Q(
        \registers[23][30] ) );
  DFFR_X1 \registers_reg[23][29]  ( .D(n4040), .CK(n4212), .RN(n3629), .Q(
        \registers[23][29] ) );
  DFFR_X1 \registers_reg[23][28]  ( .D(n4039), .CK(n4212), .RN(n3629), .Q(
        \registers[23][28] ) );
  DFFR_X1 \registers_reg[23][26]  ( .D(n4037), .CK(n4212), .RN(n3629), .Q(
        \registers[23][26] ) );
  DFFR_X1 \registers_reg[23][25]  ( .D(n4036), .CK(n4212), .RN(n3629), .Q(
        \registers[23][25] ) );
  DFFR_X1 \registers_reg[23][24]  ( .D(n4035), .CK(n4212), .RN(n3629), .Q(
        \registers[23][24] ) );
  DFFR_X1 \registers_reg[23][23]  ( .D(n4034), .CK(n4212), .RN(n3629), .Q(
        \registers[23][23] ) );
  DFFR_X1 \registers_reg[23][21]  ( .D(n4032), .CK(n4212), .RN(n3629), .Q(
        \registers[23][21] ) );
  DFFR_X1 \registers_reg[23][20]  ( .D(n4031), .CK(n4212), .RN(n3629), .Q(
        \registers[23][20] ) );
  DFFR_X1 \registers_reg[23][19]  ( .D(n4030), .CK(n4212), .RN(n3629), .Q(
        \registers[23][19] ) );
  DFFR_X1 \registers_reg[23][18]  ( .D(n4029), .CK(n4212), .RN(n3628), .Q(
        \registers[23][18] ) );
  DFFR_X1 \registers_reg[23][15]  ( .D(n4026), .CK(n4212), .RN(n3628), .Q(
        \registers[23][15] ) );
  DFFR_X1 \registers_reg[23][14]  ( .D(n4025), .CK(n4212), .RN(n3628), .Q(
        \registers[23][14] ) );
  DFFR_X1 \registers_reg[23][12]  ( .D(n4023), .CK(n4212), .RN(n3628), .Q(
        \registers[23][12] ) );
  DFFR_X1 \registers_reg[23][10]  ( .D(n4021), .CK(n4212), .RN(n3628), .Q(
        \registers[23][10] ) );
  DFFR_X1 \registers_reg[23][9]  ( .D(n4020), .CK(n4212), .RN(n3628), .Q(
        \registers[23][9] ) );
  DFFR_X1 \registers_reg[23][8]  ( .D(n4019), .CK(n4212), .RN(n3628), .Q(
        \registers[23][8] ) );
  DFFR_X1 \registers_reg[23][7]  ( .D(n4018), .CK(n4212), .RN(n3627), .Q(
        \registers[23][7] ) );
  DFFR_X1 \registers_reg[23][6]  ( .D(n4017), .CK(n4212), .RN(n3627), .Q(
        \registers[23][6] ) );
  DFFR_X1 \registers_reg[23][5]  ( .D(n4016), .CK(n4212), .RN(n3627), .Q(
        \registers[23][5] ) );
  DFFR_X1 \registers_reg[23][3]  ( .D(n4014), .CK(n4212), .RN(n3627), .Q(
        \registers[23][3] ) );
  DFFR_X1 \registers_reg[23][2]  ( .D(n4013), .CK(n4212), .RN(n3627), .Q(
        \registers[23][2] ) );
  DFFR_X1 \registers_reg[23][1]  ( .D(n4012), .CK(n4212), .RN(n3627), .Q(
        \registers[23][1] ) );
  DFFR_X1 \registers_reg[23][0]  ( .D(n4011), .CK(n4212), .RN(n3627), .Q(
        \registers[23][0] ) );
  DFFR_X1 \registers_reg[24][30]  ( .D(n4073), .CK(n4212), .RN(n3627), .Q(
        \registers[24][30] ) );
  DFFR_X1 \registers_reg[24][29]  ( .D(n4072), .CK(n4212), .RN(n3627), .Q(
        \registers[24][29] ) );
  DFFR_X1 \registers_reg[24][28]  ( .D(n4071), .CK(n4212), .RN(n3626), .Q(
        \registers[24][28] ) );
  DFFR_X1 \registers_reg[24][26]  ( .D(n4069), .CK(n4212), .RN(n3626), .Q(
        \registers[24][26] ) );
  DFFR_X1 \registers_reg[24][24]  ( .D(n4067), .CK(n4212), .RN(n3626), .Q(
        \registers[24][24] ) );
  DFFR_X1 \registers_reg[24][23]  ( .D(n4066), .CK(n4212), .RN(n3626), .Q(
        \registers[24][23] ) );
  DFFR_X1 \registers_reg[24][20]  ( .D(n4063), .CK(n4212), .RN(n3626), .Q(
        \registers[24][20] ) );
  DFFR_X1 \registers_reg[24][19]  ( .D(n4062), .CK(n4212), .RN(n3626), .Q(
        \registers[24][19] ) );
  DFFR_X1 \registers_reg[24][18]  ( .D(n4061), .CK(n4212), .RN(n3626), .Q(
        \registers[24][18] ) );
  DFFR_X1 \registers_reg[24][17]  ( .D(n4060), .CK(n4212), .RN(n3625), .Q(
        \registers[24][17] ) );
  DFFR_X1 \registers_reg[24][16]  ( .D(n4059), .CK(n4212), .RN(n3625), .Q(
        \registers[24][16] ) );
  DFFR_X1 \registers_reg[24][15]  ( .D(n4058), .CK(n4212), .RN(n3625), .Q(
        \registers[24][15] ) );
  DFFR_X1 \registers_reg[24][13]  ( .D(n4056), .CK(n4212), .RN(n3625), .Q(
        \registers[24][13] ) );
  DFFR_X1 \registers_reg[24][12]  ( .D(n4055), .CK(n4212), .RN(n3625), .Q(
        \registers[24][12] ) );
  DFFR_X1 \registers_reg[24][11]  ( .D(n4054), .CK(n4212), .RN(n3625), .Q(
        \registers[24][11] ) );
  DFFR_X1 \registers_reg[24][8]  ( .D(n4051), .CK(n4212), .RN(n3625), .Q(
        \registers[24][8] ) );
  DFFR_X1 \registers_reg[24][6]  ( .D(n4049), .CK(n4212), .RN(n3624), .Q(
        \registers[24][6] ) );
  DFFR_X1 \registers_reg[24][3]  ( .D(n4046), .CK(n4212), .RN(n3624), .Q(
        \registers[24][3] ) );
  DFFR_X1 \registers_reg[24][2]  ( .D(n4045), .CK(n4212), .RN(n3624), .Q(
        \registers[24][2] ) );
  DFFR_X1 \registers_reg[24][0]  ( .D(n4043), .CK(n4212), .RN(n3624), .Q(
        \registers[24][0] ) );
  DFFR_X1 \registers_reg[25][31]  ( .D(n4106), .CK(n4212), .RN(n3624), .Q(
        \registers[25][31] ) );
  DFFR_X1 \registers_reg[25][30]  ( .D(n4105), .CK(n4212), .RN(n3624), .Q(
        \registers[25][30] ) );
  DFFR_X1 \registers_reg[25][29]  ( .D(n4104), .CK(n4212), .RN(n3624), .Q(
        \registers[25][29] ) );
  DFFR_X1 \registers_reg[25][28]  ( .D(n4103), .CK(n4212), .RN(n3624), .Q(
        \registers[25][28] ) );
  DFFR_X1 \registers_reg[25][27]  ( .D(n4102), .CK(n4212), .RN(n3623), .Q(
        \registers[25][27] ) );
  DFFR_X1 \registers_reg[25][26]  ( .D(n4101), .CK(n4212), .RN(n3623), .Q(
        \registers[25][26] ) );
  DFFR_X1 \registers_reg[25][25]  ( .D(n4100), .CK(n4212), .RN(n3623), .Q(
        \registers[25][25] ) );
  DFFR_X1 \registers_reg[25][24]  ( .D(n4099), .CK(n4212), .RN(n3623), .Q(
        \registers[25][24] ) );
  DFFR_X1 \registers_reg[25][23]  ( .D(n4098), .CK(n4212), .RN(n3623), .Q(
        \registers[25][23] ) );
  DFFR_X1 \registers_reg[25][22]  ( .D(n4097), .CK(n4212), .RN(n3623), .Q(
        \registers[25][22] ) );
  DFFR_X1 \registers_reg[25][21]  ( .D(n4096), .CK(n4212), .RN(n3623), .Q(
        \registers[25][21] ) );
  DFFR_X1 \registers_reg[25][20]  ( .D(n4095), .CK(n4212), .RN(n3623), .Q(
        \registers[25][20] ) );
  DFFR_X1 \registers_reg[25][19]  ( .D(n4094), .CK(n4212), .RN(n3623), .Q(
        \registers[25][19] ) );
  DFFR_X1 \registers_reg[25][18]  ( .D(n4093), .CK(n4212), .RN(n3623), .Q(
        \registers[25][18] ) );
  DFFR_X1 \registers_reg[25][17]  ( .D(n4092), .CK(n4212), .RN(n3623), .Q(
        \registers[25][17] ) );
  DFFR_X1 \registers_reg[25][16]  ( .D(n4091), .CK(n4212), .RN(n3622), .Q(
        \registers[25][16] ) );
  DFFR_X1 \registers_reg[25][15]  ( .D(n4090), .CK(n4212), .RN(n3622), .Q(
        \registers[25][15] ) );
  DFFR_X1 \registers_reg[25][14]  ( .D(n4089), .CK(n4212), .RN(n3622), .Q(
        \registers[25][14] ) );
  DFFR_X1 \registers_reg[25][13]  ( .D(n4088), .CK(n4212), .RN(n3622), .Q(
        \registers[25][13] ) );
  DFFR_X1 \registers_reg[25][12]  ( .D(n4087), .CK(n4212), .RN(n3622), .Q(
        \registers[25][12] ) );
  DFFR_X1 \registers_reg[25][11]  ( .D(n4086), .CK(n4212), .RN(n3622), .Q(
        \registers[25][11] ) );
  DFFR_X1 \registers_reg[25][10]  ( .D(n4085), .CK(n4212), .RN(n3622), .Q(
        \registers[25][10] ) );
  DFFR_X1 \registers_reg[25][9]  ( .D(n4084), .CK(n4212), .RN(n3622), .Q(
        \registers[25][9] ) );
  DFFR_X1 \registers_reg[25][8]  ( .D(n4083), .CK(n4212), .RN(n3622), .Q(
        \registers[25][8] ) );
  DFFR_X1 \registers_reg[25][6]  ( .D(n4081), .CK(n4212), .RN(n3622), .Q(
        \registers[25][6] ) );
  DFFR_X1 \registers_reg[25][5]  ( .D(n4080), .CK(n4212), .RN(n3621), .Q(
        \registers[25][5] ) );
  DFFR_X1 \registers_reg[25][4]  ( .D(n4079), .CK(n4212), .RN(n3621), .Q(
        \registers[25][4] ) );
  DFFR_X1 \registers_reg[25][3]  ( .D(n4078), .CK(n4212), .RN(n3621), .Q(
        \registers[25][3] ) );
  DFFR_X1 \registers_reg[25][2]  ( .D(n4077), .CK(n4212), .RN(n3621), .Q(
        \registers[25][2] ) );
  DFFR_X1 \registers_reg[25][1]  ( .D(n4076), .CK(n4212), .RN(n3621), .Q(
        \registers[25][1] ) );
  DFFR_X1 \registers_reg[25][0]  ( .D(n4075), .CK(n4212), .RN(n3621), .Q(
        \registers[25][0] ) );
  DFFR_X1 \registers_reg[26][31]  ( .D(n2901), .CK(n4212), .RN(n3621), .QN(
        n801) );
  DFFR_X1 \registers_reg[26][4]  ( .D(n2874), .CK(n4212), .RN(n3618), .QN(n828) );
  DFFR_X1 \registers_reg[27][31]  ( .D(n2869), .CK(n4212), .RN(n3618), .QN(
        n833) );
  DFFR_X1 \registers_reg[27][30]  ( .D(n2868), .CK(n4212), .RN(n3618), .QN(
        n834) );
  DFFR_X1 \registers_reg[27][29]  ( .D(n2867), .CK(n4212), .RN(n3618), .QN(
        n835) );
  DFFR_X1 \registers_reg[27][28]  ( .D(n2866), .CK(n4212), .RN(n3618), .QN(
        n836) );
  DFFR_X1 \registers_reg[27][27]  ( .D(n2865), .CK(n4212), .RN(n3618), .QN(
        n837) );
  DFFR_X1 \registers_reg[27][26]  ( .D(n2864), .CK(n4212), .RN(n3618), .QN(
        n838) );
  DFFR_X1 \registers_reg[27][25]  ( .D(n2863), .CK(n4212), .RN(n3617), .QN(
        n839) );
  DFFR_X1 \registers_reg[27][24]  ( .D(n2862), .CK(n4212), .RN(n3617), .QN(
        n840) );
  DFFR_X1 \registers_reg[27][22]  ( .D(n2860), .CK(n4212), .RN(n3617), .QN(
        n842) );
  DFFR_X1 \registers_reg[27][21]  ( .D(n2859), .CK(n4212), .RN(n3617), .QN(
        n843) );
  DFFR_X1 \registers_reg[27][20]  ( .D(n2858), .CK(n4212), .RN(n3617), .QN(
        n844) );
  DFFR_X1 \registers_reg[27][18]  ( .D(n2856), .CK(n4212), .RN(n3617), .QN(
        n846) );
  DFFR_X1 \registers_reg[27][17]  ( .D(n2855), .CK(n4212), .RN(n3617), .QN(
        n847) );
  DFFR_X1 \registers_reg[27][16]  ( .D(n2854), .CK(n4212), .RN(n3617), .QN(
        n848) );
  DFFR_X1 \registers_reg[27][12]  ( .D(n2850), .CK(n4212), .RN(n3616), .QN(
        n852) );
  DFFR_X1 \registers_reg[27][11]  ( .D(n2849), .CK(n4212), .RN(n3616), .QN(
        n853) );
  DFFR_X1 \registers_reg[27][10]  ( .D(n2848), .CK(n4212), .RN(n3616), .QN(
        n854) );
  DFFR_X1 \registers_reg[27][9]  ( .D(n2847), .CK(n4212), .RN(n3616), .QN(n855) );
  DFFR_X1 \registers_reg[27][8]  ( .D(n2846), .CK(n4212), .RN(n3616), .QN(n856) );
  DFFR_X1 \registers_reg[27][6]  ( .D(n2844), .CK(n4212), .RN(n3616), .QN(n858) );
  DFFR_X1 \registers_reg[27][5]  ( .D(n2843), .CK(n4212), .RN(n3616), .QN(n859) );
  DFFR_X1 \registers_reg[27][4]  ( .D(n2842), .CK(n4212), .RN(n3616), .QN(n860) );
  DFFR_X1 \registers_reg[27][2]  ( .D(n2840), .CK(n4212), .RN(n3615), .QN(n862) );
  DFFR_X1 \registers_reg[27][1]  ( .D(n2839), .CK(n4212), .RN(n3615), .QN(n863) );
  DFFR_X1 \registers_reg[27][0]  ( .D(n2838), .CK(n4212), .RN(n3615), .QN(n864) );
  DFFR_X1 \registers_reg[28][31]  ( .D(n4137), .CK(n4212), .RN(n3615), .Q(
        \registers[28][31] ) );
  DFFR_X1 \registers_reg[28][30]  ( .D(n4136), .CK(n4212), .RN(n3615), .Q(
        \registers[28][30] ) );
  DFFR_X1 \registers_reg[28][28]  ( .D(n4134), .CK(n4212), .RN(n3615), .Q(
        \registers[28][28] ) );
  DFFR_X1 \registers_reg[28][27]  ( .D(n4133), .CK(n4212), .RN(n3615), .Q(
        \registers[28][27] ) );
  DFFR_X1 \registers_reg[28][24]  ( .D(n4130), .CK(n4212), .RN(n3614), .Q(
        \registers[28][24] ) );
  DFFR_X1 \registers_reg[28][23]  ( .D(n4129), .CK(n4212), .RN(n3614), .Q(
        \registers[28][23] ) );
  DFFR_X1 \registers_reg[28][22]  ( .D(n4128), .CK(n4212), .RN(n3614), .Q(
        \registers[28][22] ) );
  DFFR_X1 \registers_reg[28][20]  ( .D(n4126), .CK(n4212), .RN(n3614), .Q(
        \registers[28][20] ) );
  DFFR_X1 \registers_reg[28][19]  ( .D(n4125), .CK(n4212), .RN(n3614), .Q(
        \registers[28][19] ) );
  DFFR_X1 \registers_reg[28][18]  ( .D(n4124), .CK(n4212), .RN(n3614), .Q(
        \registers[28][18] ) );
  DFFR_X1 \registers_reg[28][16]  ( .D(n4122), .CK(n4212), .RN(n3614), .Q(
        \registers[28][16] ) );
  DFFR_X1 \registers_reg[28][12]  ( .D(n4118), .CK(n4212), .RN(n3613), .Q(
        \registers[28][12] ) );
  DFFR_X1 \registers_reg[28][10]  ( .D(n4116), .CK(n4212), .RN(n3613), .Q(
        \registers[28][10] ) );
  DFFR_X1 \registers_reg[28][8]  ( .D(n4114), .CK(n4212), .RN(n3613), .Q(
        \registers[28][8] ) );
  DFFR_X1 \registers_reg[28][6]  ( .D(n4112), .CK(n4212), .RN(n3613), .Q(
        \registers[28][6] ) );
  DFFR_X1 \registers_reg[28][5]  ( .D(n601), .CK(n4212), .RN(n3613), .Q(
        \registers[28][5] ), .QN(n602) );
  DFFR_X1 \registers_reg[28][4]  ( .D(n4111), .CK(n4212), .RN(n3613), .Q(
        \registers[28][4] ) );
  DFFR_X1 \registers_reg[28][3]  ( .D(n4110), .CK(n4212), .RN(n3613), .Q(
        \registers[28][3] ) );
  DFFR_X1 \registers_reg[28][2]  ( .D(n4109), .CK(n4212), .RN(n3612), .Q(
        \registers[28][2] ) );
  DFFR_X1 \registers_reg[28][0]  ( .D(n4107), .CK(n4212), .RN(n3612), .Q(
        \registers[28][0] ) );
  DFFR_X1 \registers_reg[29][19]  ( .D(n4157), .CK(n4212), .RN(n3611), .Q(
        \registers[29][19] ) );
  DFFR_X1 \registers_reg[29][3]  ( .D(n4141), .CK(n4212), .RN(n3610), .Q(
        \registers[29][3] ) );
  DFFR_X1 \registers_reg[30][31]  ( .D(n2837), .CK(n4212), .RN(n3609), .QN(
        n929) );
  DFFR_X1 \registers_reg[30][28]  ( .D(n2834), .CK(n4212), .RN(n3609), .QN(
        n932) );
  DFFR_X1 \registers_reg[30][26]  ( .D(n2832), .CK(n4212), .RN(n3609), .QN(
        n934) );
  DFFR_X1 \registers_reg[30][23]  ( .D(n2829), .CK(n4212), .RN(n3609), .QN(
        n937) );
  DFFR_X1 \registers_reg[30][21]  ( .D(n2827), .CK(n4212), .RN(n3608), .QN(
        n939) );
  DFFR_X1 \registers_reg[30][20]  ( .D(n2826), .CK(n4212), .RN(n3608), .QN(
        n940) );
  DFFR_X1 \registers_reg[30][16]  ( .D(n2822), .CK(n4212), .RN(n3608), .QN(
        n944) );
  DFFR_X1 \registers_reg[30][13]  ( .D(n2819), .CK(n4212), .RN(n3608), .QN(
        n947) );
  DFFR_X1 \registers_reg[30][6]  ( .D(n2812), .CK(n4212), .RN(n3607), .QN(n954) );
  DFFR_X1 \registers_reg[30][4]  ( .D(n2810), .CK(n4212), .RN(n3607), .QN(n956) );
  DFFR_X1 \registers_reg[30][2]  ( .D(n2808), .CK(n4212), .RN(n3607), .QN(n958) );
  DFFR_X1 \registers_reg[30][0]  ( .D(n2806), .CK(n4212), .RN(n3606), .Q(n30), 
        .QN(n960) );
  DFFR_X1 \registers_reg[31][31]  ( .D(n2805), .CK(n4212), .RN(n3606), .QN(
        n961) );
  DFFR_X1 \registers_reg[31][30]  ( .D(n2804), .CK(n4212), .RN(n3606), .QN(
        n962) );
  DFFR_X1 \registers_reg[31][29]  ( .D(n2803), .CK(n4212), .RN(n3606), .QN(
        n963) );
  DFFR_X1 \registers_reg[31][28]  ( .D(n2802), .CK(n4212), .RN(n3606), .QN(
        n964) );
  DFFR_X1 \registers_reg[31][27]  ( .D(n2801), .CK(n4212), .RN(n3606), .QN(
        n965) );
  DFFR_X1 \registers_reg[31][26]  ( .D(n2800), .CK(n4212), .RN(n3606), .QN(
        n966) );
  DFFR_X1 \registers_reg[31][25]  ( .D(n2799), .CK(n4212), .RN(n3606), .QN(
        n967) );
  DFFR_X1 \registers_reg[31][24]  ( .D(n2798), .CK(n4212), .RN(n3606), .QN(
        n968) );
  DFFR_X1 \registers_reg[31][23]  ( .D(n2797), .CK(n4212), .RN(n3606), .QN(
        n969) );
  DFFR_X1 \registers_reg[31][21]  ( .D(n2795), .CK(n4212), .RN(n3605), .QN(
        n971) );
  DFFR_X1 \registers_reg[31][20]  ( .D(n2794), .CK(n4212), .RN(n3605), .QN(
        n972) );
  DFFR_X1 \registers_reg[31][9]  ( .D(n2783), .CK(n4212), .RN(n3604), .QN(n983) );
  DFFR_X1 \registers_reg[31][4]  ( .D(n2778), .CK(n4212), .RN(n3604), .QN(n988) );
  DFFR_X1 \registers_reg[31][3]  ( .D(n2777), .CK(n4212), .RN(n3604), .QN(n989) );
  DFFR_X1 \registers_reg[31][2]  ( .D(n2776), .CK(n4212), .RN(n3604), .QN(n990) );
  DLH_X1 \OUT1_reg[31]  ( .G(n3589), .D(N217), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n3589), .D(N216), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n3589), .D(N215), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n3589), .D(N214), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n3589), .D(N213), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n3589), .D(N212), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n3589), .D(N211), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n3589), .D(N210), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n3589), .D(N209), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n3589), .D(N208), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n3590), .D(N207), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n3590), .D(N206), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n3590), .D(N205), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n3590), .D(N204), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n3590), .D(N203), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n3590), .D(N202), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n3590), .D(N201), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n3590), .D(N200), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n3590), .D(N199), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n3590), .D(N198), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n3591), .D(N197), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n3591), .D(N196), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n3591), .D(N195), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n3591), .D(N194), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n3591), .D(N193), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n3591), .D(N192), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n3591), .D(N191), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n3591), .D(N190), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n3591), .D(N189), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n3591), .D(N188), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n3592), .D(N187), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n3592), .D(N186), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(n3585), .D(N352), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n3585), .D(N351), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n3585), .D(N350), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n3585), .D(N349), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n3585), .D(N348), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n3585), .D(N347), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n3585), .D(N346), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n3585), .D(N345), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n3585), .D(N344), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n3585), .D(N343), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n3586), .D(N342), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n3586), .D(N341), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n3586), .D(N340), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n3586), .D(N339), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n3586), .D(N338), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n3586), .D(N337), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n3586), .D(N336), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n3586), .D(N335), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n3586), .D(N334), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n3586), .D(N333), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n3587), .D(N332), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n3587), .D(N331), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n3587), .D(N330), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n3587), .D(N329), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n3587), .D(N328), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n3587), .D(N327), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n3587), .D(N326), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n3587), .D(N325), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n3587), .D(N324), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n3587), .D(N323), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n3588), .D(N322), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n3588), .D(N321), .Q(OUT2[0]) );
  AND3_X2 U531 ( .A1(n4170), .A2(ADD_WR[4]), .A3(n1213), .ZN(n1247) );
  AND3_X2 U796 ( .A1(n3923), .A2(n1213), .A3(n265), .ZN(n1352) );
  NOR3_X2 U898 ( .A1(n4173), .A2(n4171), .A3(ADD_WR[1]), .ZN(n1106) );
  NOR3_X2 U932 ( .A1(n4171), .A2(ADD_WR[1]), .A3(ADD_WR[0]), .ZN(n1140) );
  NOR3_X2 U1034 ( .A1(ADD_WR[2]), .A2(n4173), .A3(ADD_WR[1]), .ZN(n1178) );
  AND3_X2 U1036 ( .A1(n3923), .A2(n4170), .A3(n1213), .ZN(n1521) );
  AND2_X2 U1037 ( .A1(WR), .A2(ENABLE), .ZN(n1213) );
  DFFR_X2 \registers_reg[1][18]  ( .D(n3845), .CK(n4212), .RN(n3692), .Q(
        \registers[1][18] ) );
  DFFR_X2 \registers_reg[27][3]  ( .D(n2841), .CK(n4212), .RN(n3615), .QN(n861) );
  DFFR_X2 \registers_reg[27][7]  ( .D(n2845), .CK(n4212), .RN(n3616), .QN(n857) );
  DFFR_X2 \registers_reg[26][3]  ( .D(n2873), .CK(n4212), .RN(n3618), .QN(n829) );
  DFFR_X2 \registers_reg[5][1]  ( .D(n3159), .CK(n4212), .RN(n3679), .QN(n159)
         );
  DFFR_X2 \registers_reg[5][2]  ( .D(n3160), .CK(n4212), .RN(n3679), .QN(n158)
         );
  DFFR_X2 \registers_reg[5][3]  ( .D(n3161), .CK(n4212), .RN(n3679), .QN(n157)
         );
  DFFR_X2 \registers_reg[5][7]  ( .D(n3165), .CK(n4212), .RN(n3680), .QN(n153)
         );
  DFFR_X2 \registers_reg[5][9]  ( .D(n3167), .CK(n4212), .RN(n3680), .QN(n151)
         );
  DFFR_X2 \registers_reg[5][19]  ( .D(n3177), .CK(n4212), .RN(n3681), .QN(n141) );
  DFFR_X2 \registers_reg[5][20]  ( .D(n3178), .CK(n4212), .RN(n3681), .QN(n140) );
  DFFR_X2 \registers_reg[5][21]  ( .D(n3179), .CK(n4212), .RN(n3681), .QN(n139) );
  DFFR_X2 \registers_reg[5][25]  ( .D(n3183), .CK(n4212), .RN(n3681), .QN(n135) );
  DFFR_X2 \registers_reg[5][26]  ( .D(n3184), .CK(n4212), .RN(n3682), .QN(n134) );
  DFFR_X2 \registers_reg[26][2]  ( .D(n2872), .CK(n4212), .RN(n3618), .QN(n830) );
  DFFR_X2 \registers_reg[26][9]  ( .D(n2879), .CK(n4212), .RN(n3619), .QN(n823) );
  DFFR_X2 \registers_reg[26][23]  ( .D(n2893), .CK(n4212), .RN(n3620), .QN(
        n809) );
  DFFR_X2 \registers_reg[26][25]  ( .D(n2895), .CK(n4212), .RN(n3620), .QN(
        n807) );
  DFFR_X2 \registers_reg[26][27]  ( .D(n2897), .CK(n4212), .RN(n3621), .QN(
        n805) );
  DFFR_X2 \registers_reg[10][1]  ( .D(n3127), .CK(n4212), .RN(n3665), .QN(n319) );
  DFFR_X2 \registers_reg[10][3]  ( .D(n3129), .CK(n4212), .RN(n3665), .QN(n317) );
  DFFR_X2 \registers_reg[10][7]  ( .D(n3133), .CK(n4212), .RN(n3665), .QN(n313) );
  DFFR_X2 \registers_reg[10][9]  ( .D(n3135), .CK(n4212), .RN(n3665), .QN(n311) );
  DFFR_X2 \registers_reg[10][19]  ( .D(n3145), .CK(n4212), .RN(n3666), .QN(
        n301) );
  DFFR_X2 \registers_reg[10][20]  ( .D(n3146), .CK(n4212), .RN(n3666), .QN(
        n300) );
  DFFR_X2 \registers_reg[10][21]  ( .D(n3147), .CK(n4212), .RN(n3667), .QN(
        n299) );
  DFFR_X2 \registers_reg[10][25]  ( .D(n3151), .CK(n4212), .RN(n3667), .QN(
        n295) );
  DFFR_X2 \registers_reg[10][26]  ( .D(n3152), .CK(n4212), .RN(n3667), .QN(
        n294) );
  DFFR_X2 \registers_reg[2][1]  ( .D(n3255), .CK(n4212), .RN(n3688), .QN(n63)
         );
  DFFR_X2 \registers_reg[2][2]  ( .D(n3256), .CK(n4212), .RN(n3688), .QN(n62)
         );
  DFFR_X2 \registers_reg[2][3]  ( .D(n3257), .CK(n4212), .RN(n3688), .QN(n61)
         );
  DFFR_X2 \registers_reg[2][7]  ( .D(n3261), .CK(n4212), .RN(n3689), .QN(n57)
         );
  DFFR_X2 \registers_reg[2][9]  ( .D(n3263), .CK(n4212), .RN(n3689), .QN(n55)
         );
  DFFR_X2 \registers_reg[2][19]  ( .D(n3273), .CK(n4212), .RN(n3690), .QN(n45)
         );
  DFFR_X2 \registers_reg[2][20]  ( .D(n3274), .CK(n4212), .RN(n3690), .QN(n44)
         );
  DFFR_X2 \registers_reg[2][25]  ( .D(n3279), .CK(n4212), .RN(n3690), .QN(n39)
         );
  DFFR_X2 \registers_reg[2][26]  ( .D(n3280), .CK(n4212), .RN(n3690), .QN(n38)
         );
  DFFR_X1 \registers_reg[26][17]  ( .D(n2887), .CK(n4212), .RN(n3620), .QN(
        n815) );
  DFFR_X1 \registers_reg[26][16]  ( .D(n2886), .CK(n4212), .RN(n3620), .QN(
        n816) );
  DFFR_X1 \registers_reg[26][8]  ( .D(n2878), .CK(n4212), .RN(n3619), .QN(n824) );
  DFFR_X1 \registers_reg[2][17]  ( .D(n3271), .CK(n4212), .RN(n3689), .QN(n47)
         );
  DFFR_X1 \registers_reg[2][16]  ( .D(n3270), .CK(n4212), .RN(n3689), .QN(n48)
         );
  DFFR_X1 \registers_reg[2][13]  ( .D(n3267), .CK(n4212), .RN(n3689), .QN(n51)
         );
  DFFR_X1 \registers_reg[26][13]  ( .D(n2883), .CK(n4212), .RN(n3619), .QN(
        n819) );
  DFFR_X1 \registers_reg[26][18]  ( .D(n2888), .CK(n4212), .RN(n3620), .QN(
        n814) );
  DFFR_X1 \registers_reg[26][14]  ( .D(n2884), .CK(n4212), .RN(n3619), .QN(
        n818) );
  DFFR_X1 \registers_reg[26][12]  ( .D(n2882), .CK(n4212), .RN(n3619), .QN(
        n820) );
  DFFR_X1 \registers_reg[2][14]  ( .D(n3268), .CK(n4212), .RN(n3689), .QN(n50)
         );
  DFFR_X1 \registers_reg[26][0]  ( .D(n2870), .CK(n4212), .RN(n3618), .QN(n832) );
  DFFR_X1 \registers_reg[2][18]  ( .D(n3272), .CK(n4212), .RN(n3690), .QN(n46)
         );
  DFFR_X1 \registers_reg[2][15]  ( .D(n3269), .CK(n4212), .RN(n3689), .QN(n49)
         );
  DFFR_X1 \registers_reg[2][12]  ( .D(n3266), .CK(n4212), .RN(n3689), .QN(n52)
         );
  DFFR_X1 \registers_reg[26][19]  ( .D(n2889), .CK(n4212), .RN(n3620), .QN(
        n813) );
  DFFR_X1 \registers_reg[26][22]  ( .D(n2892), .CK(n4212), .RN(n3620), .QN(
        n810) );
  DFFR_X1 \registers_reg[5][14]  ( .D(n3172), .CK(n4212), .RN(n3680), .QN(n146) );
  DFFR_X1 \registers_reg[5][13]  ( .D(n3171), .CK(n4212), .RN(n3680), .QN(n147) );
  DFFR_X1 \registers_reg[26][11]  ( .D(n2881), .CK(n4212), .RN(n3619), .QN(
        n821) );
  DFFR_X1 \registers_reg[31][8]  ( .D(n2782), .CK(n4212), .RN(n3604), .QN(n984) );
  DFFR_X1 \registers_reg[31][7]  ( .D(n2781), .CK(n4212), .RN(n3604), .QN(n985) );
  DFFR_X1 \registers_reg[31][0]  ( .D(n2774), .CK(n4212), .RN(n3604), .QN(n992) );
  DFFR_X1 \registers_reg[26][10]  ( .D(n2880), .CK(n4212), .RN(n3619), .QN(
        n822) );
  DFFR_X1 \registers_reg[26][5]  ( .D(n2875), .CK(n4212), .RN(n3619), .QN(n827) );
  DFFR_X1 \registers_reg[11][0]  ( .D(n3094), .CK(n4212), .RN(n3662), .QN(n352) );
  DFFR_X1 \registers_reg[3][0]  ( .D(n3222), .CK(n4212), .RN(n3685), .QN(n96)
         );
  DFFR_X1 \registers_reg[26][1]  ( .D(n2871), .CK(n4212), .RN(n3618), .QN(n831) );
  DFFR_X1 \registers_reg[14][0]  ( .D(n3062), .CK(n4212), .RN(n3653), .QN(n448) );
  DFFR_X1 \registers_reg[30][22]  ( .D(n2828), .CK(n4212), .RN(n3608), .QN(
        n938) );
  DFFR_X1 \registers_reg[30][7]  ( .D(n2813), .CK(n4212), .RN(n3607), .QN(n953) );
  DFFR_X1 \registers_reg[30][5]  ( .D(n2811), .CK(n4212), .RN(n3607), .QN(n955) );
  DFFR_X1 \registers_reg[5][6]  ( .D(n3164), .CK(n4212), .RN(n3680), .QN(n154)
         );
  DFFR_X1 \registers_reg[5][18]  ( .D(n3176), .CK(n4212), .RN(n3681), .QN(n142) );
  DFFR_X1 \registers_reg[5][17]  ( .D(n3175), .CK(n4212), .RN(n3681), .QN(n143) );
  DFFR_X1 \registers_reg[5][16]  ( .D(n3174), .CK(n4212), .RN(n3681), .QN(n144) );
  DFFR_X1 \registers_reg[5][15]  ( .D(n3173), .CK(n4212), .RN(n3681), .QN(n145) );
  DFFR_X1 \registers_reg[5][12]  ( .D(n3170), .CK(n4212), .RN(n3680), .QN(n148) );
  DFFR_X1 \registers_reg[31][1]  ( .D(n2775), .CK(n4212), .RN(n3604), .QN(n991) );
  DFFR_X1 \registers_reg[31][5]  ( .D(n2779), .CK(n4212), .RN(n3604), .QN(n987) );
  DFFR_X1 \registers_reg[30][18]  ( .D(n2824), .CK(n4212), .RN(n3608), .QN(
        n942) );
  DFFR_X1 \registers_reg[30][14]  ( .D(n2820), .CK(n4212), .RN(n3608), .QN(
        n946) );
  DFFR_X1 \registers_reg[14][18]  ( .D(n3080), .CK(n4212), .RN(n3655), .QN(
        n430) );
  DFFR_X1 \registers_reg[14][14]  ( .D(n3076), .CK(n4212), .RN(n3654), .QN(
        n434) );
  DFFR_X1 \registers_reg[11][14]  ( .D(n3108), .CK(n4212), .RN(n3663), .QN(
        n338) );
  DFFR_X1 \registers_reg[4][18]  ( .D(n3208), .CK(n4212), .RN(n3684), .QN(n110) );
  DFFR_X1 \registers_reg[4][14]  ( .D(n3204), .CK(n4212), .RN(n3683), .QN(n114) );
  DFFR_X1 \registers_reg[4][22]  ( .D(n3212), .CK(n4212), .RN(n3684), .QN(n106) );
  DFFR_X1 \registers_reg[4][15]  ( .D(n3205), .CK(n4212), .RN(n3683), .QN(n113) );
  DFFR_X1 \registers_reg[4][12]  ( .D(n3202), .CK(n4212), .RN(n3683), .QN(n116) );
  DFFR_X1 \registers_reg[4][10]  ( .D(n3200), .CK(n4212), .RN(n3683), .QN(n118) );
  DFFR_X1 \registers_reg[4][1]  ( .D(n3191), .CK(n4212), .RN(n3682), .QN(n127)
         );
  DFFR_X1 \registers_reg[4][0]  ( .D(n3190), .CK(n4212), .RN(n3682), .QN(n128)
         );
  DFFR_X1 \registers_reg[31][22]  ( .D(n2796), .CK(n4212), .RN(n3606), .QN(
        n970) );
  DFFR_X1 \registers_reg[31][19]  ( .D(n2793), .CK(n4212), .RN(n3605), .QN(
        n973) );
  DFFR_X1 \registers_reg[31][18]  ( .D(n2792), .CK(n4212), .RN(n3605), .QN(
        n974) );
  DFFR_X1 \registers_reg[31][17]  ( .D(n2791), .CK(n4212), .RN(n3605), .QN(
        n975) );
  DFFR_X1 \registers_reg[31][16]  ( .D(n2790), .CK(n4212), .RN(n3605), .QN(
        n976) );
  DFFR_X1 \registers_reg[31][15]  ( .D(n2789), .CK(n4212), .RN(n3605), .QN(
        n977) );
  DFFR_X1 \registers_reg[31][14]  ( .D(n2788), .CK(n4212), .RN(n3605), .QN(
        n978) );
  DFFR_X1 \registers_reg[31][13]  ( .D(n2787), .CK(n4212), .RN(n3605), .QN(
        n979) );
  DFFR_X1 \registers_reg[31][12]  ( .D(n2786), .CK(n4212), .RN(n3605), .QN(
        n980) );
  DFFR_X1 \registers_reg[31][11]  ( .D(n2785), .CK(n4212), .RN(n3605), .QN(
        n981) );
  DFFR_X1 \registers_reg[31][10]  ( .D(n2784), .CK(n4212), .RN(n3604), .QN(
        n982) );
  DFFR_X1 \registers_reg[31][6]  ( .D(n2780), .CK(n4212), .RN(n3604), .QN(n986) );
  DFFR_X1 \registers_reg[5][22]  ( .D(n3180), .CK(n4212), .RN(n3681), .QN(n138) );
  DFFR_X1 \registers_reg[2][22]  ( .D(n3276), .CK(n4212), .RN(n3690), .QN(n42)
         );
  DFFR_X1 \registers_reg[4][11]  ( .D(n3201), .CK(n4212), .RN(n3683), .QN(n117) );
  DFFR_X1 \registers_reg[5][5]  ( .D(n3163), .CK(n4212), .RN(n3680), .QN(n155)
         );
  DFFR_X1 \registers_reg[14][22]  ( .D(n3084), .CK(n4212), .RN(n3655), .QN(
        n426) );
  DFFR_X1 \registers_reg[30][17]  ( .D(n2823), .CK(n4212), .RN(n3608), .QN(
        n943) );
  DFFR_X1 \registers_reg[4][17]  ( .D(n3207), .CK(n4212), .RN(n3684), .QN(n111) );
  DFFR_X1 \registers_reg[30][19]  ( .D(n2825), .CK(n4212), .RN(n3608), .QN(
        n941) );
  DFFR_X1 \registers_reg[30][15]  ( .D(n2821), .CK(n4212), .RN(n3608), .QN(
        n945) );
  DFFR_X1 \registers_reg[30][10]  ( .D(n2816), .CK(n4212), .RN(n3607), .QN(
        n950) );
  DFFR_X1 \registers_reg[30][8]  ( .D(n2814), .CK(n4212), .RN(n3607), .QN(n952) );
  DFFR_X1 \registers_reg[30][1]  ( .D(n2807), .CK(n4212), .RN(n3607), .QN(n959) );
  DFFR_X1 \registers_reg[14][17]  ( .D(n3079), .CK(n4212), .RN(n3655), .QN(
        n431) );
  DFFR_X1 \registers_reg[14][15]  ( .D(n3077), .CK(n4212), .RN(n3654), .QN(
        n433) );
  DFFR_X1 \registers_reg[14][12]  ( .D(n3074), .CK(n4212), .RN(n3654), .QN(
        n436) );
  DFFR_X1 \registers_reg[14][11]  ( .D(n3073), .CK(n4212), .RN(n3654), .QN(
        n437) );
  DFFR_X1 \registers_reg[14][10]  ( .D(n3072), .CK(n4212), .RN(n3654), .QN(
        n438) );
  DFFR_X1 \registers_reg[5][11]  ( .D(n3169), .CK(n4212), .RN(n3680), .QN(n149) );
  DFFR_X1 \registers_reg[26][30]  ( .D(n2900), .CK(n4212), .RN(n3621), .QN(
        n802) );
  DFFR_X1 \registers_reg[30][30]  ( .D(n2836), .CK(n4212), .RN(n3609), .QN(
        n930) );
  DFFR_X1 \registers_reg[10][30]  ( .D(n3156), .CK(n4212), .RN(n3667), .QN(
        n290) );
  DFFR_X2 \registers_reg[20][5]  ( .D(n2939), .CK(n4212), .RN(n3636), .QN(n635) );
  DFFR_X2 \registers_reg[20][6]  ( .D(n2940), .CK(n4212), .RN(n3636), .QN(n634) );
  DFFR_X2 \registers_reg[21][1]  ( .D(n2903), .CK(n4212), .RN(n3633), .QN(n671) );
  DFFR_X2 \registers_reg[21][2]  ( .D(n2904), .CK(n4212), .RN(n3633), .QN(n670) );
  DFFR_X2 \registers_reg[21][3]  ( .D(n2905), .CK(n4212), .RN(n3633), .QN(n669) );
  DFFR_X2 \registers_reg[21][7]  ( .D(n2909), .CK(n4212), .RN(n3633), .QN(n665) );
  DFFR_X2 \registers_reg[21][9]  ( .D(n2911), .CK(n4212), .RN(n3633), .QN(n663) );
  DFFR_X2 \registers_reg[21][10]  ( .D(n2912), .CK(n4212), .RN(n3634), .QN(
        n662) );
  DFFR_X2 \registers_reg[21][11]  ( .D(n2913), .CK(n4212), .RN(n3634), .QN(
        n661) );
  DFFR_X2 \registers_reg[21][12]  ( .D(n2914), .CK(n4212), .RN(n3634), .QN(
        n660) );
  DFFR_X2 \registers_reg[21][15]  ( .D(n2917), .CK(n4212), .RN(n3634), .QN(
        n657) );
  DFFR_X2 \registers_reg[21][16]  ( .D(n2918), .CK(n4212), .RN(n3634), .QN(
        n656) );
  DFFR_X2 \registers_reg[21][17]  ( .D(n2919), .CK(n4212), .RN(n3634), .QN(
        n655) );
  DFFR_X2 \registers_reg[21][18]  ( .D(n2920), .CK(n4212), .RN(n3634), .QN(
        n654) );
  DFFR_X2 \registers_reg[21][19]  ( .D(n2921), .CK(n4212), .RN(n3634), .QN(
        n653) );
  DFFR_X2 \registers_reg[21][20]  ( .D(n2922), .CK(n4212), .RN(n3634), .QN(
        n652) );
  DFFR_X2 \registers_reg[21][21]  ( .D(n2923), .CK(n4212), .RN(n3635), .QN(
        n651) );
  DFFR_X2 \registers_reg[21][22]  ( .D(n2924), .CK(n4212), .RN(n3635), .QN(
        n650) );
  DFFR_X2 \registers_reg[21][25]  ( .D(n2927), .CK(n4212), .RN(n3635), .QN(
        n647) );
  DFFR_X2 \registers_reg[21][26]  ( .D(n2928), .CK(n4212), .RN(n3635), .QN(
        n646) );
  DFFR_X2 \registers_reg[21][28]  ( .D(n2930), .CK(n4212), .RN(n3635), .QN(
        n644) );
  DFFR_X2 \registers_reg[15][2]  ( .D(n3032), .CK(n4212), .RN(n3650), .QN(n478) );
  DFFR_X2 \registers_reg[15][3]  ( .D(n3033), .CK(n4212), .RN(n3650), .QN(n477) );
  DFFR_X2 \registers_reg[15][6]  ( .D(n3036), .CK(n4212), .RN(n3651), .QN(n474) );
  DFFR_X2 \registers_reg[15][7]  ( .D(n3037), .CK(n4212), .RN(n3651), .QN(n473) );
  DFFR_X2 \registers_reg[15][8]  ( .D(n3038), .CK(n4212), .RN(n3651), .QN(n472) );
  DFFR_X2 \registers_reg[15][9]  ( .D(n3039), .CK(n4212), .RN(n3651), .QN(n471) );
  DFFR_X2 \registers_reg[15][13]  ( .D(n3043), .CK(n4212), .RN(n3651), .QN(
        n467) );
  DFFR_X2 \registers_reg[15][14]  ( .D(n3044), .CK(n4212), .RN(n3651), .QN(
        n466) );
  DFFR_X2 \registers_reg[15][15]  ( .D(n3045), .CK(n4212), .RN(n3651), .QN(
        n465) );
  DFFR_X2 \registers_reg[15][16]  ( .D(n3046), .CK(n4212), .RN(n3652), .QN(
        n464) );
  DFFR_X2 \registers_reg[15][17]  ( .D(n3047), .CK(n4212), .RN(n3652), .QN(
        n463) );
  DFFR_X2 \registers_reg[15][19]  ( .D(n3049), .CK(n4212), .RN(n3652), .QN(
        n461) );
  DFFR_X2 \registers_reg[15][20]  ( .D(n3050), .CK(n4212), .RN(n3652), .QN(
        n460) );
  DFFR_X2 \registers_reg[15][21]  ( .D(n3051), .CK(n4212), .RN(n3652), .QN(
        n459) );
  DFFR_X2 \registers_reg[15][23]  ( .D(n3053), .CK(n4212), .RN(n3652), .QN(
        n457) );
  DFFR_X2 \registers_reg[15][27]  ( .D(n3057), .CK(n4212), .RN(n3653), .QN(
        n453) );
  DFFR_X2 \registers_reg[15][29]  ( .D(n3059), .CK(n4212), .RN(n3653), .QN(
        n451) );
  DFFR_X2 \registers_reg[16][13]  ( .D(n3011), .CK(n4212), .RN(n3648), .QN(
        n499) );
  DFFR_X2 \registers_reg[16][30]  ( .D(n3028), .CK(n4212), .RN(n3650), .QN(
        n482) );
  DFFR_X2 \registers_reg[16][1]  ( .D(n2999), .CK(n4212), .RN(n3647), .QN(n511) );
  DFFR_X2 \registers_reg[16][4]  ( .D(n3002), .CK(n4212), .RN(n3648), .QN(n508) );
  DFFR_X2 \registers_reg[16][8]  ( .D(n3006), .CK(n4212), .RN(n3648), .QN(n504) );
  DFFR_X2 \registers_reg[16][22]  ( .D(n3020), .CK(n4212), .RN(n3649), .QN(
        n490) );
  DFFR_X1 \registers_reg[11][2]  ( .D(n3096), .CK(n4212), .RN(n3662), .QN(n350) );
  DFFR_X2 \registers_reg[17][0]  ( .D(n2966), .CK(n4212), .RN(n3644), .QN(n544) );
  DFFR_X2 \registers_reg[17][3]  ( .D(n2969), .CK(n4212), .RN(n3645), .QN(n541) );
  DFFR_X2 \registers_reg[17][12]  ( .D(n2978), .CK(n4212), .RN(n3645), .QN(
        n532) );
  DFFR_X2 \registers_reg[17][19]  ( .D(n2985), .CK(n4212), .RN(n3646), .QN(
        n525) );
  DFFR_X2 \registers_reg[17][30]  ( .D(n2996), .CK(n4212), .RN(n3647), .QN(
        n514) );
  DFFR_X2 \registers_reg[17][1]  ( .D(n2967), .CK(n4212), .RN(n3644), .QN(n543) );
  DFFR_X2 \registers_reg[17][9]  ( .D(n2975), .CK(n4212), .RN(n3645), .QN(n535) );
  DFFR_X2 \registers_reg[17][16]  ( .D(n2982), .CK(n4212), .RN(n3646), .QN(
        n528) );
  DFFR_X2 \registers_reg[17][21]  ( .D(n2987), .CK(n4212), .RN(n3646), .QN(
        n523) );
  DFFR_X2 \registers_reg[17][22]  ( .D(n2988), .CK(n4212), .RN(n3646), .QN(
        n522) );
  DFFR_X2 \registers_reg[17][29]  ( .D(n2995), .CK(n4212), .RN(n3647), .QN(
        n515) );
  DFFR_X2 \registers_reg[17][2]  ( .D(n2968), .CK(n4212), .RN(n3644), .QN(n542) );
  DFFR_X2 \registers_reg[17][4]  ( .D(n2970), .CK(n4212), .RN(n3645), .QN(n540) );
  DFFR_X2 \registers_reg[17][7]  ( .D(n2973), .CK(n4212), .RN(n3645), .QN(n537) );
  DFFR_X2 \registers_reg[17][8]  ( .D(n2974), .CK(n4212), .RN(n3645), .QN(n536) );
  DFFR_X2 \registers_reg[17][11]  ( .D(n2977), .CK(n4212), .RN(n3645), .QN(
        n533) );
  DFFR_X2 \registers_reg[17][14]  ( .D(n2980), .CK(n4212), .RN(n3646), .QN(
        n530) );
  DFFR_X2 \registers_reg[17][15]  ( .D(n2981), .CK(n4212), .RN(n3646), .QN(
        n529) );
  DFFR_X2 \registers_reg[17][23]  ( .D(n2989), .CK(n4212), .RN(n3646), .QN(
        n521) );
  DFFR_X2 \registers_reg[17][25]  ( .D(n2991), .CK(n4212), .RN(n3647), .QN(
        n519) );
  DFFR_X2 \registers_reg[17][27]  ( .D(n2993), .CK(n4212), .RN(n3647), .QN(
        n517) );
  DFFR_X2 \registers_reg[17][28]  ( .D(n2994), .CK(n4212), .RN(n3647), .QN(
        n516) );
  DFFR_X1 \registers_reg[11][19]  ( .D(n3113), .CK(n4212), .RN(n3663), .QN(
        n333) );
  DFFR_X2 \registers_reg[17][6]  ( .D(n2972), .CK(n4212), .RN(n3645), .QN(n538) );
  DFFR_X2 \registers_reg[17][13]  ( .D(n2979), .CK(n4212), .RN(n3645), .QN(
        n531) );
  DFFR_X2 \registers_reg[17][18]  ( .D(n2984), .CK(n4212), .RN(n3646), .QN(
        n526) );
  DFFR_X2 \registers_reg[17][26]  ( .D(n2992), .CK(n4212), .RN(n3647), .QN(
        n518) );
  DFFR_X2 \registers_reg[17][5]  ( .D(n2971), .CK(n4212), .RN(n3645), .QN(n539) );
  DFFR_X2 \registers_reg[17][17]  ( .D(n2983), .CK(n4212), .RN(n3646), .QN(
        n527) );
  DFFR_X2 \registers_reg[17][20]  ( .D(n2986), .CK(n4212), .RN(n3646), .QN(
        n524) );
  DFFR_X2 \registers_reg[17][31]  ( .D(n2997), .CK(n4212), .RN(n3647), .QN(
        n513) );
  DFFR_X1 \registers_reg[5][28]  ( .D(n3186), .CK(n4212), .RN(n3682), .QN(n132) );
  DFFR_X1 \registers_reg[2][28]  ( .D(n3282), .CK(n4212), .RN(n3690), .QN(n36)
         );
  DFFR_X1 \registers_reg[15][24]  ( .D(n3054), .CK(n4212), .RN(n3652), .QN(
        n456) );
  DFFR_X1 \registers_reg[2][21]  ( .D(n3275), .CK(n4212), .RN(n3690), .QN(n43)
         );
  DFFR_X1 \registers_reg[26][21]  ( .D(n2891), .CK(n4212), .RN(n3620), .QN(
        n811) );
  DFFR_X1 \registers_reg[11][21]  ( .D(n3115), .CK(n4212), .RN(n3664), .QN(
        n331) );
  DFFR_X1 \registers_reg[11][17]  ( .D(n3111), .CK(n4212), .RN(n3663), .QN(
        n335) );
  DFFR_X1 \registers_reg[11][20]  ( .D(n3114), .CK(n4212), .RN(n3664), .QN(
        n332) );
  DFFR_X1 \registers_reg[11][15]  ( .D(n3109), .CK(n4212), .RN(n3663), .QN(
        n337) );
  DFFR_X1 \registers_reg[11][26]  ( .D(n3120), .CK(n4212), .RN(n3664), .QN(
        n326) );
  DFFR_X1 \registers_reg[11][9]  ( .D(n3103), .CK(n4212), .RN(n3663), .QN(n343) );
  DFFR_X1 \registers_reg[11][18]  ( .D(n3112), .CK(n4212), .RN(n3663), .QN(
        n334) );
  DFFR_X1 \registers_reg[11][3]  ( .D(n3097), .CK(n4212), .RN(n3662), .QN(n349) );
  DFFR_X1 \registers_reg[11][10]  ( .D(n3104), .CK(n4212), .RN(n3663), .QN(
        n342) );
  DFFR_X1 \registers_reg[11][1]  ( .D(n3095), .CK(n4212), .RN(n3662), .QN(n351) );
  DFFR_X1 \registers_reg[11][25]  ( .D(n3119), .CK(n4212), .RN(n3664), .QN(
        n327) );
  DFFR_X1 \registers_reg[11][28]  ( .D(n3122), .CK(n4212), .RN(n3664), .QN(
        n324) );
  DFFR_X1 \registers_reg[3][18]  ( .D(n3240), .CK(n4212), .RN(n3687), .QN(n78)
         );
  DFFR_X1 \registers_reg[3][25]  ( .D(n3247), .CK(n4212), .RN(n3687), .QN(n71)
         );
  DFFR_X1 \registers_reg[3][17]  ( .D(n3239), .CK(n4212), .RN(n3687), .QN(n79)
         );
  DFFR_X1 \registers_reg[3][26]  ( .D(n3248), .CK(n4212), .RN(n3687), .QN(n70)
         );
  DFFR_X1 \registers_reg[3][1]  ( .D(n3223), .CK(n4212), .RN(n3685), .QN(n95)
         );
  DFFR_X1 \registers_reg[3][10]  ( .D(n3232), .CK(n4212), .RN(n3686), .QN(n86)
         );
  DFFR_X1 \registers_reg[3][9]  ( .D(n3231), .CK(n4212), .RN(n3686), .QN(n87)
         );
  DFFR_X1 \registers_reg[3][7]  ( .D(n3229), .CK(n4212), .RN(n3686), .QN(n89)
         );
  DFFR_X1 \registers_reg[3][3]  ( .D(n3225), .CK(n4212), .RN(n3685), .QN(n93)
         );
  DFFR_X1 \registers_reg[3][20]  ( .D(n3242), .CK(n4212), .RN(n3687), .QN(n76)
         );
  DFFR_X1 \registers_reg[11][11]  ( .D(n3105), .CK(n4212), .RN(n3663), .QN(
        n341) );
  DFFR_X1 \registers_reg[3][11]  ( .D(n3233), .CK(n4212), .RN(n3686), .QN(n85)
         );
  DFFR_X1 \registers_reg[17][24]  ( .D(n2990), .CK(n4212), .RN(n3646), .QN(
        n520) );
  DFFR_X1 \registers_reg[11][22]  ( .D(n3116), .CK(n4212), .RN(n3664), .QN(
        n330) );
  DFFR_X1 \registers_reg[3][12]  ( .D(n3234), .CK(n4212), .RN(n3686), .QN(n84)
         );
  DFFR_X2 \registers_reg[13][8]  ( .D(n3804), .CK(n4212), .RN(n3657), .Q(
        \registers[13][8] ) );
  DFFR_X2 \registers_reg[13][21]  ( .D(n3816), .CK(n4212), .RN(n3658), .Q(
        \registers[13][21] ) );
  DFFR_X1 \registers_reg[17][10]  ( .D(n2976), .CK(n4212), .RN(n3645), .QN(
        n534) );
  DFFR_X1 \registers_reg[5][10]  ( .D(n3168), .CK(n4212), .RN(n3680), .QN(n150) );
  DFFR_X2 \registers_reg[20][7]  ( .D(n2941), .CK(n4212), .RN(n3636), .QN(n633) );
  DFFR_X2 \registers_reg[20][8]  ( .D(n2942), .CK(n4212), .RN(n3636), .QN(n632) );
  DFFR_X2 \registers_reg[20][9]  ( .D(n2943), .CK(n4212), .RN(n3636), .QN(n631) );
  DFFR_X2 \registers_reg[29][20]  ( .D(n4158), .CK(n4212), .RN(n3611), .Q(
        \registers[29][20] ) );
  DFFR_X2 \registers_reg[29][26]  ( .D(n4164), .CK(n4212), .RN(n3612), .Q(
        \registers[29][26] ) );
  DFFR_X2 \registers_reg[22][1]  ( .D(n234), .CK(n4212), .RN(n3630), .Q(
        \registers[22][1] ), .QN(n235) );
  DFFR_X2 \registers_reg[22][5]  ( .D(n213), .CK(n4212), .RN(n3630), .Q(
        \registers[22][5] ), .QN(n214) );
  DFFR_X2 \registers_reg[22][9]  ( .D(n389), .CK(n4212), .RN(n3631), .Q(
        \registers[22][9] ), .QN(n390) );
  DFFR_X2 \registers_reg[22][17]  ( .D(n200), .CK(n4212), .RN(n3631), .Q(
        \registers[22][17] ), .QN(n201) );
  DFFR_X2 \registers_reg[29][5]  ( .D(n4143), .CK(n4212), .RN(n3610), .Q(
        \registers[29][5] ) );
  DFFR_X2 \registers_reg[9][17]  ( .D(n3755), .CK(n4212), .RN(n3669), .Q(
        \registers[9][17] ) );
  DFFR_X2 \registers_reg[9][24]  ( .D(n3761), .CK(n4212), .RN(n3670), .Q(
        \registers[9][24] ) );
  DFFR_X2 \registers_reg[9][29]  ( .D(n3766), .CK(n4212), .RN(n3670), .Q(
        \registers[9][29] ) );
  DFFR_X2 \registers_reg[9][1]  ( .D(n218), .CK(n4212), .RN(n3668), .Q(
        \registers[9][1] ), .QN(n219) );
  DFFR_X2 \registers_reg[29][14]  ( .D(n4152), .CK(n4212), .RN(n3611), .Q(
        \registers[29][14] ) );
  DFFR_X2 \registers_reg[29][18]  ( .D(n4156), .CK(n4212), .RN(n3611), .Q(
        \registers[29][18] ) );
  DFFR_X2 \registers_reg[29][13]  ( .D(n4151), .CK(n4212), .RN(n3611), .Q(
        \registers[29][13] ) );
  DFFR_X2 \registers_reg[29][1]  ( .D(n4139), .CK(n4212), .RN(n3609), .Q(
        \registers[29][1] ) );
  DFFR_X2 \registers_reg[29][16]  ( .D(n4154), .CK(n4212), .RN(n3611), .Q(
        \registers[29][16] ) );
  DFFR_X2 \registers_reg[29][12]  ( .D(n4150), .CK(n4212), .RN(n3610), .Q(
        \registers[29][12] ) );
  DFFR_X2 \registers_reg[9][23]  ( .D(n3760), .CK(n4212), .RN(n3670), .Q(
        \registers[9][23] ) );
  DFFR_X2 \registers_reg[9][25]  ( .D(n3762), .CK(n4212), .RN(n3670), .Q(
        \registers[9][25] ) );
  DFFR_X2 \registers_reg[9][28]  ( .D(n3765), .CK(n4212), .RN(n3670), .Q(
        \registers[9][28] ) );
  DFFR_X2 \registers_reg[9][18]  ( .D(n3756), .CK(n4212), .RN(n3669), .Q(
        \registers[9][18] ) );
  DFFR_X2 \registers_reg[29][15]  ( .D(n4153), .CK(n4212), .RN(n3611), .Q(
        \registers[29][15] ) );
  DFFR_X2 \registers_reg[9][26]  ( .D(n3763), .CK(n4212), .RN(n3670), .Q(
        \registers[9][26] ) );
  DFFR_X2 \registers_reg[29][2]  ( .D(n4140), .CK(n4212), .RN(n3610), .Q(
        \registers[29][2] ) );
  DFFR_X2 \registers_reg[29][4]  ( .D(n4142), .CK(n4212), .RN(n3610), .Q(
        \registers[29][4] ) );
  DFFR_X2 \registers_reg[29][6]  ( .D(n4144), .CK(n4212), .RN(n3610), .Q(
        \registers[29][6] ) );
  DFFR_X2 \registers_reg[29][7]  ( .D(n4145), .CK(n4212), .RN(n3610), .Q(
        \registers[29][7] ) );
  DFFR_X2 \registers_reg[29][8]  ( .D(n4146), .CK(n4212), .RN(n3610), .Q(
        \registers[29][8] ) );
  DFFR_X2 \registers_reg[29][9]  ( .D(n4147), .CK(n4212), .RN(n3610), .Q(
        \registers[29][9] ) );
  DFFR_X2 \registers_reg[29][10]  ( .D(n4148), .CK(n4212), .RN(n3610), .Q(
        \registers[29][10] ) );
  DFFR_X2 \registers_reg[29][11]  ( .D(n4149), .CK(n4212), .RN(n3610), .Q(
        \registers[29][11] ) );
  DFFR_X2 \registers_reg[29][17]  ( .D(n4155), .CK(n4212), .RN(n3611), .Q(
        \registers[29][17] ) );
  DFFR_X2 \registers_reg[29][21]  ( .D(n4159), .CK(n4212), .RN(n3611), .Q(
        \registers[29][21] ) );
  DFFR_X2 \registers_reg[29][22]  ( .D(n4160), .CK(n4212), .RN(n3611), .Q(
        \registers[29][22] ) );
  DFFR_X2 \registers_reg[29][23]  ( .D(n4161), .CK(n4212), .RN(n3611), .Q(
        \registers[29][23] ) );
  DFFR_X2 \registers_reg[29][24]  ( .D(n4162), .CK(n4212), .RN(n3612), .Q(
        \registers[29][24] ) );
  DFFR_X2 \registers_reg[29][25]  ( .D(n4163), .CK(n4212), .RN(n3612), .Q(
        \registers[29][25] ) );
  DFFR_X2 \registers_reg[29][27]  ( .D(n4165), .CK(n4212), .RN(n3612), .Q(
        \registers[29][27] ) );
  DFFR_X2 \registers_reg[29][28]  ( .D(n4166), .CK(n4212), .RN(n3612), .Q(
        \registers[29][28] ) );
  DFFR_X2 \registers_reg[29][29]  ( .D(n4167), .CK(n4212), .RN(n3612), .Q(
        \registers[29][29] ) );
  DFFR_X2 \registers_reg[29][31]  ( .D(n4169), .CK(n4212), .RN(n3612), .Q(
        \registers[29][31] ) );
  DFFR_X2 \registers_reg[10][2]  ( .D(n3128), .CK(n4212), .RN(n3665), .QN(n318) );
  DFFR_X2 \registers_reg[10][10]  ( .D(n3136), .CK(n4212), .RN(n3666), .QN(
        n310) );
  DFFR_X2 \registers_reg[10][5]  ( .D(n3131), .CK(n4212), .RN(n3665), .QN(n315) );
  DFFR_X2 \registers_reg[10][0]  ( .D(n3126), .CK(n4212), .RN(n3665), .QN(n320) );
  DFFR_X2 \registers_reg[10][4]  ( .D(n3130), .CK(n4212), .RN(n3665), .QN(n316) );
  DFFR_X2 \registers_reg[10][8]  ( .D(n3134), .CK(n4212), .RN(n3665), .QN(n312) );
  DFFR_X2 \registers_reg[10][23]  ( .D(n3149), .CK(n4212), .RN(n3667), .QN(
        n297) );
  DFFR_X2 \registers_reg[10][24]  ( .D(n3150), .CK(n4212), .RN(n3667), .QN(
        n296) );
  DFFR_X2 \registers_reg[10][27]  ( .D(n3153), .CK(n4212), .RN(n3667), .QN(
        n293) );
  DFFR_X2 \registers_reg[10][29]  ( .D(n3155), .CK(n4212), .RN(n3667), .QN(
        n291) );
  DFFR_X2 \registers_reg[10][28]  ( .D(n3154), .CK(n4212), .RN(n3667), .QN(
        n292) );
  DFFR_X2 \registers_reg[10][6]  ( .D(n3132), .CK(n4212), .RN(n3665), .QN(n314) );
  DFFR_X2 \registers_reg[10][22]  ( .D(n3148), .CK(n4212), .RN(n3667), .QN(
        n298) );
  DFFR_X2 \registers_reg[10][15]  ( .D(n3141), .CK(n4212), .RN(n3666), .QN(
        n305) );
  DFFR_X2 \registers_reg[10][12]  ( .D(n3138), .CK(n4212), .RN(n3666), .QN(
        n308) );
  DFFR_X2 \registers_reg[10][14]  ( .D(n3140), .CK(n4212), .RN(n3666), .QN(
        n306) );
  DFFR_X2 \registers_reg[10][13]  ( .D(n3139), .CK(n4212), .RN(n3666), .QN(
        n307) );
  DFFR_X2 \registers_reg[10][16]  ( .D(n3142), .CK(n4212), .RN(n3666), .QN(
        n304) );
  DFFR_X2 \registers_reg[10][17]  ( .D(n3143), .CK(n4212), .RN(n3666), .QN(
        n303) );
  DFFR_X2 \registers_reg[10][18]  ( .D(n3144), .CK(n4212), .RN(n3666), .QN(
        n302) );
  DFFR_X2 \registers_reg[10][11]  ( .D(n3137), .CK(n4212), .RN(n3666), .QN(
        n309) );
  DFFR_X2 \registers_reg[29][0]  ( .D(n4138), .CK(n4212), .RN(n3609), .Q(
        \registers[29][0] ) );
  DFFR_X2 \registers_reg[29][30]  ( .D(n4168), .CK(n4212), .RN(n3612), .Q(
        \registers[29][30] ) );
  DFFR_X2 \registers_reg[13][4]  ( .D(n3800), .CK(n4212), .RN(n3656), .Q(
        \registers[13][4] ) );
  DFFR_X2 \registers_reg[13][14]  ( .D(n3809), .CK(n4212), .RN(n3657), .Q(
        \registers[13][14] ) );
  DFFR_X2 \registers_reg[18][0]  ( .D(n3924), .CK(n4212), .RN(n3641), .Q(
        \registers[18][0] ) );
  DFFR_X2 \registers_reg[18][1]  ( .D(n3925), .CK(n4212), .RN(n3641), .Q(
        \registers[18][1] ) );
  DFFR_X2 \registers_reg[18][4]  ( .D(n3927), .CK(n4212), .RN(n3642), .Q(
        \registers[18][4] ) );
  DFFR_X2 \registers_reg[18][10]  ( .D(n3933), .CK(n4212), .RN(n3642), .Q(
        \registers[18][10] ) );
  DFFR_X2 \registers_reg[18][12]  ( .D(n3935), .CK(n4212), .RN(n3642), .Q(
        \registers[18][12] ) );
  DFFR_X2 \registers_reg[18][13]  ( .D(n3936), .CK(n4212), .RN(n3643), .Q(
        \registers[18][13] ) );
  DFFR_X2 \registers_reg[18][15]  ( .D(n3938), .CK(n4212), .RN(n3643), .Q(
        \registers[18][15] ) );
  DFFR_X2 \registers_reg[18][17]  ( .D(n3940), .CK(n4212), .RN(n3643), .Q(
        \registers[18][17] ) );
  DFFR_X2 \registers_reg[18][18]  ( .D(n3941), .CK(n4212), .RN(n3643), .Q(
        \registers[18][18] ) );
  DFFR_X2 \registers_reg[18][20]  ( .D(n3943), .CK(n4212), .RN(n3643), .Q(
        \registers[18][20] ) );
  DFFR_X2 \registers_reg[18][21]  ( .D(n3944), .CK(n4212), .RN(n3643), .Q(
        \registers[18][21] ) );
  DFFR_X2 \registers_reg[18][22]  ( .D(n3945), .CK(n4212), .RN(n3643), .Q(
        \registers[18][22] ) );
  DFFR_X2 \registers_reg[18][23]  ( .D(n3946), .CK(n4212), .RN(n3643), .Q(
        \registers[18][23] ) );
  DFFR_X2 \registers_reg[18][24]  ( .D(n3947), .CK(n4212), .RN(n3644), .Q(
        \registers[18][24] ) );
  DFFR_X2 \registers_reg[18][2]  ( .D(n3926), .CK(n4212), .RN(n3642), .Q(
        \registers[18][2] ) );
  DFFR_X2 \registers_reg[28][26]  ( .D(n4132), .CK(n4212), .RN(n3615), .Q(
        \registers[28][26] ) );
  DFFR_X2 \registers_reg[6][17]  ( .D(n3876), .CK(n4212), .RN(n3678), .Q(
        \registers[6][17] ) );
  DFFR_X2 \registers_reg[6][21]  ( .D(n3880), .CK(n4212), .RN(n3678), .Q(
        \registers[6][21] ) );
  DFFR_X2 \registers_reg[6][25]  ( .D(n3884), .CK(n4212), .RN(n3679), .Q(
        \registers[6][25] ) );
  DFFR_X2 \registers_reg[6][28]  ( .D(n3887), .CK(n4212), .RN(n3679), .Q(
        \registers[6][28] ) );
  DFFR_X2 \registers_reg[6][1]  ( .D(n3860), .CK(n4212), .RN(n3676), .Q(
        \registers[6][1] ) );
  DFFR_X2 \registers_reg[6][4]  ( .D(n3863), .CK(n4212), .RN(n3677), .Q(
        \registers[6][4] ) );
  DFFR_X2 \registers_reg[6][5]  ( .D(n3864), .CK(n4212), .RN(n3677), .Q(
        \registers[6][5] ) );
  DFFR_X2 \registers_reg[6][9]  ( .D(n3868), .CK(n4212), .RN(n3677), .Q(
        \registers[6][9] ) );
  DFFR_X2 \registers_reg[6][10]  ( .D(n3869), .CK(n4212), .RN(n3677), .Q(
        \registers[6][10] ) );
  DFFR_X2 \registers_reg[6][12]  ( .D(n3871), .CK(n4212), .RN(n3677), .Q(
        \registers[6][12] ) );
  DFFR_X2 \registers_reg[6][16]  ( .D(n3875), .CK(n4212), .RN(n3678), .Q(
        \registers[6][16] ) );
  DFFR_X2 \registers_reg[6][18]  ( .D(n3877), .CK(n4212), .RN(n3678), .Q(
        \registers[6][18] ) );
  DFFR_X2 \registers_reg[6][30]  ( .D(n3889), .CK(n4212), .RN(n3679), .Q(
        \registers[6][30] ) );
  DFFR_X2 \registers_reg[28][25]  ( .D(n4131), .CK(n4212), .RN(n3615), .Q(
        \registers[28][25] ) );
  DFFR_X2 \registers_reg[24][4]  ( .D(n4047), .CK(n4212), .RN(n3624), .Q(
        \registers[24][4] ) );
  DFFR_X2 \registers_reg[24][31]  ( .D(n4074), .CK(n4212), .RN(n3627), .Q(
        \registers[24][31] ) );
  DFFR_X2 \registers_reg[6][13]  ( .D(n3872), .CK(n4212), .RN(n3677), .Q(
        \registers[6][13] ) );
  DFFR_X2 \registers_reg[28][7]  ( .D(n4113), .CK(n4212), .RN(n3613), .Q(
        \registers[28][7] ) );
  DFFR_X2 \registers_reg[18][5]  ( .D(n3928), .CK(n4212), .RN(n3642), .Q(
        \registers[18][5] ) );
  DFFR_X2 \registers_reg[18][6]  ( .D(n3929), .CK(n4212), .RN(n3642), .Q(
        \registers[18][6] ) );
  DFFR_X2 \registers_reg[18][7]  ( .D(n3930), .CK(n4212), .RN(n3642), .Q(
        \registers[18][7] ) );
  DFFR_X2 \registers_reg[18][8]  ( .D(n3931), .CK(n4212), .RN(n3642), .Q(
        \registers[18][8] ) );
  DFFR_X2 \registers_reg[18][9]  ( .D(n3932), .CK(n4212), .RN(n3642), .Q(
        \registers[18][9] ) );
  DFFR_X2 \registers_reg[18][14]  ( .D(n3937), .CK(n4212), .RN(n3643), .Q(
        \registers[18][14] ) );
  DFFR_X2 \registers_reg[18][16]  ( .D(n3939), .CK(n4212), .RN(n3643), .Q(
        \registers[18][16] ) );
  DFFR_X2 \registers_reg[18][25]  ( .D(n3948), .CK(n4212), .RN(n3644), .Q(
        \registers[18][25] ) );
  DFFR_X2 \registers_reg[18][26]  ( .D(n3949), .CK(n4212), .RN(n3644), .Q(
        \registers[18][26] ) );
  DFFR_X2 \registers_reg[18][27]  ( .D(n3950), .CK(n4212), .RN(n3644), .Q(
        \registers[18][27] ) );
  DFFR_X2 \registers_reg[18][28]  ( .D(n3951), .CK(n4212), .RN(n3644), .Q(
        \registers[18][28] ) );
  DFFR_X2 \registers_reg[18][29]  ( .D(n3952), .CK(n4212), .RN(n3644), .Q(
        \registers[18][29] ) );
  DFFR_X2 \registers_reg[18][11]  ( .D(n3934), .CK(n4212), .RN(n3642), .Q(
        \registers[18][11] ) );
  DFFR_X2 \registers_reg[24][10]  ( .D(n4053), .CK(n4212), .RN(n3625), .Q(
        \registers[24][10] ) );
  DFFR_X2 \registers_reg[24][21]  ( .D(n4064), .CK(n4212), .RN(n3626), .Q(
        \registers[24][21] ) );
  DFFR_X2 \registers_reg[6][0]  ( .D(n3859), .CK(n4212), .RN(n3676), .Q(
        \registers[6][0] ) );
  DFFR_X2 \registers_reg[6][14]  ( .D(n3873), .CK(n4212), .RN(n3678), .Q(
        \registers[6][14] ) );
  DFFR_X2 \registers_reg[6][27]  ( .D(n3886), .CK(n4212), .RN(n3679), .Q(
        \registers[6][27] ) );
  DFFR_X2 \registers_reg[6][31]  ( .D(n3890), .CK(n4212), .RN(n3679), .Q(
        \registers[6][31] ) );
  DFFR_X2 \registers_reg[28][13]  ( .D(n4119), .CK(n4212), .RN(n3613), .Q(
        \registers[28][13] ) );
  DFFR_X2 \registers_reg[28][15]  ( .D(n4121), .CK(n4212), .RN(n3614), .Q(
        \registers[28][15] ) );
  DFFR_X2 \registers_reg[6][23]  ( .D(n3882), .CK(n4212), .RN(n3678), .Q(
        \registers[6][23] ) );
  DFFR_X2 \registers_reg[6][26]  ( .D(n3885), .CK(n4212), .RN(n3679), .Q(
        \registers[6][26] ) );
  DFFR_X2 \registers_reg[6][6]  ( .D(n3865), .CK(n4212), .RN(n3677), .Q(
        \registers[6][6] ) );
  DFFR_X2 \registers_reg[6][20]  ( .D(n3879), .CK(n4212), .RN(n3678), .Q(
        \registers[6][20] ) );
  DFFR_X2 \registers_reg[24][5]  ( .D(n4048), .CK(n4212), .RN(n3624), .Q(
        \registers[24][5] ) );
  DFFR_X2 \registers_reg[26][26]  ( .D(n2896), .CK(n4212), .RN(n3620), .QN(
        n806) );
  DFFR_X2 \registers_reg[26][24]  ( .D(n2894), .CK(n4212), .RN(n3620), .QN(
        n808) );
  DFFR_X2 \registers_reg[26][28]  ( .D(n2898), .CK(n4212), .RN(n3621), .QN(
        n804) );
  DFFR_X2 \registers_reg[26][29]  ( .D(n2899), .CK(n4212), .RN(n3621), .QN(
        n803) );
  DFFR_X2 \registers_reg[26][20]  ( .D(n2890), .CK(n4212), .RN(n3620), .QN(
        n812) );
  DFFR_X2 \registers_reg[26][6]  ( .D(n2876), .CK(n4212), .RN(n3619), .QN(n826) );
  DFFR_X2 \registers_reg[26][7]  ( .D(n2877), .CK(n4212), .RN(RST_AN), .QN(
        n825) );
  DFFR_X2 \registers_reg[24][1]  ( .D(n4044), .CK(n4212), .RN(n3624), .Q(
        \registers[24][1] ) );
  DFFR_X2 \registers_reg[24][7]  ( .D(n4050), .CK(n4212), .RN(n3625), .Q(
        \registers[24][7] ) );
  DFFR_X2 \registers_reg[24][9]  ( .D(n4052), .CK(n4212), .RN(n3625), .Q(
        \registers[24][9] ) );
  DFFR_X2 \registers_reg[24][14]  ( .D(n4057), .CK(n4212), .RN(n3625), .Q(
        \registers[24][14] ) );
  DFFR_X2 \registers_reg[24][22]  ( .D(n4065), .CK(n4212), .RN(n3626), .Q(
        \registers[24][22] ) );
  DFFR_X2 \registers_reg[24][27]  ( .D(n4070), .CK(n4212), .RN(n3626), .Q(
        \registers[24][27] ) );
  DFFR_X2 \registers_reg[6][15]  ( .D(n3874), .CK(n4212), .RN(n3678), .Q(
        \registers[6][15] ) );
  DFFR_X2 \registers_reg[6][11]  ( .D(n3870), .CK(n4212), .RN(n3677), .Q(
        \registers[6][11] ) );
  DFFR_X2 \registers_reg[6][24]  ( .D(n3883), .CK(n4212), .RN(n3678), .Q(
        \registers[6][24] ) );
  DFFR_X2 \registers_reg[6][2]  ( .D(n3861), .CK(n4212), .RN(n3676), .Q(
        \registers[6][2] ) );
  DFFR_X2 \registers_reg[13][2]  ( .D(n404), .CK(n4212), .RN(n3656), .Q(
        \registers[13][2] ) );
  DFFR_X2 \registers_reg[13][12]  ( .D(n394), .CK(n4212), .RN(n3657), .Q(
        \registers[13][12] ) );
  DFFR_X2 \registers_reg[27][13]  ( .D(n2851), .CK(n4212), .RN(n3616), .QN(
        n851) );
  DFFR_X2 \registers_reg[27][14]  ( .D(n2852), .CK(n4212), .RN(n3616), .QN(
        n850) );
  DFFR_X2 \registers_reg[27][15]  ( .D(n2853), .CK(n4212), .RN(n3617), .QN(
        n849) );
  DFFR_X2 \registers_reg[27][19]  ( .D(n2857), .CK(n4212), .RN(n3617), .QN(
        n845) );
  DFFR_X2 \registers_reg[27][23]  ( .D(n2861), .CK(n4212), .RN(n3617), .QN(
        n841) );
  DFFR_X2 \registers_reg[6][29]  ( .D(n3888), .CK(n4212), .RN(n3679), .Q(
        \registers[6][29] ) );
  DFFR_X2 \registers_reg[23][4]  ( .D(n4015), .CK(n4212), .RN(n3627), .Q(
        \registers[23][4] ) );
  DFFR_X2 \registers_reg[23][11]  ( .D(n4022), .CK(n4212), .RN(n3628), .Q(
        \registers[23][11] ) );
  DFFR_X2 \registers_reg[23][13]  ( .D(n4024), .CK(n4212), .RN(n3628), .Q(
        \registers[23][13] ) );
  DFFR_X2 \registers_reg[23][16]  ( .D(n4027), .CK(n4212), .RN(n3628), .Q(
        \registers[23][16] ) );
  DFFR_X2 \registers_reg[23][17]  ( .D(n4028), .CK(n4212), .RN(n3628), .Q(
        \registers[23][17] ) );
  DFFR_X2 \registers_reg[11][7]  ( .D(n3101), .CK(n4212), .RN(n3662), .QN(n345) );
  DFFR_X2 \registers_reg[11][5]  ( .D(n3099), .CK(n4212), .RN(n3662), .QN(n347) );
  DFFR_X2 \registers_reg[11][6]  ( .D(n3100), .CK(n4212), .RN(n3662), .QN(n346) );
  DFFR_X2 \registers_reg[11][8]  ( .D(n3102), .CK(n4212), .RN(n3662), .QN(n344) );
  DFFR_X2 \registers_reg[30][11]  ( .D(n2817), .CK(n4212), .RN(n3607), .QN(
        n949) );
  DFFR_X2 \registers_reg[30][3]  ( .D(n2809), .CK(n4212), .RN(n3607), .QN(n957) );
  DFFR_X2 \registers_reg[30][9]  ( .D(n2815), .CK(n4212), .RN(n3607), .QN(n951) );
  DFFR_X2 \registers_reg[30][12]  ( .D(n2818), .CK(n4212), .RN(n3608), .QN(
        n948) );
  DFFR_X2 \registers_reg[30][24]  ( .D(n2830), .CK(n4212), .RN(n3609), .QN(
        n936) );
  DFFR_X2 \registers_reg[30][25]  ( .D(n2831), .CK(n4212), .RN(n3609), .QN(
        n935) );
  DFFR_X2 \registers_reg[30][27]  ( .D(n2833), .CK(n4212), .RN(n3609), .QN(
        n933) );
  DFFR_X2 \registers_reg[30][29]  ( .D(n2835), .CK(n4212), .RN(n3609), .QN(
        n931) );
  DFFR_X2 \registers_reg[26][15]  ( .D(n2885), .CK(n4212), .RN(n3619), .QN(
        n817) );
  DFFR_X2 \registers_reg[23][22]  ( .D(n4033), .CK(n4212), .RN(n3629), .Q(
        \registers[23][22] ) );
  DFFR_X2 \registers_reg[28][17]  ( .D(n4123), .CK(n4212), .RN(n3614), .Q(
        \registers[28][17] ) );
  DFFR_X2 \registers_reg[28][11]  ( .D(n4117), .CK(n4212), .RN(n3613), .Q(
        \registers[28][11] ) );
  DFFR_X2 \registers_reg[28][21]  ( .D(n4127), .CK(n4212), .RN(n3614), .Q(
        \registers[28][21] ) );
  DFFR_X2 \registers_reg[28][29]  ( .D(n4135), .CK(n4212), .RN(n3615), .Q(
        \registers[28][29] ) );
  DFFR_X2 \registers_reg[14][1]  ( .D(n3063), .CK(n4212), .RN(n3653), .QN(n447) );
  DFFR_X2 \registers_reg[23][27]  ( .D(n4038), .CK(n4212), .RN(n3629), .Q(
        \registers[23][27] ) );
  DFFR_X2 \registers_reg[25][7]  ( .D(n4082), .CK(n4212), .RN(n3622), .Q(
        \registers[25][7] ) );
  DFFR_X2 \registers_reg[13][5]  ( .D(n3801), .CK(n4212), .RN(n3656), .Q(
        \registers[13][5] ) );
  DFFR_X2 \registers_reg[13][10]  ( .D(n3806), .CK(n4212), .RN(n3657), .Q(
        \registers[13][10] ) );
  DFFR_X2 \registers_reg[13][11]  ( .D(n3807), .CK(n4212), .RN(n3657), .Q(
        \registers[13][11] ) );
  DFFR_X2 \registers_reg[13][18]  ( .D(n3813), .CK(n4212), .RN(n3658), .Q(
        \registers[13][18] ) );
  DFFR_X2 \registers_reg[13][22]  ( .D(n3817), .CK(n4212), .RN(n3658), .Q(
        \registers[13][22] ) );
  DFFR_X2 \registers_reg[13][31]  ( .D(n3826), .CK(n4212), .RN(n3659), .Q(
        \registers[13][31] ) );
  DFFR_X2 \registers_reg[21][5]  ( .D(n2907), .CK(n4212), .RN(n3633), .QN(n667) );
  DFFR_X2 \registers_reg[19][12]  ( .D(n3966), .CK(n4212), .RN(n3640), .Q(
        \registers[19][12] ) );
  DFFR_X2 \registers_reg[19][14]  ( .D(n3968), .CK(n4212), .RN(n3640), .Q(
        \registers[19][14] ) );
  DFFR_X2 \registers_reg[2][10]  ( .D(n3264), .CK(n4212), .RN(n3689), .QN(n54)
         );
  DFFR_X2 \registers_reg[2][5]  ( .D(n3259), .CK(n4212), .RN(n3688), .QN(n59)
         );
  DFFR_X2 \registers_reg[2][11]  ( .D(n3265), .CK(n4212), .RN(n3689), .QN(n53)
         );
  DFFR_X2 \registers_reg[2][6]  ( .D(n3260), .CK(n4212), .RN(n3688), .QN(n58)
         );
  DFFR_X2 \registers_reg[2][8]  ( .D(n3262), .CK(n4212), .RN(n3689), .QN(n56)
         );
  DFFR_X2 \registers_reg[28][9]  ( .D(n4115), .CK(n4212), .RN(n3613), .Q(
        \registers[28][9] ) );
  DFFR_X2 \registers_reg[1][6]  ( .D(n3833), .CK(n4212), .RN(n3691), .Q(
        \registers[1][6] ) );
  DFFR_X2 \registers_reg[1][7]  ( .D(n3834), .CK(n4212), .RN(n3691), .Q(
        \registers[1][7] ) );
  DFFR_X2 \registers_reg[1][22]  ( .D(n3849), .CK(n4212), .RN(n3693), .Q(
        \registers[1][22] ) );
  DFFR_X2 \registers_reg[28][14]  ( .D(n4120), .CK(n4212), .RN(n3614), .Q(
        \registers[28][14] ) );
  DFFR_X2 \registers_reg[6][8]  ( .D(n3867), .CK(n4212), .RN(n3677), .Q(
        \registers[6][8] ) );
  DFFR_X2 \registers_reg[6][7]  ( .D(n3866), .CK(n4212), .RN(n3677), .Q(
        \registers[6][7] ) );
  DFFR_X2 \registers_reg[3][2]  ( .D(n3224), .CK(n4212), .RN(n3685), .QN(n94)
         );
  DFFR_X2 \registers_reg[3][15]  ( .D(n3237), .CK(n4212), .RN(n3686), .QN(n81)
         );
  DFFR_X2 \registers_reg[3][28]  ( .D(n3250), .CK(n4212), .RN(n3688), .QN(n68)
         );
  DFFR_X2 \registers_reg[3][16]  ( .D(n3238), .CK(n4212), .RN(n3686), .QN(n80)
         );
  DFFR_X2 \registers_reg[3][22]  ( .D(n3244), .CK(n4212), .RN(n3687), .QN(n74)
         );
  DFFR_X2 \registers_reg[3][19]  ( .D(n3241), .CK(n4212), .RN(n3687), .QN(n77)
         );
  DFFR_X2 \registers_reg[3][21]  ( .D(n3243), .CK(n4212), .RN(n3687), .QN(n75)
         );
  DFFR_X2 \registers_reg[3][14]  ( .D(n3236), .CK(n4212), .RN(n3686), .QN(n82)
         );
  DFFR_X2 \registers_reg[3][29]  ( .D(n3251), .CK(n4212), .RN(n3688), .QN(n67)
         );
  DFFR_X2 \registers_reg[6][3]  ( .D(n3862), .CK(n4212), .RN(n3677), .Q(
        \registers[6][3] ) );
  DFFR_X2 \registers_reg[19][18]  ( .D(n3972), .CK(n4212), .RN(n3640), .Q(
        \registers[19][18] ) );
  DFFR_X2 \registers_reg[19][13]  ( .D(n3967), .CK(n4212), .RN(n3640), .Q(
        \registers[19][13] ) );
  DFFR_X2 \registers_reg[20][1]  ( .D(n2935), .CK(n4212), .RN(n3636), .QN(n639) );
  DFFR_X2 \registers_reg[20][2]  ( .D(n2936), .CK(n4212), .RN(n3636), .QN(n638) );
  DFFR_X2 \registers_reg[20][10]  ( .D(n2944), .CK(n4212), .RN(n3636), .QN(
        n630) );
  DFFR_X2 \registers_reg[20][14]  ( .D(n2948), .CK(n4212), .RN(n3637), .QN(
        n626) );
  DFFR_X2 \registers_reg[20][15]  ( .D(n2949), .CK(n4212), .RN(n3637), .QN(
        n625) );
  DFFR_X2 \registers_reg[20][16]  ( .D(n2950), .CK(n4212), .RN(n3637), .QN(
        n624) );
  DFFR_X2 \registers_reg[20][21]  ( .D(n2955), .CK(n4212), .RN(n3637), .QN(
        n619) );
  DFFR_X2 \registers_reg[20][24]  ( .D(n2958), .CK(n4212), .RN(n3638), .QN(
        n616) );
  DFFR_X2 \registers_reg[20][25]  ( .D(n2959), .CK(n4212), .RN(n3638), .QN(
        n615) );
  DFFR_X2 \registers_reg[20][26]  ( .D(n2960), .CK(n4212), .RN(n3638), .QN(
        n614) );
  DFFR_X2 \registers_reg[1][2]  ( .D(n3829), .CK(n4212), .RN(n3691), .Q(
        \registers[1][2] ) );
  DFFR_X2 \registers_reg[1][8]  ( .D(n3835), .CK(n4212), .RN(n3692), .Q(
        \registers[1][8] ) );
  DFFR_X2 \registers_reg[1][23]  ( .D(n3850), .CK(n4212), .RN(n3693), .Q(
        \registers[1][23] ) );
  DFFR_X2 \registers_reg[1][31]  ( .D(n3858), .CK(n4212), .RN(n3694), .Q(
        \registers[1][31] ) );
  DFFR_X2 \registers_reg[19][25]  ( .D(n3979), .CK(n4212), .RN(n3641), .Q(
        \registers[19][25] ) );
  DFFR_X2 \registers_reg[19][30]  ( .D(n3984), .CK(n4212), .RN(n3641), .Q(
        \registers[19][30] ) );
  DFFR_X2 \registers_reg[24][25]  ( .D(n4068), .CK(n4212), .RN(n3626), .Q(
        \registers[24][25] ) );
  DFFR_X2 \registers_reg[19][6]  ( .D(n3960), .CK(n4212), .RN(n3639), .Q(
        \registers[19][6] ) );
  DFFR_X2 \registers_reg[19][8]  ( .D(n3962), .CK(n4212), .RN(n3639), .Q(
        \registers[19][8] ) );
  DFFR_X2 \registers_reg[19][23]  ( .D(n3977), .CK(n4212), .RN(n3641), .Q(
        \registers[19][23] ) );
  DFFR_X2 \registers_reg[19][29]  ( .D(n3983), .CK(n4212), .RN(n3641), .Q(
        \registers[19][29] ) );
  DFFR_X2 \registers_reg[12][6]  ( .D(n3774), .CK(n4212), .RN(n3659), .Q(
        \registers[12][6] ) );
  DFFR_X2 \registers_reg[12][27]  ( .D(n3792), .CK(n4212), .RN(n3661), .Q(
        \registers[12][27] ) );
  DFFR_X2 \registers_reg[12][28]  ( .D(n3793), .CK(n4212), .RN(n3661), .Q(
        \registers[12][28] ) );
  DFFR_X2 \registers_reg[11][16]  ( .D(n3110), .CK(n4212), .RN(n3663), .QN(
        n336) );
  DFFR_X2 \registers_reg[11][12]  ( .D(n3106), .CK(n4212), .RN(n3663), .QN(
        n340) );
  DFFR_X2 \registers_reg[9][4]  ( .D(n258), .CK(n4212), .RN(n3668), .Q(
        \registers[9][4] ), .QN(n259) );
  DFFR_X2 \registers_reg[9][22]  ( .D(n242), .CK(n4212), .RN(n3670), .Q(
        \registers[9][22] ), .QN(n243) );
  DFFR_X2 \registers_reg[12][0]  ( .D(n266), .CK(n4212), .RN(n3659), .Q(
        \registers[12][0] ), .QN(n267) );
  DFFR_X2 \registers_reg[28][1]  ( .D(n4108), .CK(n4212), .RN(n3612), .Q(
        \registers[28][1] ) );
  BUF_X1 U2 ( .A(n3341), .Z(n1) );
  CLKBUF_X3 U3 ( .A(n208), .Z(n3357) );
  BUF_X1 U4 ( .A(n3488), .Z(n2) );
  BUF_X1 U5 ( .A(n3488), .Z(n3) );
  BUF_X1 U6 ( .A(n3488), .Z(n4) );
  INV_X1 U7 ( .A(n877), .ZN(n5) );
  INV_X1 U8 ( .A(n877), .ZN(n6) );
  INV_X1 U9 ( .A(n877), .ZN(n272) );
  INV_X1 U10 ( .A(n277), .ZN(n7) );
  INV_X1 U11 ( .A(n880), .ZN(n8) );
  INV_X1 U12 ( .A(n880), .ZN(n9) );
  BUF_X1 U13 ( .A(n563), .Z(n3506) );
  INV_X1 U14 ( .A(n237), .ZN(n10) );
  INV_X1 U15 ( .A(n3532), .ZN(n3526) );
  BUF_X1 U16 ( .A(n575), .Z(n3500) );
  BUF_X2 U17 ( .A(n898), .Z(n575) );
  BUF_X1 U18 ( .A(n3501), .Z(n359) );
  BUF_X1 U19 ( .A(n3442), .Z(n11) );
  BUF_X2 U20 ( .A(n3442), .Z(n12) );
  BUF_X1 U21 ( .A(n3442), .Z(n13) );
  BUF_X1 U22 ( .A(n1355), .Z(n3442) );
  BUF_X2 U23 ( .A(n178), .Z(n3545) );
  BUF_X1 U24 ( .A(n3362), .Z(n269) );
  CLKBUF_X3 U25 ( .A(n897), .Z(n563) );
  CLKBUF_X3 U26 ( .A(n897), .Z(n3511) );
  BUF_X1 U27 ( .A(n278), .Z(n14) );
  INV_X1 U28 ( .A(n867), .ZN(n15) );
  INV_X1 U29 ( .A(n867), .ZN(n16) );
  INV_X1 U30 ( .A(n3532), .ZN(n17) );
  INV_X1 U31 ( .A(n3532), .ZN(n3524) );
  BUF_X1 U32 ( .A(n3489), .Z(n18) );
  BUF_X2 U33 ( .A(n3489), .Z(n19) );
  BUF_X1 U34 ( .A(n1284), .Z(n3489) );
  CLKBUF_X3 U35 ( .A(n549), .Z(n3351) );
  BUF_X2 U36 ( .A(DATAIN[25]), .Z(n367) );
  BUF_X1 U37 ( .A(n1388), .Z(n3436) );
  BUF_X1 U38 ( .A(n207), .Z(n270) );
  CLKBUF_X3 U39 ( .A(n902), .Z(n3432) );
  CLKBUF_X2 U40 ( .A(n552), .Z(n3427) );
  BUF_X1 U41 ( .A(n904), .Z(n20) );
  BUF_X1 U42 ( .A(n904), .Z(n21) );
  BUF_X1 U43 ( .A(n21), .Z(n22) );
  AND2_X2 U44 ( .A1(n360), .A2(n1521), .ZN(n904) );
  BUF_X1 U45 ( .A(n600), .Z(n23) );
  BUF_X1 U46 ( .A(n1560), .Z(n3341) );
  INV_X1 U47 ( .A(n884), .ZN(n24) );
  INV_X1 U48 ( .A(n884), .ZN(n25) );
  BUF_X2 U49 ( .A(n1523), .Z(n3386) );
  BUF_X2 U50 ( .A(n1523), .Z(n3385) );
  BUF_X2 U51 ( .A(n1523), .Z(n3388) );
  CLKBUF_X3 U52 ( .A(n549), .Z(n3349) );
  BUF_X1 U53 ( .A(n549), .Z(n3347) );
  BUF_X1 U54 ( .A(n592), .Z(n361) );
  BUF_X1 U55 ( .A(n901), .Z(n3474) );
  CLKBUF_X3 U56 ( .A(n1068), .Z(n3582) );
  CLKBUF_X1 U57 ( .A(n1068), .Z(n3584) );
  CLKBUF_X1 U58 ( .A(n1068), .Z(n3583) );
  BUF_X1 U59 ( .A(n1074), .Z(n692) );
  CLKBUF_X3 U60 ( .A(n1074), .Z(n3572) );
  OAI22_X1 U61 ( .A1(n4211), .A2(n186), .B1(n185), .B2(n27), .ZN(n26) );
  CLKBUF_X1 U62 ( .A(n3512), .Z(n363) );
  CLKBUF_X3 U63 ( .A(n595), .Z(n185) );
  CLKBUF_X1 U64 ( .A(n3576), .Z(n28) );
  CLKBUF_X3 U65 ( .A(n3576), .Z(n29) );
  BUF_X1 U66 ( .A(n411), .Z(n3576) );
  BUF_X2 U67 ( .A(n551), .Z(n3420) );
  BUF_X2 U68 ( .A(n903), .Z(n551) );
  NOR2_X1 U69 ( .A1(n4178), .A2(ADD_RD2[2]), .ZN(n2160) );
  NOR2_X1 U70 ( .A1(n4175), .A2(ADD_RD1[2]), .ZN(n2751) );
  BUF_X2 U71 ( .A(n407), .Z(n3449) );
  BUF_X1 U72 ( .A(n1523), .Z(n3387) );
  BUF_X1 U73 ( .A(n899), .Z(n562) );
  BUF_X1 U74 ( .A(n904), .Z(n3362) );
  BUF_X1 U75 ( .A(DATAIN[8]), .Z(n793) );
  BUF_X2 U76 ( .A(n895), .Z(n3557) );
  BUF_X2 U77 ( .A(n896), .Z(n178) );
  BUF_X1 U78 ( .A(DATAIN[6]), .Z(n227) );
  BUF_X1 U79 ( .A(n1388), .Z(n3438) );
  BUF_X1 U80 ( .A(DATAIN[6]), .Z(n228) );
  INV_X1 U81 ( .A(n3535), .ZN(n31) );
  BUF_X1 U82 ( .A(n1456), .Z(n32) );
  INV_X1 U83 ( .A(n797), .ZN(n678) );
  BUF_X1 U84 ( .A(DATAIN[0]), .Z(n165) );
  BUF_X1 U85 ( .A(DATAIN[0]), .Z(n180) );
  BUF_X1 U86 ( .A(DATAIN[24]), .Z(n871) );
  BUF_X1 U87 ( .A(DATAIN[24]), .Z(n236) );
  INV_X2 U88 ( .A(n1068), .ZN(n3579) );
  BUF_X1 U89 ( .A(n3490), .Z(n161) );
  BUF_X1 U90 ( .A(n3490), .Z(n162) );
  BUF_X1 U91 ( .A(n3490), .Z(n163) );
  OR2_X1 U92 ( .A1(n447), .A2(n3448), .ZN(n405) );
  BUF_X1 U93 ( .A(DATAIN[7]), .Z(n795) );
  CLKBUF_X1 U94 ( .A(n874), .Z(n374) );
  BUF_X1 U95 ( .A(n32), .Z(n189) );
  INV_X1 U96 ( .A(n3523), .ZN(n3519) );
  BUF_X1 U97 ( .A(DATAIN[30]), .Z(n288) );
  BUF_X2 U98 ( .A(n164), .Z(n3346) );
  INV_X1 U99 ( .A(n880), .ZN(n714) );
  BUF_X1 U100 ( .A(DATAIN[4]), .Z(n882) );
  INV_X1 U101 ( .A(n791), .ZN(n192) );
  CLKBUF_X3 U102 ( .A(n553), .Z(n3541) );
  BUF_X2 U103 ( .A(n1180), .Z(n3532) );
  CLKBUF_X3 U104 ( .A(n4188), .Z(n286) );
  BUF_X1 U105 ( .A(n563), .Z(n3508) );
  BUF_X1 U106 ( .A(n563), .Z(n3507) );
  BUF_X1 U107 ( .A(n563), .Z(n3509) );
  CLKBUF_X3 U108 ( .A(n905), .Z(n164) );
  INV_X1 U109 ( .A(n871), .ZN(n166) );
  INV_X1 U110 ( .A(n871), .ZN(n167) );
  INV_X1 U111 ( .A(n871), .ZN(n4187) );
  BUF_X1 U112 ( .A(DATAIN[17]), .Z(n193) );
  CLKBUF_X1 U113 ( .A(DATAIN[17]), .Z(n709) );
  INV_X1 U114 ( .A(DATAIN[11]), .ZN(n168) );
  INV_X1 U115 ( .A(DATAIN[11]), .ZN(n169) );
  INV_X1 U116 ( .A(n880), .ZN(n170) );
  BUF_X1 U117 ( .A(DATAIN[6]), .Z(n880) );
  BUF_X1 U118 ( .A(n575), .Z(n3497) );
  BUF_X1 U119 ( .A(n575), .Z(n3496) );
  BUF_X1 U120 ( .A(n575), .Z(n3498) );
  BUF_X1 U121 ( .A(n575), .Z(n3499) );
  INV_X1 U122 ( .A(n869), .ZN(n171) );
  INV_X1 U123 ( .A(n875), .ZN(n172) );
  INV_X1 U124 ( .A(n3523), .ZN(n173) );
  INV_X1 U125 ( .A(n3523), .ZN(n3517) );
  BUF_X1 U126 ( .A(DATAIN[21]), .Z(n237) );
  CLKBUF_X3 U127 ( .A(n4186), .Z(n283) );
  INV_X1 U128 ( .A(n867), .ZN(n683) );
  BUF_X1 U129 ( .A(DATAIN[28]), .Z(n867) );
  BUF_X1 U130 ( .A(n207), .Z(n174) );
  BUF_X1 U131 ( .A(n550), .Z(n175) );
  CLKBUF_X3 U132 ( .A(n4207), .Z(n356) );
  INV_X1 U133 ( .A(n884), .ZN(n271) );
  BUF_X1 U134 ( .A(DATAIN[27]), .Z(n884) );
  INV_X1 U135 ( .A(n3422), .ZN(n176) );
  INV_X1 U136 ( .A(n237), .ZN(n257) );
  INV_X1 U137 ( .A(n237), .ZN(n744) );
  INV_X1 U138 ( .A(DATAIN[31]), .ZN(n713) );
  BUF_X1 U139 ( .A(DATAIN[31]), .Z(n877) );
  BUF_X1 U140 ( .A(n895), .Z(n177) );
  BUF_X2 U141 ( .A(n573), .Z(n3556) );
  BUF_X2 U142 ( .A(n3547), .Z(n3543) );
  INV_X1 U143 ( .A(n871), .ZN(n686) );
  BUF_X1 U144 ( .A(n3474), .Z(n205) );
  BUF_X1 U145 ( .A(n3472), .Z(n179) );
  CLKBUF_X1 U146 ( .A(n901), .Z(n3472) );
  INV_X1 U147 ( .A(n791), .ZN(n677) );
  INV_X1 U148 ( .A(n227), .ZN(n4205) );
  BUF_X1 U149 ( .A(n3437), .Z(n277) );
  BUF_X1 U150 ( .A(n553), .Z(n3542) );
  BUF_X1 U151 ( .A(n553), .Z(n3546) );
  BUF_X2 U152 ( .A(DATAIN[22]), .Z(n874) );
  INV_X1 U153 ( .A(n867), .ZN(n682) );
  INV_X1 U154 ( .A(n867), .ZN(n4183) );
  BUF_X2 U155 ( .A(n3352), .Z(n3350) );
  INV_X1 U156 ( .A(n884), .ZN(n716) );
  BUF_X1 U157 ( .A(n3435), .Z(n181) );
  BUF_X1 U158 ( .A(n1456), .Z(n3407) );
  BUF_X2 U159 ( .A(n1317), .Z(n3484) );
  CLKBUF_X3 U160 ( .A(n407), .Z(n225) );
  CLKBUF_X3 U161 ( .A(n407), .Z(n226) );
  BUF_X1 U162 ( .A(n3560), .Z(n182) );
  BUF_X1 U163 ( .A(n1180), .Z(n3527) );
  BUF_X1 U164 ( .A(n551), .Z(n3416) );
  BUF_X1 U165 ( .A(n551), .Z(n3418) );
  BUF_X1 U166 ( .A(n551), .Z(n3421) );
  BUF_X1 U167 ( .A(n551), .Z(n3419) );
  BUF_X1 U168 ( .A(n1215), .Z(n3521) );
  BUF_X1 U169 ( .A(n1215), .Z(n3520) );
  BUF_X1 U170 ( .A(n1215), .Z(n3522) );
  INV_X1 U171 ( .A(n3532), .ZN(n3525) );
  BUF_X1 U172 ( .A(n3341), .Z(n264) );
  BUF_X1 U173 ( .A(n595), .Z(n183) );
  BUF_X2 U174 ( .A(n595), .Z(n184) );
  INV_X1 U175 ( .A(n183), .ZN(n186) );
  BUF_X1 U176 ( .A(n756), .Z(n595) );
  BUF_X1 U177 ( .A(DATAIN[3]), .Z(n799) );
  INV_X1 U178 ( .A(n891), .ZN(n187) );
  INV_X1 U179 ( .A(n891), .ZN(n188) );
  BUF_X1 U180 ( .A(n1247), .Z(n548) );
  BUF_X1 U181 ( .A(DATAIN[30]), .Z(n190) );
  BUF_X1 U182 ( .A(DATAIN[30]), .Z(n866) );
  BUF_X1 U183 ( .A(DATAIN[13]), .Z(n191) );
  CLKBUF_X1 U184 ( .A(DATAIN[13]), .Z(n705) );
  BUF_X1 U185 ( .A(n1423), .Z(n3412) );
  BUF_X1 U186 ( .A(n901), .Z(n3475) );
  BUF_X1 U187 ( .A(n901), .Z(n3476) );
  BUF_X1 U188 ( .A(n901), .Z(n3471) );
  BUF_X1 U189 ( .A(n901), .Z(n3470) );
  BUF_X1 U190 ( .A(n901), .Z(n3473) );
  BUF_X1 U191 ( .A(n3512), .Z(n194) );
  INV_X1 U192 ( .A(n3386), .ZN(n195) );
  INV_X1 U193 ( .A(n3388), .ZN(n196) );
  INV_X1 U194 ( .A(n3572), .ZN(n197) );
  BUF_X1 U195 ( .A(DATAIN[7]), .Z(n198) );
  BUF_X1 U196 ( .A(DATAIN[7]), .Z(n199) );
  BUF_X1 U197 ( .A(DATAIN[7]), .Z(n796) );
  CLKBUF_X1 U198 ( .A(n1317), .Z(n3480) );
  CLKBUF_X1 U199 ( .A(n1317), .Z(n3482) );
  OAI22_X1 U200 ( .A1(n773), .A2(n221), .B1(n185), .B2(n201), .ZN(n200) );
  INV_X1 U201 ( .A(n18), .ZN(n202) );
  BUF_X1 U202 ( .A(DATAIN[8]), .Z(n203) );
  BUF_X1 U203 ( .A(DATAIN[8]), .Z(n204) );
  BUF_X1 U204 ( .A(DATAIN[8]), .Z(n794) );
  BUF_X1 U205 ( .A(n709), .Z(n206) );
  BUF_X1 U206 ( .A(n902), .Z(n207) );
  BUF_X1 U207 ( .A(n904), .Z(n208) );
  OAI22_X1 U208 ( .A1(n776), .A2(n3434), .B1(n222), .B2(n210), .ZN(n209) );
  BUF_X2 U209 ( .A(n1284), .Z(n3491) );
  BUF_X1 U210 ( .A(n1249), .Z(n211) );
  INV_X1 U211 ( .A(n3342), .ZN(n380) );
  INV_X1 U212 ( .A(n3342), .ZN(n3338) );
  BUF_X1 U213 ( .A(n3471), .Z(n212) );
  OAI22_X1 U214 ( .A1(n679), .A2(n221), .B1(n184), .B2(n214), .ZN(n213) );
  INV_X1 U215 ( .A(n797), .ZN(n4206) );
  NAND2_X1 U216 ( .A1(n1521), .A2(n1069), .ZN(n215) );
  NAND2_X1 U217 ( .A1(n1521), .A2(n1069), .ZN(n1489) );
  INV_X1 U218 ( .A(n3434), .ZN(n216) );
  INV_X1 U219 ( .A(n3434), .ZN(n217) );
  OAI22_X1 U220 ( .A1(n694), .A2(n385), .B1(n561), .B2(n219), .ZN(n218) );
  BUF_X1 U221 ( .A(n3437), .Z(n220) );
  BUF_X1 U222 ( .A(DATAIN[16]), .Z(n711) );
  INV_X1 U223 ( .A(n183), .ZN(n221) );
  INV_X1 U224 ( .A(n181), .ZN(n222) );
  CLKBUF_X3 U225 ( .A(n4202), .Z(n370) );
  CLKBUF_X3 U226 ( .A(n4202), .Z(n369) );
  BUF_X1 U227 ( .A(n3476), .Z(n223) );
  BUF_X1 U228 ( .A(n3474), .Z(n224) );
  BUF_X1 U229 ( .A(n3341), .Z(n263) );
  BUF_X1 U230 ( .A(n3560), .Z(n229) );
  BUF_X1 U231 ( .A(n3560), .Z(n230) );
  BUF_X1 U232 ( .A(n3560), .Z(n231) );
  BUF_X1 U233 ( .A(n1108), .Z(n3560) );
  BUF_X1 U234 ( .A(n1249), .Z(n3514) );
  OAI22_X1 U235 ( .A1(n6), .A2(n221), .B1(n185), .B2(n233), .ZN(n232) );
  BUF_X1 U236 ( .A(n4182), .Z(n376) );
  CLKBUF_X3 U237 ( .A(n563), .Z(n3505) );
  BUF_X1 U238 ( .A(n4182), .Z(n377) );
  BUF_X1 U239 ( .A(n563), .Z(n3510) );
  BUF_X1 U240 ( .A(n1388), .Z(n3435) );
  OAI22_X1 U241 ( .A1(n4210), .A2(n186), .B1(n185), .B2(n235), .ZN(n234) );
  INV_X1 U242 ( .A(n891), .ZN(n694) );
  CLKBUF_X1 U243 ( .A(ADD_WR[3]), .Z(n265) );
  INV_X1 U244 ( .A(n869), .ZN(n4185) );
  INV_X1 U245 ( .A(n869), .ZN(n684) );
  INV_X1 U246 ( .A(n869), .ZN(n685) );
  INV_X1 U247 ( .A(n875), .ZN(n4191) );
  INV_X1 U248 ( .A(n875), .ZN(n687) );
  INV_X1 U249 ( .A(n875), .ZN(n688) );
  INV_X1 U250 ( .A(n3577), .ZN(n238) );
  INV_X1 U251 ( .A(n238), .ZN(n239) );
  INV_X1 U252 ( .A(n238), .ZN(n240) );
  INV_X1 U253 ( .A(n238), .ZN(n241) );
  OAI22_X1 U254 ( .A1(n608), .A2(n381), .B1(n244), .B2(n243), .ZN(n242) );
  INV_X1 U255 ( .A(n354), .ZN(n244) );
  OAI22_X1 U256 ( .A1(n368), .A2(n385), .B1(n384), .B2(n246), .ZN(n245) );
  BUF_X2 U257 ( .A(DATAIN[9]), .Z(n589) );
  INV_X1 U258 ( .A(n865), .ZN(n247) );
  INV_X1 U259 ( .A(n795), .ZN(n248) );
  INV_X1 U260 ( .A(n795), .ZN(n249) );
  INV_X1 U261 ( .A(n795), .ZN(n690) );
  CLKBUF_X3 U262 ( .A(n1388), .Z(n3434) );
  BUF_X2 U263 ( .A(DATAIN[28]), .Z(n250) );
  BUF_X2 U264 ( .A(DATAIN[27]), .Z(n251) );
  BUF_X1 U265 ( .A(n3362), .Z(n3356) );
  BUF_X1 U266 ( .A(n21), .Z(n3358) );
  BUF_X1 U267 ( .A(n208), .Z(n3360) );
  BUF_X1 U268 ( .A(n550), .Z(n3361) );
  BUF_X1 U269 ( .A(n20), .Z(n3359) );
  BUF_X1 U270 ( .A(n207), .Z(n3426) );
  BUF_X1 U271 ( .A(n552), .Z(n3428) );
  BUF_X1 U272 ( .A(n207), .Z(n3430) );
  BUF_X1 U273 ( .A(n3432), .Z(n3431) );
  BUF_X1 U274 ( .A(n207), .Z(n3429) );
  BUF_X2 U275 ( .A(DATAIN[31]), .Z(n252) );
  INV_X1 U276 ( .A(n3445), .ZN(n3439) );
  INV_X1 U277 ( .A(n793), .ZN(n253) );
  INV_X1 U278 ( .A(n793), .ZN(n254) );
  INV_X1 U279 ( .A(n793), .ZN(n689) );
  BUF_X1 U280 ( .A(n3341), .Z(n262) );
  OAI22_X1 U281 ( .A1(n715), .A2(n385), .B1(n256), .B2(n382), .ZN(n255) );
  INV_X1 U282 ( .A(n880), .ZN(n715) );
  OAI22_X1 U283 ( .A1(n355), .A2(n3410), .B1(n244), .B2(n259), .ZN(n258) );
  OAI22_X1 U284 ( .A1(n767), .A2(n385), .B1(n384), .B2(n261), .ZN(n260) );
  OAI22_X1 U285 ( .A1(n14), .A2(n4211), .B1(n222), .B2(n267), .ZN(n266) );
  BUF_X1 U286 ( .A(n894), .Z(n268) );
  INV_X1 U287 ( .A(n865), .ZN(n681) );
  INV_X1 U288 ( .A(n3464), .ZN(n273) );
  BUF_X1 U289 ( .A(n3435), .Z(n274) );
  BUF_X1 U290 ( .A(n3435), .Z(n275) );
  BUF_X1 U291 ( .A(n3435), .Z(n276) );
  BUF_X1 U292 ( .A(n3437), .Z(n278) );
  BUF_X1 U293 ( .A(n585), .Z(n3530) );
  BUF_X1 U294 ( .A(n585), .Z(n3531) );
  INV_X1 U295 ( .A(n799), .ZN(n279) );
  INV_X1 U296 ( .A(n799), .ZN(n280) );
  INV_X1 U297 ( .A(n799), .ZN(n691) );
  BUF_X1 U298 ( .A(n692), .Z(n554) );
  BUF_X1 U299 ( .A(n692), .Z(n3567) );
  BUF_X1 U300 ( .A(n692), .Z(n3569) );
  BUF_X1 U301 ( .A(n692), .Z(n3570) );
  BUF_X1 U302 ( .A(n692), .Z(n3571) );
  CLKBUF_X1 U303 ( .A(n3511), .Z(n281) );
  CLKBUF_X1 U304 ( .A(n4186), .Z(n282) );
  CLKBUF_X1 U305 ( .A(n4186), .Z(n284) );
  INV_X1 U306 ( .A(DATAIN[25]), .ZN(n4186) );
  BUF_X1 U307 ( .A(n600), .Z(n3401) );
  BUF_X1 U308 ( .A(n32), .Z(n3402) );
  BUF_X1 U309 ( .A(n600), .Z(n3404) );
  BUF_X1 U310 ( .A(n3407), .Z(n3405) );
  BUF_X1 U311 ( .A(n600), .Z(n3406) );
  BUF_X1 U312 ( .A(n600), .Z(n3403) );
  CLKBUF_X1 U313 ( .A(n4188), .Z(n285) );
  CLKBUF_X1 U314 ( .A(n4188), .Z(n287) );
  INV_X1 U315 ( .A(DATAIN[23]), .ZN(n4188) );
  BUF_X2 U316 ( .A(n893), .Z(n353) );
  INV_X1 U317 ( .A(n865), .ZN(n680) );
  BUF_X2 U318 ( .A(n1146), .Z(n386) );
  BUF_X2 U319 ( .A(n1146), .Z(n3537) );
  INV_X1 U320 ( .A(n757), .ZN(n721) );
  INV_X1 U321 ( .A(n865), .ZN(n4181) );
  BUF_X1 U322 ( .A(n1423), .Z(n354) );
  CLKBUF_X1 U323 ( .A(n4207), .Z(n355) );
  CLKBUF_X1 U324 ( .A(n4207), .Z(n357) );
  INV_X1 U325 ( .A(DATAIN[4]), .ZN(n4207) );
  INV_X1 U326 ( .A(n215), .ZN(n358) );
  BUF_X1 U327 ( .A(n1142), .Z(n360) );
  NOR3_X1 U328 ( .A1(n4172), .A2(n4173), .A3(ADD_WR[2]), .ZN(n1142) );
  BUF_X1 U329 ( .A(n592), .Z(n3516) );
  INV_X1 U330 ( .A(n1249), .ZN(n3513) );
  BUF_X1 U331 ( .A(n1249), .Z(n387) );
  BUF_X1 U332 ( .A(n3512), .Z(n362) );
  BUF_X1 U333 ( .A(n3512), .Z(n364) );
  BUF_X1 U334 ( .A(DATAIN[15]), .Z(n780) );
  BUF_X1 U335 ( .A(DATAIN[14]), .Z(n783) );
  BUF_X1 U336 ( .A(DATAIN[12]), .Z(n788) );
  INV_X1 U337 ( .A(n3342), .ZN(n365) );
  INV_X1 U338 ( .A(n3342), .ZN(n366) );
  INV_X1 U339 ( .A(n3342), .ZN(n3337) );
  CLKBUF_X1 U340 ( .A(n4202), .Z(n368) );
  INV_X1 U341 ( .A(DATAIN[9]), .ZN(n4202) );
  BUF_X2 U342 ( .A(DATAIN[23]), .Z(n371) );
  INV_X1 U343 ( .A(n3458), .ZN(n372) );
  BUF_X1 U344 ( .A(n874), .Z(n373) );
  BUF_X1 U345 ( .A(n575), .Z(n3495) );
  BUF_X2 U346 ( .A(DATAIN[2]), .Z(n375) );
  BUF_X2 U347 ( .A(n4182), .Z(n378) );
  INV_X1 U348 ( .A(DATAIN[29]), .ZN(n4182) );
  BUF_X1 U349 ( .A(n1144), .Z(n379) );
  NOR3_X1 U350 ( .A1(n4172), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n1144) );
  BUF_X1 U351 ( .A(DATAIN[18]), .Z(n771) );
  INV_X1 U352 ( .A(n3342), .ZN(n3339) );
  BUF_X1 U353 ( .A(n1423), .Z(n381) );
  INV_X1 U354 ( .A(n721), .ZN(n382) );
  BUF_X1 U355 ( .A(n585), .Z(n3529) );
  INV_X1 U356 ( .A(n3467), .ZN(n383) );
  INV_X1 U357 ( .A(n721), .ZN(n384) );
  INV_X1 U358 ( .A(n757), .ZN(n385) );
  BUF_X2 U359 ( .A(n1146), .Z(n3535) );
  INV_X1 U360 ( .A(n1249), .ZN(n388) );
  OAI22_X1 U361 ( .A1(n369), .A2(n186), .B1(n184), .B2(n390), .ZN(n389) );
  INV_X1 U362 ( .A(n3445), .ZN(n391) );
  INV_X1 U363 ( .A(n3445), .ZN(n3441) );
  NAND2_X1 U364 ( .A1(n718), .A2(n708), .ZN(n392) );
  NAND2_X1 U365 ( .A1(n3444), .A2(\registers[13][12] ), .ZN(n393) );
  NAND2_X1 U366 ( .A1(n392), .A2(n393), .ZN(n394) );
  INV_X1 U367 ( .A(n3563), .ZN(n395) );
  INV_X1 U368 ( .A(n3491), .ZN(n396) );
  BUF_X2 U369 ( .A(DATAIN[29]), .Z(n397) );
  INV_X1 U370 ( .A(n3387), .ZN(n398) );
  INV_X2 U371 ( .A(n215), .ZN(n3390) );
  NAND2_X1 U372 ( .A1(n400), .A2(n401), .ZN(n399) );
  NAND2_X1 U373 ( .A1(n702), .A2(n695), .ZN(n400) );
  NAND2_X1 U374 ( .A1(n277), .A2(\registers[12][15] ), .ZN(n401) );
  NAND2_X1 U375 ( .A1(n717), .A2(n890), .ZN(n402) );
  NAND2_X1 U376 ( .A1(n3444), .A2(\registers[13][2] ), .ZN(n403) );
  NAND2_X1 U377 ( .A1(n402), .A2(n403), .ZN(n404) );
  INV_X1 U378 ( .A(n3445), .ZN(n3440) );
  NAND2_X1 U379 ( .A1(n405), .A2(n406), .ZN(n3063) );
  AND2_X1 U380 ( .A1(n1072), .A2(n1352), .ZN(n407) );
  NAND2_X1 U381 ( .A1(n3448), .A2(n891), .ZN(n406) );
  CLKBUF_X3 U382 ( .A(n407), .Z(n3448) );
  BUF_X2 U383 ( .A(DATAIN[1]), .Z(n891) );
  INV_X1 U384 ( .A(n891), .ZN(n4210) );
  NAND2_X1 U385 ( .A1(n408), .A2(n409), .ZN(n2806) );
  INV_X1 U386 ( .A(n28), .ZN(n410) );
  NAND2_X1 U387 ( .A1(n30), .A2(n410), .ZN(n408) );
  AND2_X1 U388 ( .A1(n1072), .A2(n1070), .ZN(n411) );
  NAND2_X1 U389 ( .A1(n3578), .A2(n180), .ZN(n409) );
  BUF_X1 U390 ( .A(n411), .Z(n3577) );
  INV_X1 U391 ( .A(n3474), .ZN(n412) );
  OAI22_X1 U392 ( .A1(n168), .A2(n220), .B1(n7), .B2(n414), .ZN(n413) );
  CLKBUF_X1 U393 ( .A(n1388), .Z(n3437) );
  OAI22_X1 U394 ( .A1(n691), .A2(n387), .B1(n184), .B2(n416), .ZN(n415) );
  INV_X1 U395 ( .A(n3563), .ZN(n545) );
  INV_X1 U396 ( .A(n3491), .ZN(n546) );
  INV_X1 U397 ( .A(n3387), .ZN(n547) );
  BUF_X1 U398 ( .A(n905), .Z(n549) );
  BUF_X1 U399 ( .A(n904), .Z(n550) );
  BUF_X1 U400 ( .A(n902), .Z(n552) );
  BUF_X1 U401 ( .A(n896), .Z(n553) );
  BUF_X2 U402 ( .A(n1146), .Z(n3536) );
  BUF_X1 U403 ( .A(n692), .Z(n3568) );
  INV_X1 U404 ( .A(n3471), .ZN(n555) );
  INV_X1 U405 ( .A(n3472), .ZN(n556) );
  INV_X1 U406 ( .A(n3563), .ZN(n3559) );
  BUF_X1 U407 ( .A(n585), .Z(n557) );
  BUF_X1 U408 ( .A(n585), .Z(n3528) );
  INV_X1 U409 ( .A(n3449), .ZN(n558) );
  INV_X1 U410 ( .A(n3449), .ZN(n559) );
  INV_X1 U411 ( .A(n3578), .ZN(n560) );
  BUF_X2 U412 ( .A(n1215), .Z(n3523) );
  INV_X1 U413 ( .A(n721), .ZN(n561) );
  INV_X1 U414 ( .A(n721), .ZN(n3409) );
  INV_X1 U415 ( .A(n3352), .ZN(n564) );
  INV_X1 U416 ( .A(n164), .ZN(n565) );
  INV_X1 U417 ( .A(n3362), .ZN(n566) );
  INV_X1 U418 ( .A(n20), .ZN(n567) );
  INV_X1 U419 ( .A(n3422), .ZN(n568) );
  INV_X1 U420 ( .A(n3422), .ZN(n569) );
  INV_X1 U421 ( .A(n3432), .ZN(n570) );
  INV_X1 U422 ( .A(n552), .ZN(n571) );
  INV_X1 U423 ( .A(n178), .ZN(n572) );
  BUF_X1 U424 ( .A(n895), .Z(n573) );
  INV_X1 U425 ( .A(n721), .ZN(n3408) );
  BUF_X2 U426 ( .A(n900), .Z(n574) );
  INV_X1 U427 ( .A(n891), .ZN(n693) );
  CLKBUF_X3 U428 ( .A(n411), .Z(n3578) );
  INV_X1 U429 ( .A(n3387), .ZN(n576) );
  BUF_X1 U430 ( .A(n1284), .Z(n3488) );
  BUF_X1 U431 ( .A(n1284), .Z(n3490) );
  INV_X1 U432 ( .A(n3511), .ZN(n577) );
  INV_X1 U433 ( .A(n3371), .ZN(n578) );
  INV_X1 U434 ( .A(n3501), .ZN(n579) );
  OAI22_X1 U435 ( .A1(n691), .A2(n3481), .B1(n3479), .B2(n581), .ZN(n580) );
  CLKBUF_X1 U436 ( .A(n1317), .Z(n3481) );
  OAI22_X1 U437 ( .A1(n693), .A2(n3), .B1(n202), .B2(n583), .ZN(n582) );
  BUF_X1 U438 ( .A(n1423), .Z(n3410) );
  BUF_X1 U439 ( .A(n1423), .Z(n3411) );
  INV_X1 U440 ( .A(n3434), .ZN(n584) );
  BUF_X1 U441 ( .A(n1180), .Z(n585) );
  BUF_X1 U442 ( .A(n709), .Z(n774) );
  BUF_X1 U443 ( .A(n874), .Z(n586) );
  BUF_X1 U444 ( .A(n874), .Z(n587) );
  BUF_X1 U445 ( .A(n874), .Z(n588) );
  BUF_X2 U446 ( .A(DATAIN[4]), .Z(n590) );
  INV_X1 U447 ( .A(n3537), .ZN(n591) );
  INV_X1 U448 ( .A(n756), .ZN(n592) );
  NOR3_X1 U449 ( .A1(n4172), .A2(ADD_WR[0]), .A3(n768), .ZN(n1072) );
  BUF_X1 U450 ( .A(n592), .Z(n3515) );
  INV_X1 U451 ( .A(n3458), .ZN(n593) );
  INV_X1 U452 ( .A(n3458), .ZN(n594) );
  CLKBUF_X3 U453 ( .A(n893), .Z(n3458) );
  INV_X1 U454 ( .A(n3484), .ZN(n596) );
  INV_X1 U455 ( .A(n18), .ZN(n597) );
  INV_X1 U456 ( .A(n3387), .ZN(n598) );
  INV_X1 U457 ( .A(n3387), .ZN(n599) );
  BUF_X1 U458 ( .A(DATAIN[18]), .Z(n699) );
  BUF_X1 U459 ( .A(DATAIN[14]), .Z(n703) );
  BUF_X1 U460 ( .A(n1355), .Z(n3444) );
  BUF_X2 U461 ( .A(n1560), .Z(n3340) );
  BUF_X1 U462 ( .A(n1456), .Z(n600) );
  OAI22_X1 U463 ( .A1(n679), .A2(n3561), .B1(n753), .B2(n602), .ZN(n601) );
  INV_X1 U464 ( .A(n797), .ZN(n679) );
  INV_X1 U465 ( .A(n3563), .ZN(n3558) );
  INV_X1 U466 ( .A(n3532), .ZN(n603) );
  INV_X1 U467 ( .A(n3532), .ZN(n604) );
  INV_X1 U468 ( .A(n3467), .ZN(n605) );
  INV_X1 U469 ( .A(n3467), .ZN(n606) );
  CLKBUF_X3 U470 ( .A(n894), .Z(n3467) );
  CLKBUF_X1 U471 ( .A(n353), .Z(n3452) );
  CLKBUF_X1 U472 ( .A(n353), .Z(n3453) );
  CLKBUF_X1 U473 ( .A(n353), .Z(n3454) );
  CLKBUF_X1 U474 ( .A(n353), .Z(n3455) );
  CLKBUF_X1 U475 ( .A(n353), .Z(n3456) );
  CLKBUF_X1 U476 ( .A(n353), .Z(n3457) );
  INV_X1 U477 ( .A(n873), .ZN(n607) );
  INV_X1 U478 ( .A(n873), .ZN(n608) );
  INV_X1 U479 ( .A(n873), .ZN(n4189) );
  INV_X1 U480 ( .A(n3578), .ZN(n673) );
  INV_X1 U481 ( .A(n3578), .ZN(n674) );
  INV_X1 U482 ( .A(n32), .ZN(n675) );
  INV_X1 U483 ( .A(n3407), .ZN(n676) );
  INV_X1 U484 ( .A(n791), .ZN(n4192) );
  BUF_X1 U485 ( .A(n711), .Z(n777) );
  INV_X1 U486 ( .A(n793), .ZN(n4203) );
  INV_X1 U487 ( .A(n795), .ZN(n4204) );
  INV_X1 U488 ( .A(n799), .ZN(n4208) );
  BUF_X1 U489 ( .A(DATAIN[15]), .Z(n701) );
  BUF_X1 U490 ( .A(DATAIN[12]), .Z(n707) );
  NOR3_X1 U491 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(ADD_WR[1]), .ZN(n1212) );
  BUF_X2 U492 ( .A(DATAIN[23]), .Z(n887) );
  INV_X1 U493 ( .A(n3438), .ZN(n695) );
  INV_X1 U494 ( .A(n3438), .ZN(n696) );
  INV_X1 U495 ( .A(n3438), .ZN(n3433) );
  INV_X1 U496 ( .A(n3449), .ZN(n697) );
  INV_X1 U497 ( .A(n3449), .ZN(n698) );
  BUF_X2 U498 ( .A(DATAIN[18]), .Z(n700) );
  BUF_X2 U499 ( .A(DATAIN[15]), .Z(n702) );
  BUF_X2 U500 ( .A(DATAIN[14]), .Z(n704) );
  BUF_X2 U501 ( .A(DATAIN[13]), .Z(n706) );
  BUF_X2 U502 ( .A(DATAIN[12]), .Z(n708) );
  BUF_X2 U503 ( .A(DATAIN[17]), .Z(n710) );
  BUF_X2 U504 ( .A(DATAIN[16]), .Z(n712) );
  INV_X1 U505 ( .A(n877), .ZN(n4180) );
  INV_X1 U506 ( .A(n884), .ZN(n4184) );
  INV_X1 U507 ( .A(n3445), .ZN(n717) );
  INV_X1 U508 ( .A(n3445), .ZN(n718) );
  BUF_X2 U509 ( .A(n1355), .Z(n3445) );
  INV_X1 U510 ( .A(n3537), .ZN(n719) );
  INV_X1 U511 ( .A(n3535), .ZN(n720) );
  INV_X1 U512 ( .A(n757), .ZN(n1423) );
  AND3_X1 U513 ( .A1(ADD_WR[3]), .A2(ADD_WR[4]), .A3(n1213), .ZN(n1070) );
  CLKBUF_X1 U514 ( .A(n215), .Z(n3397) );
  INV_X1 U515 ( .A(n3476), .ZN(n722) );
  INV_X1 U516 ( .A(n3472), .ZN(n723) );
  INV_X1 U517 ( .A(n3491), .ZN(n724) );
  INV_X1 U518 ( .A(n3491), .ZN(n725) );
  INV_X1 U519 ( .A(n552), .ZN(n726) );
  INV_X1 U520 ( .A(n3557), .ZN(n727) );
  INV_X1 U521 ( .A(n3557), .ZN(n728) );
  INV_X1 U522 ( .A(n3484), .ZN(n729) );
  INV_X1 U523 ( .A(n3484), .ZN(n730) );
  INV_X1 U524 ( .A(n3547), .ZN(n731) );
  INV_X1 U525 ( .A(n178), .ZN(n732) );
  CLKBUF_X3 U526 ( .A(n896), .Z(n3547) );
  INV_X1 U527 ( .A(n3371), .ZN(n733) );
  INV_X1 U528 ( .A(n3371), .ZN(n734) );
  CLKBUF_X3 U529 ( .A(n900), .Z(n3371) );
  INV_X1 U530 ( .A(n3501), .ZN(n735) );
  CLKBUF_X3 U532 ( .A(n898), .Z(n3501) );
  INV_X1 U533 ( .A(n3381), .ZN(n736) );
  INV_X1 U534 ( .A(n3381), .ZN(n737) );
  CLKBUF_X3 U535 ( .A(n899), .Z(n3381) );
  INV_X1 U536 ( .A(n3511), .ZN(n738) );
  INV_X1 U537 ( .A(n208), .ZN(n739) );
  INV_X1 U538 ( .A(n164), .ZN(n740) );
  INV_X1 U539 ( .A(n3352), .ZN(n741) );
  CLKBUF_X3 U540 ( .A(n905), .Z(n3352) );
  INV_X1 U541 ( .A(n3422), .ZN(n742) );
  INV_X1 U542 ( .A(n3422), .ZN(n743) );
  CLKBUF_X3 U543 ( .A(n903), .Z(n3422) );
  INV_X1 U544 ( .A(n237), .ZN(n4190) );
  BUF_X1 U545 ( .A(DATAIN[19]), .Z(n791) );
  BUF_X1 U546 ( .A(n1108), .Z(n3561) );
  INV_X1 U547 ( .A(n3572), .ZN(n745) );
  INV_X1 U548 ( .A(n3572), .ZN(n746) );
  INV_X1 U549 ( .A(n3434), .ZN(n747) );
  INV_X1 U550 ( .A(n3537), .ZN(n3533) );
  BUF_X1 U551 ( .A(DATAIN[30]), .Z(n865) );
  BUF_X1 U552 ( .A(DATAIN[5]), .Z(n797) );
  BUF_X1 U553 ( .A(DATAIN[26]), .Z(n869) );
  BUF_X1 U554 ( .A(DATAIN[22]), .Z(n873) );
  INV_X1 U555 ( .A(n3572), .ZN(n3564) );
  INV_X1 U556 ( .A(n3572), .ZN(n3565) );
  INV_X1 U557 ( .A(n3563), .ZN(n748) );
  INV_X1 U558 ( .A(n3523), .ZN(n749) );
  INV_X1 U559 ( .A(n3523), .ZN(n750) );
  INV_X1 U560 ( .A(n3438), .ZN(n751) );
  INV_X1 U561 ( .A(n3563), .ZN(n752) );
  INV_X1 U562 ( .A(n3563), .ZN(n753) );
  INV_X1 U563 ( .A(n3572), .ZN(n754) );
  INV_X1 U564 ( .A(n3572), .ZN(n755) );
  INV_X1 U565 ( .A(n3572), .ZN(n3566) );
  AND2_X1 U566 ( .A1(n1247), .A2(n1072), .ZN(n756) );
  INV_X1 U567 ( .A(n756), .ZN(n1249) );
  AND2_X1 U568 ( .A1(n1247), .A2(n1212), .ZN(n894) );
  AND2_X1 U569 ( .A1(n1178), .A2(n1352), .ZN(n757) );
  BUF_X1 U570 ( .A(DATAIN[20]), .Z(n875) );
  BUF_X1 U571 ( .A(DATAIN[21]), .Z(n888) );
  INV_X1 U572 ( .A(DATAIN[10]), .ZN(n758) );
  INV_X1 U573 ( .A(DATAIN[10]), .ZN(n759) );
  INV_X1 U574 ( .A(DATAIN[10]), .ZN(n4201) );
  INV_X1 U575 ( .A(n32), .ZN(n760) );
  INV_X1 U576 ( .A(n3537), .ZN(n761) );
  INV_X1 U577 ( .A(n3537), .ZN(n762) );
  INV_X1 U578 ( .A(n3537), .ZN(n3534) );
  INV_X1 U579 ( .A(n3484), .ZN(n763) );
  INV_X1 U580 ( .A(n3484), .ZN(n764) );
  INV_X1 U581 ( .A(n3491), .ZN(n765) );
  INV_X1 U582 ( .A(DATAIN[0]), .ZN(n766) );
  INV_X1 U583 ( .A(DATAIN[0]), .ZN(n767) );
  INV_X1 U584 ( .A(DATAIN[0]), .ZN(n4211) );
  INV_X1 U585 ( .A(ADD_WR[2]), .ZN(n768) );
  BUF_X2 U586 ( .A(n1108), .Z(n3563) );
  BUF_X2 U587 ( .A(n1560), .Z(n3342) );
  AND3_X1 U588 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n1069) );
  INV_X1 U589 ( .A(n699), .ZN(n769) );
  INV_X1 U590 ( .A(n699), .ZN(n770) );
  INV_X1 U591 ( .A(n699), .ZN(n4193) );
  INV_X1 U592 ( .A(n193), .ZN(n772) );
  INV_X1 U593 ( .A(n193), .ZN(n773) );
  INV_X1 U594 ( .A(n193), .ZN(n4194) );
  INV_X1 U595 ( .A(n711), .ZN(n775) );
  INV_X1 U596 ( .A(n711), .ZN(n776) );
  INV_X1 U597 ( .A(DATAIN[16]), .ZN(n4195) );
  INV_X1 U598 ( .A(n701), .ZN(n778) );
  INV_X1 U599 ( .A(n701), .ZN(n779) );
  INV_X1 U600 ( .A(n701), .ZN(n4196) );
  INV_X1 U601 ( .A(n703), .ZN(n781) );
  INV_X1 U602 ( .A(n703), .ZN(n782) );
  INV_X1 U603 ( .A(n703), .ZN(n4197) );
  INV_X1 U604 ( .A(n191), .ZN(n784) );
  INV_X1 U605 ( .A(n191), .ZN(n785) );
  INV_X1 U606 ( .A(n191), .ZN(n4198) );
  INV_X1 U607 ( .A(n707), .ZN(n786) );
  INV_X1 U608 ( .A(n707), .ZN(n787) );
  INV_X1 U609 ( .A(n707), .ZN(n4199) );
  INV_X1 U610 ( .A(DATAIN[11]), .ZN(n789) );
  INV_X1 U611 ( .A(DATAIN[11]), .ZN(n790) );
  INV_X1 U612 ( .A(DATAIN[11]), .ZN(n4200) );
  BUF_X2 U613 ( .A(DATAIN[19]), .Z(n792) );
  BUF_X2 U614 ( .A(DATAIN[5]), .Z(n798) );
  BUF_X2 U615 ( .A(DATAIN[3]), .Z(n800) );
  BUF_X2 U616 ( .A(DATAIN[28]), .Z(n868) );
  BUF_X2 U617 ( .A(DATAIN[26]), .Z(n870) );
  BUF_X2 U618 ( .A(DATAIN[24]), .Z(n872) );
  BUF_X2 U619 ( .A(DATAIN[20]), .Z(n876) );
  BUF_X2 U620 ( .A(DATAIN[31]), .Z(n878) );
  BUF_X2 U621 ( .A(DATAIN[9]), .Z(n879) );
  BUF_X2 U622 ( .A(DATAIN[6]), .Z(n881) );
  BUF_X2 U623 ( .A(DATAIN[29]), .Z(n883) );
  BUF_X2 U624 ( .A(DATAIN[27]), .Z(n885) );
  BUF_X2 U625 ( .A(DATAIN[25]), .Z(n886) );
  BUF_X2 U626 ( .A(DATAIN[21]), .Z(n889) );
  BUF_X2 U627 ( .A(DATAIN[2]), .Z(n890) );
  BUF_X2 U628 ( .A(DATAIN[1]), .Z(n892) );
  CLKBUF_X1 U629 ( .A(n177), .Z(n3551) );
  CLKBUF_X1 U630 ( .A(n177), .Z(n3552) );
  CLKBUF_X1 U631 ( .A(n177), .Z(n3553) );
  CLKBUF_X1 U632 ( .A(n573), .Z(n3554) );
  CLKBUF_X1 U633 ( .A(n573), .Z(n3555) );
  CLKBUF_X1 U634 ( .A(n553), .Z(n3544) );
  CLKBUF_X1 U635 ( .A(n551), .Z(n3417) );
  CLKBUF_X1 U636 ( .A(n562), .Z(n3375) );
  CLKBUF_X1 U637 ( .A(n562), .Z(n3376) );
  CLKBUF_X1 U638 ( .A(n562), .Z(n3377) );
  CLKBUF_X1 U639 ( .A(n562), .Z(n3378) );
  CLKBUF_X1 U640 ( .A(n562), .Z(n3379) );
  CLKBUF_X1 U641 ( .A(n562), .Z(n3380) );
  CLKBUF_X1 U642 ( .A(n574), .Z(n3365) );
  CLKBUF_X1 U643 ( .A(n574), .Z(n3366) );
  CLKBUF_X1 U644 ( .A(n574), .Z(n3367) );
  CLKBUF_X1 U645 ( .A(n574), .Z(n3368) );
  CLKBUF_X1 U646 ( .A(n574), .Z(n3369) );
  CLKBUF_X1 U647 ( .A(n574), .Z(n3370) );
  CLKBUF_X1 U648 ( .A(n549), .Z(n3348) );
  CLKBUF_X1 U649 ( .A(n268), .Z(n3461) );
  CLKBUF_X1 U650 ( .A(n268), .Z(n3462) );
  CLKBUF_X1 U651 ( .A(n268), .Z(n3463) );
  CLKBUF_X1 U652 ( .A(n894), .Z(n3464) );
  CLKBUF_X1 U653 ( .A(n268), .Z(n3465) );
  CLKBUF_X1 U654 ( .A(n268), .Z(n3466) );
  CLKBUF_X1 U655 ( .A(n1489), .Z(n3393) );
  CLKBUF_X1 U656 ( .A(n1489), .Z(n3394) );
  CLKBUF_X1 U657 ( .A(n1489), .Z(n3395) );
  CLKBUF_X1 U658 ( .A(n1489), .Z(n3396) );
  CLKBUF_X1 U659 ( .A(n1489), .Z(n3392) );
  CLKBUF_X1 U660 ( .A(n1489), .Z(n3391) );
  CLKBUF_X1 U661 ( .A(n1108), .Z(n3562) );
  CLKBUF_X1 U662 ( .A(n1317), .Z(n3483) );
  CLKBUF_X1 U663 ( .A(n1355), .Z(n3443) );
  AND2_X1 U664 ( .A1(n1352), .A2(n1069), .ZN(n893) );
  INV_X2 U665 ( .A(DATAIN[2]), .ZN(n4209) );
  INV_X1 U666 ( .A(n3523), .ZN(n3518) );
  INV_X1 U667 ( .A(n592), .ZN(n3512) );
  INV_X1 U668 ( .A(n215), .ZN(n3389) );
  INV_X1 U669 ( .A(n3385), .ZN(n3383) );
  INV_X1 U670 ( .A(n3385), .ZN(n3382) );
  INV_X1 U671 ( .A(n3491), .ZN(n3486) );
  INV_X1 U672 ( .A(n18), .ZN(n3485) );
  INV_X1 U673 ( .A(n3484), .ZN(n3478) );
  INV_X1 U674 ( .A(n3484), .ZN(n3477) );
  INV_X1 U675 ( .A(n32), .ZN(n3399) );
  INV_X1 U676 ( .A(n3407), .ZN(n3398) );
  INV_X1 U677 ( .A(n3578), .ZN(n3574) );
  INV_X1 U678 ( .A(n3578), .ZN(n3573) );
  INV_X1 U679 ( .A(n3557), .ZN(n3549) );
  INV_X1 U680 ( .A(n3557), .ZN(n3548) );
  INV_X1 U681 ( .A(n178), .ZN(n3539) );
  INV_X1 U682 ( .A(n3547), .ZN(n3538) );
  INV_X1 U683 ( .A(n3511), .ZN(n3503) );
  INV_X1 U684 ( .A(n3511), .ZN(n3502) );
  INV_X1 U685 ( .A(n3501), .ZN(n3493) );
  INV_X1 U686 ( .A(n3501), .ZN(n3492) );
  INV_X1 U687 ( .A(n3458), .ZN(n3450) );
  INV_X1 U688 ( .A(n3449), .ZN(n3447) );
  INV_X1 U689 ( .A(n3449), .ZN(n3446) );
  INV_X1 U690 ( .A(n3381), .ZN(n3373) );
  INV_X1 U691 ( .A(n3381), .ZN(n3372) );
  INV_X1 U692 ( .A(n3371), .ZN(n3363) );
  INV_X1 U693 ( .A(n3476), .ZN(n3468) );
  INV_X1 U694 ( .A(n3432), .ZN(n3424) );
  INV_X1 U695 ( .A(n3432), .ZN(n3423) );
  INV_X1 U696 ( .A(n3422), .ZN(n3414) );
  INV_X1 U697 ( .A(n3422), .ZN(n3413) );
  INV_X1 U698 ( .A(n550), .ZN(n3354) );
  INV_X1 U699 ( .A(n21), .ZN(n3353) );
  INV_X1 U700 ( .A(n164), .ZN(n3344) );
  INV_X1 U701 ( .A(n3352), .ZN(n3343) );
  INV_X1 U702 ( .A(n3467), .ZN(n3459) );
  INV_X1 U703 ( .A(n1068), .ZN(n3580) );
  INV_X1 U704 ( .A(n1068), .ZN(n3581) );
  BUF_X1 U705 ( .A(n3600), .Z(n3710) );
  BUF_X1 U706 ( .A(n3600), .Z(n3709) );
  BUF_X1 U707 ( .A(n3599), .Z(n3708) );
  BUF_X1 U708 ( .A(n3599), .Z(n3707) );
  BUF_X1 U709 ( .A(n3598), .Z(n3706) );
  BUF_X1 U710 ( .A(n3598), .Z(n3705) );
  BUF_X1 U711 ( .A(n3597), .Z(n3704) );
  BUF_X1 U712 ( .A(n3597), .Z(n3703) );
  BUF_X1 U713 ( .A(n3596), .Z(n3702) );
  BUF_X1 U714 ( .A(n3596), .Z(n3701) );
  BUF_X1 U715 ( .A(n3595), .Z(n3700) );
  BUF_X1 U716 ( .A(n3595), .Z(n3699) );
  BUF_X1 U717 ( .A(n3594), .Z(n3698) );
  BUF_X1 U718 ( .A(n3594), .Z(n3697) );
  BUF_X1 U719 ( .A(n3593), .Z(n3696) );
  BUF_X1 U720 ( .A(n3593), .Z(n3695) );
  BUF_X1 U721 ( .A(n1630), .Z(n1350) );
  BUF_X1 U722 ( .A(n1635), .Z(n1248) );
  BUF_X1 U723 ( .A(n1630), .Z(n1351) );
  BUF_X1 U724 ( .A(n1635), .Z(n1250) );
  BUF_X1 U725 ( .A(n2221), .Z(n927) );
  BUF_X1 U726 ( .A(n2226), .Z(n915) );
  BUF_X1 U727 ( .A(n2221), .Z(n928) );
  BUF_X1 U728 ( .A(n2226), .Z(n916) );
  BUF_X1 U729 ( .A(n1620), .Z(n3286) );
  BUF_X1 U730 ( .A(n1620), .Z(n3287) );
  BUF_X1 U731 ( .A(n2211), .Z(n1012) );
  BUF_X1 U732 ( .A(n2211), .Z(n1013) );
  BUF_X1 U733 ( .A(n1603), .Z(n3328) );
  BUF_X1 U734 ( .A(n1608), .Z(n3316) );
  BUF_X1 U735 ( .A(n1618), .Z(n3292) );
  BUF_X1 U736 ( .A(n1603), .Z(n3329) );
  BUF_X1 U737 ( .A(n1608), .Z(n3317) );
  BUF_X1 U738 ( .A(n1618), .Z(n3293) );
  BUF_X1 U739 ( .A(n2194), .Z(n1054) );
  BUF_X1 U740 ( .A(n2199), .Z(n1042) );
  BUF_X1 U741 ( .A(n2194), .Z(n1055) );
  BUF_X1 U742 ( .A(n2199), .Z(n1043) );
  BUF_X1 U743 ( .A(n1613), .Z(n3304) );
  BUF_X1 U744 ( .A(n1628), .Z(n1399) );
  BUF_X1 U745 ( .A(n1613), .Z(n3305) );
  BUF_X1 U746 ( .A(n1628), .Z(n1403) );
  BUF_X1 U747 ( .A(n2204), .Z(n1030) );
  BUF_X1 U748 ( .A(n2209), .Z(n1018) );
  BUF_X1 U749 ( .A(n2219), .Z(n997) );
  BUF_X1 U750 ( .A(n2204), .Z(n1031) );
  BUF_X1 U751 ( .A(n2209), .Z(n1019) );
  BUF_X1 U752 ( .A(n2219), .Z(n998) );
  BUF_X1 U753 ( .A(n1631), .Z(n1285) );
  BUF_X1 U754 ( .A(n1636), .Z(n1113) );
  BUF_X1 U755 ( .A(n1631), .Z(n1320) );
  BUF_X1 U756 ( .A(n1636), .Z(n1141) );
  BUF_X1 U757 ( .A(n2222), .Z(n924) );
  BUF_X1 U758 ( .A(n2227), .Z(n912) );
  BUF_X1 U759 ( .A(n2222), .Z(n925) );
  BUF_X1 U760 ( .A(n2227), .Z(n913) );
  BUF_X1 U761 ( .A(n1600), .Z(n3334) );
  BUF_X1 U762 ( .A(n1605), .Z(n3322) );
  BUF_X1 U763 ( .A(n1610), .Z(n3310) );
  BUF_X1 U764 ( .A(n1615), .Z(n3298) );
  BUF_X1 U765 ( .A(n1625), .Z(n1424) );
  BUF_X1 U766 ( .A(n2191), .Z(n1060) );
  BUF_X1 U767 ( .A(n2196), .Z(n1048) );
  BUF_X1 U768 ( .A(n2201), .Z(n1036) );
  BUF_X1 U769 ( .A(n2206), .Z(n1024) );
  BUF_X1 U770 ( .A(n2216), .Z(n1003) );
  BUF_X1 U771 ( .A(n1604), .Z(n3325) );
  BUF_X1 U772 ( .A(n1609), .Z(n3313) );
  BUF_X1 U773 ( .A(n1614), .Z(n3301) );
  BUF_X1 U774 ( .A(n1619), .Z(n3289) );
  BUF_X1 U775 ( .A(n1629), .Z(n1357) );
  BUF_X1 U776 ( .A(n1604), .Z(n3326) );
  BUF_X1 U777 ( .A(n1609), .Z(n3314) );
  BUF_X1 U778 ( .A(n1614), .Z(n3302) );
  BUF_X1 U779 ( .A(n1619), .Z(n3290) );
  BUF_X1 U780 ( .A(n1629), .Z(n1367) );
  BUF_X1 U781 ( .A(n2195), .Z(n1051) );
  BUF_X1 U782 ( .A(n2200), .Z(n1039) );
  BUF_X1 U783 ( .A(n2205), .Z(n1027) );
  BUF_X1 U784 ( .A(n2195), .Z(n1052) );
  BUF_X1 U785 ( .A(n2200), .Z(n1040) );
  BUF_X1 U786 ( .A(n2205), .Z(n1028) );
  BUF_X1 U787 ( .A(n2210), .Z(n1015) );
  BUF_X1 U788 ( .A(n2220), .Z(n994) );
  BUF_X1 U789 ( .A(n2210), .Z(n1016) );
  BUF_X1 U790 ( .A(n2220), .Z(n995) );
  BUF_X1 U791 ( .A(n1601), .Z(n3333) );
  BUF_X1 U792 ( .A(n1606), .Z(n3321) );
  BUF_X1 U793 ( .A(n1611), .Z(n3309) );
  BUF_X1 U794 ( .A(n1616), .Z(n3297) );
  BUF_X1 U795 ( .A(n1626), .Z(n1422) );
  BUF_X1 U797 ( .A(n2192), .Z(n1059) );
  BUF_X1 U798 ( .A(n2197), .Z(n1047) );
  BUF_X1 U799 ( .A(n2202), .Z(n1035) );
  BUF_X1 U800 ( .A(n2207), .Z(n1023) );
  BUF_X1 U801 ( .A(n2217), .Z(n1002) );
  BUF_X1 U802 ( .A(n1630), .Z(n1353) );
  BUF_X1 U803 ( .A(n1635), .Z(n1252) );
  BUF_X1 U804 ( .A(n2221), .Z(n993) );
  BUF_X1 U805 ( .A(n2226), .Z(n917) );
  BUF_X1 U806 ( .A(n1620), .Z(n3288) );
  BUF_X1 U807 ( .A(n2211), .Z(n1014) );
  BUF_X1 U808 ( .A(n1603), .Z(n3330) );
  BUF_X1 U809 ( .A(n1608), .Z(n3318) );
  BUF_X1 U810 ( .A(n2194), .Z(n1056) );
  BUF_X1 U811 ( .A(n2199), .Z(n1044) );
  BUF_X1 U812 ( .A(n1613), .Z(n3306) );
  BUF_X1 U813 ( .A(n1618), .Z(n3294) );
  BUF_X1 U814 ( .A(n1628), .Z(n1404) );
  BUF_X1 U815 ( .A(n2204), .Z(n1032) );
  BUF_X1 U816 ( .A(n2209), .Z(n1020) );
  BUF_X1 U817 ( .A(n2219), .Z(n999) );
  BUF_X1 U818 ( .A(n1631), .Z(n1349) );
  BUF_X1 U819 ( .A(n1636), .Z(n1143) );
  BUF_X1 U820 ( .A(n2222), .Z(n926) );
  BUF_X1 U821 ( .A(n2227), .Z(n914) );
  BUF_X1 U822 ( .A(n1600), .Z(n3336) );
  BUF_X1 U823 ( .A(n1605), .Z(n3324) );
  BUF_X1 U824 ( .A(n1610), .Z(n3312) );
  BUF_X1 U825 ( .A(n1615), .Z(n3300) );
  BUF_X1 U826 ( .A(n1625), .Z(n1429) );
  BUF_X1 U827 ( .A(n2191), .Z(n1062) );
  BUF_X1 U828 ( .A(n2196), .Z(n1050) );
  BUF_X1 U829 ( .A(n2201), .Z(n1038) );
  BUF_X1 U830 ( .A(n2206), .Z(n1026) );
  BUF_X1 U831 ( .A(n2216), .Z(n1005) );
  BUF_X1 U832 ( .A(n1604), .Z(n3327) );
  BUF_X1 U833 ( .A(n1609), .Z(n3315) );
  BUF_X1 U834 ( .A(n1614), .Z(n3303) );
  BUF_X1 U835 ( .A(n1619), .Z(n3291) );
  BUF_X1 U836 ( .A(n1629), .Z(n1387) );
  BUF_X1 U837 ( .A(n2195), .Z(n1053) );
  BUF_X1 U838 ( .A(n2200), .Z(n1041) );
  BUF_X1 U839 ( .A(n2205), .Z(n1029) );
  BUF_X1 U840 ( .A(n2210), .Z(n1017) );
  BUF_X1 U841 ( .A(n2220), .Z(n996) );
  BUF_X1 U842 ( .A(n1623), .Z(n1556) );
  BUF_X1 U843 ( .A(n1638), .Z(n1066) );
  BUF_X1 U844 ( .A(n1623), .Z(n1557) );
  BUF_X1 U845 ( .A(n1638), .Z(n1067) );
  BUF_X1 U846 ( .A(n2214), .Z(n1009) );
  BUF_X1 U847 ( .A(n2229), .Z(n909) );
  BUF_X1 U848 ( .A(n2214), .Z(n1010) );
  BUF_X1 U849 ( .A(n2229), .Z(n910) );
  BUF_X1 U850 ( .A(n1633), .Z(n1280) );
  BUF_X1 U851 ( .A(n1633), .Z(n1281) );
  BUF_X1 U852 ( .A(n2224), .Z(n921) );
  BUF_X1 U853 ( .A(n2224), .Z(n922) );
  BUF_X1 U854 ( .A(n1624), .Z(n1432) );
  BUF_X1 U855 ( .A(n1639), .Z(n1063) );
  BUF_X1 U856 ( .A(n1624), .Z(n1445) );
  BUF_X1 U857 ( .A(n1639), .Z(n1064) );
  BUF_X1 U858 ( .A(n2215), .Z(n1006) );
  BUF_X1 U859 ( .A(n2230), .Z(n906) );
  BUF_X1 U860 ( .A(n2215), .Z(n1007) );
  BUF_X1 U861 ( .A(n2230), .Z(n907) );
  BUF_X1 U862 ( .A(n1634), .Z(n1254) );
  BUF_X1 U863 ( .A(n1634), .Z(n1258) );
  BUF_X1 U864 ( .A(n2225), .Z(n918) );
  BUF_X1 U865 ( .A(n2225), .Z(n919) );
  BUF_X1 U866 ( .A(n1623), .Z(n1558) );
  BUF_X1 U867 ( .A(n1638), .Z(n1071) );
  BUF_X1 U868 ( .A(n2214), .Z(n1011) );
  BUF_X1 U869 ( .A(n2229), .Z(n911) );
  BUF_X1 U870 ( .A(n1633), .Z(n1282) );
  BUF_X1 U871 ( .A(n2224), .Z(n923) );
  NAND2_X1 U872 ( .A1(n1106), .A2(n1070), .ZN(n1074) );
  NAND2_X1 U873 ( .A1(n1140), .A2(n1070), .ZN(n1108) );
  NAND2_X1 U874 ( .A1(n1178), .A2(n1070), .ZN(n1146) );
  NAND2_X1 U875 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
  BUF_X1 U876 ( .A(n1624), .Z(n1555) );
  BUF_X1 U877 ( .A(n1639), .Z(n1065) );
  BUF_X1 U878 ( .A(n2215), .Z(n1008) );
  BUF_X1 U879 ( .A(n2230), .Z(n908) );
  BUF_X1 U880 ( .A(n1634), .Z(n1266) );
  BUF_X1 U881 ( .A(n2225), .Z(n920) );
  BUF_X1 U882 ( .A(n1601), .Z(n3331) );
  BUF_X1 U883 ( .A(n1606), .Z(n3319) );
  BUF_X1 U884 ( .A(n1611), .Z(n3307) );
  BUF_X1 U885 ( .A(n1616), .Z(n3295) );
  BUF_X1 U886 ( .A(n1626), .Z(n1420) );
  BUF_X1 U887 ( .A(n1601), .Z(n3332) );
  BUF_X1 U888 ( .A(n1606), .Z(n3320) );
  BUF_X1 U889 ( .A(n1611), .Z(n3308) );
  BUF_X1 U890 ( .A(n1616), .Z(n3296) );
  BUF_X1 U891 ( .A(n1626), .Z(n1421) );
  BUF_X1 U892 ( .A(n2192), .Z(n1057) );
  BUF_X1 U893 ( .A(n2197), .Z(n1045) );
  BUF_X1 U894 ( .A(n2202), .Z(n1033) );
  BUF_X1 U895 ( .A(n2207), .Z(n1021) );
  BUF_X1 U896 ( .A(n2217), .Z(n1000) );
  BUF_X1 U897 ( .A(n2192), .Z(n1058) );
  BUF_X1 U899 ( .A(n2197), .Z(n1046) );
  BUF_X1 U900 ( .A(n2202), .Z(n1034) );
  BUF_X1 U901 ( .A(n2207), .Z(n1022) );
  BUF_X1 U902 ( .A(n2217), .Z(n1001) );
  BUF_X1 U903 ( .A(n1600), .Z(n3335) );
  BUF_X1 U904 ( .A(n1605), .Z(n3323) );
  BUF_X1 U905 ( .A(n1610), .Z(n3311) );
  BUF_X1 U906 ( .A(n1615), .Z(n3299) );
  BUF_X1 U907 ( .A(n1625), .Z(n1427) );
  BUF_X1 U908 ( .A(n2191), .Z(n1061) );
  BUF_X1 U909 ( .A(n2196), .Z(n1049) );
  BUF_X1 U910 ( .A(n2201), .Z(n1037) );
  BUF_X1 U911 ( .A(n2206), .Z(n1025) );
  BUF_X1 U912 ( .A(n2216), .Z(n1004) );
  NAND2_X1 U913 ( .A1(n1070), .A2(n1212), .ZN(n1180) );
  NAND2_X1 U914 ( .A1(n1247), .A2(n1069), .ZN(n1215) );
  NAND2_X1 U915 ( .A1(n1352), .A2(n1106), .ZN(n1355) );
  NAND2_X1 U916 ( .A1(n1352), .A2(n1140), .ZN(n1388) );
  NAND2_X1 U917 ( .A1(n1521), .A2(n1072), .ZN(n1523) );
  NAND2_X1 U918 ( .A1(n1178), .A2(n1521), .ZN(n1560) );
  NAND2_X1 U919 ( .A1(n1142), .A2(n1247), .ZN(n1284) );
  NAND2_X1 U920 ( .A1(n1247), .A2(n1144), .ZN(n1317) );
  NAND2_X1 U921 ( .A1(n1352), .A2(n1212), .ZN(n1456) );
  AND2_X1 U922 ( .A1(n1142), .A2(n1070), .ZN(n895) );
  AND2_X1 U923 ( .A1(n379), .A2(n1070), .ZN(n896) );
  AND2_X1 U924 ( .A1(n1106), .A2(n548), .ZN(n897) );
  AND2_X1 U925 ( .A1(n548), .A2(n1140), .ZN(n898) );
  AND2_X1 U926 ( .A1(n1106), .A2(n1521), .ZN(n899) );
  AND2_X1 U927 ( .A1(n1140), .A2(n1521), .ZN(n900) );
  AND2_X1 U928 ( .A1(n1247), .A2(n1178), .ZN(n901) );
  AND2_X1 U929 ( .A1(n360), .A2(n1352), .ZN(n902) );
  AND2_X1 U930 ( .A1(n379), .A2(n1352), .ZN(n903) );
  AND2_X1 U931 ( .A1(n379), .A2(n1521), .ZN(n905) );
  BUF_X1 U933 ( .A(n3601), .Z(n3600) );
  BUF_X1 U934 ( .A(n3601), .Z(n3599) );
  BUF_X1 U935 ( .A(n3601), .Z(n3598) );
  BUF_X1 U936 ( .A(n3602), .Z(n3597) );
  BUF_X1 U937 ( .A(n3602), .Z(n3596) );
  BUF_X1 U938 ( .A(n3602), .Z(n3595) );
  BUF_X1 U939 ( .A(n3603), .Z(n3594) );
  BUF_X1 U940 ( .A(n3603), .Z(n3593) );
  NAND2_X1 U941 ( .A1(n2160), .A2(n2168), .ZN(n1611) );
  NAND2_X1 U942 ( .A1(n2751), .A2(n2759), .ZN(n2202) );
  NAND2_X1 U943 ( .A1(n2160), .A2(n2169), .ZN(n1610) );
  NAND2_X1 U944 ( .A1(n2751), .A2(n2760), .ZN(n2201) );
  INV_X1 U945 ( .A(ADD_WR[2]), .ZN(n4171) );
  INV_X1 U946 ( .A(ADD_WR[1]), .ZN(n4172) );
  INV_X1 U947 ( .A(ADD_WR[0]), .ZN(n4173) );
  NAND2_X1 U948 ( .A1(n2174), .A2(n2160), .ZN(n1624) );
  NAND2_X1 U949 ( .A1(n2175), .A2(n2160), .ZN(n1623) );
  NAND2_X1 U950 ( .A1(n2179), .A2(n2160), .ZN(n1639) );
  NAND2_X1 U951 ( .A1(n2180), .A2(n2160), .ZN(n1638) );
  NAND2_X1 U952 ( .A1(n2765), .A2(n2751), .ZN(n2215) );
  NAND2_X1 U953 ( .A1(n2766), .A2(n2751), .ZN(n2214) );
  NAND2_X1 U954 ( .A1(n2770), .A2(n2751), .ZN(n2230) );
  NAND2_X1 U955 ( .A1(n2771), .A2(n2751), .ZN(n2229) );
  AND2_X1 U956 ( .A1(n2171), .A2(n4179), .ZN(n2168) );
  AND2_X1 U957 ( .A1(n2762), .A2(n4176), .ZN(n2759) );
  NAND2_X1 U958 ( .A1(n2159), .A2(n2162), .ZN(n1601) );
  AND2_X1 U959 ( .A1(n2182), .A2(n4179), .ZN(n2180) );
  AND2_X1 U960 ( .A1(n2773), .A2(n4176), .ZN(n2771) );
  AND2_X1 U961 ( .A1(n2166), .A2(n4179), .ZN(n2159) );
  AND2_X1 U962 ( .A1(n2757), .A2(n4176), .ZN(n2750) );
  NAND2_X1 U963 ( .A1(n2750), .A2(n2753), .ZN(n2192) );
  NAND2_X1 U964 ( .A1(n2159), .A2(n2165), .ZN(n1606) );
  NAND2_X1 U965 ( .A1(n2175), .A2(n2165), .ZN(n1626) );
  NAND2_X1 U966 ( .A1(n2750), .A2(n2756), .ZN(n2197) );
  NAND2_X1 U967 ( .A1(n2766), .A2(n2756), .ZN(n2217) );
  NAND2_X1 U968 ( .A1(n2168), .A2(n2164), .ZN(n1616) );
  NAND2_X1 U969 ( .A1(n2180), .A2(n2164), .ZN(n1633) );
  NAND2_X1 U970 ( .A1(n2179), .A2(n2164), .ZN(n1634) );
  NAND2_X1 U971 ( .A1(n2759), .A2(n2755), .ZN(n2207) );
  NAND2_X1 U972 ( .A1(n2771), .A2(n2755), .ZN(n2224) );
  NAND2_X1 U973 ( .A1(n2770), .A2(n2755), .ZN(n2225) );
  NAND2_X1 U974 ( .A1(n2161), .A2(n2162), .ZN(n1600) );
  NAND2_X1 U975 ( .A1(n2752), .A2(n2753), .ZN(n2191) );
  NAND2_X1 U976 ( .A1(n2164), .A2(n2169), .ZN(n1615) );
  NAND2_X1 U977 ( .A1(n2755), .A2(n2760), .ZN(n2206) );
  AND2_X1 U978 ( .A1(n2177), .A2(n4179), .ZN(n2175) );
  AND2_X1 U979 ( .A1(n2768), .A2(n4176), .ZN(n2766) );
  NAND2_X1 U980 ( .A1(n2161), .A2(n2165), .ZN(n1605) );
  NAND2_X1 U981 ( .A1(n2174), .A2(n2165), .ZN(n1625) );
  NAND2_X1 U982 ( .A1(n2752), .A2(n2756), .ZN(n2196) );
  NAND2_X1 U983 ( .A1(n2765), .A2(n2756), .ZN(n2216) );
  AND2_X1 U984 ( .A1(n2159), .A2(n2160), .ZN(n1604) );
  AND2_X1 U985 ( .A1(n2161), .A2(n2160), .ZN(n1603) );
  AND2_X1 U986 ( .A1(n2750), .A2(n2751), .ZN(n2195) );
  AND2_X1 U987 ( .A1(n2752), .A2(n2751), .ZN(n2194) );
  AND2_X1 U988 ( .A1(n2162), .A2(n2168), .ZN(n1614) );
  AND2_X1 U989 ( .A1(n2162), .A2(n2169), .ZN(n1613) );
  AND2_X1 U990 ( .A1(n2753), .A2(n2759), .ZN(n2205) );
  AND2_X1 U991 ( .A1(n2753), .A2(n2760), .ZN(n2204) );
  AND2_X1 U992 ( .A1(n2174), .A2(n2162), .ZN(n1620) );
  AND2_X1 U993 ( .A1(n2179), .A2(n2162), .ZN(n1635) );
  AND2_X1 U994 ( .A1(n2180), .A2(n2162), .ZN(n1636) );
  AND2_X1 U995 ( .A1(n2765), .A2(n2753), .ZN(n2211) );
  AND2_X1 U996 ( .A1(n2770), .A2(n2753), .ZN(n2226) );
  AND2_X1 U997 ( .A1(n2771), .A2(n2753), .ZN(n2227) );
  AND2_X1 U998 ( .A1(n2165), .A2(n2168), .ZN(n1619) );
  AND2_X1 U999 ( .A1(n2165), .A2(n2169), .ZN(n1618) );
  AND2_X1 U1000 ( .A1(n2756), .A2(n2759), .ZN(n2210) );
  AND2_X1 U1001 ( .A1(n2756), .A2(n2760), .ZN(n2209) );
  AND2_X1 U1002 ( .A1(n2179), .A2(n2165), .ZN(n1630) );
  AND2_X1 U1003 ( .A1(n2180), .A2(n2165), .ZN(n1631) );
  AND2_X1 U1004 ( .A1(n2770), .A2(n2756), .ZN(n2221) );
  AND2_X1 U1005 ( .A1(n2771), .A2(n2756), .ZN(n2222) );
  AND2_X1 U1006 ( .A1(n2159), .A2(n2164), .ZN(n1609) );
  AND2_X1 U1007 ( .A1(n2161), .A2(n2164), .ZN(n1608) );
  AND2_X1 U1008 ( .A1(n2175), .A2(n2164), .ZN(n1629) );
  AND2_X1 U1009 ( .A1(n2174), .A2(n2164), .ZN(n1628) );
  AND2_X1 U1010 ( .A1(n2750), .A2(n2755), .ZN(n2200) );
  AND2_X1 U1011 ( .A1(n2752), .A2(n2755), .ZN(n2199) );
  AND2_X1 U1012 ( .A1(n2766), .A2(n2755), .ZN(n2220) );
  AND2_X1 U1013 ( .A1(n2765), .A2(n2755), .ZN(n2219) );
  INV_X1 U1014 ( .A(ADD_WR[4]), .ZN(n3923) );
  INV_X1 U1015 ( .A(ADD_WR[3]), .ZN(n4170) );
  BUF_X1 U1016 ( .A(RST_AN), .Z(n3601) );
  BUF_X1 U1017 ( .A(RST_AN), .Z(n3602) );
  BUF_X1 U1018 ( .A(RST_AN), .Z(n3603) );
  NOR2_X1 U1019 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n2162) );
  NOR2_X1 U1020 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2753) );
  NOR4_X1 U1021 ( .A1(n1780), .A2(n1781), .A3(n1782), .A4(n1783), .ZN(n1779)
         );
  OAI221_X1 U1022 ( .B1(n970), .B2(n3300), .C1(n938), .C2(n3297), .A(n1787), 
        .ZN(n1780) );
  OAI221_X1 U1023 ( .B1(n842), .B2(n3312), .C1(n810), .C2(n3309), .A(n1786), 
        .ZN(n1781) );
  OAI221_X1 U1024 ( .B1(n650), .B2(n3324), .C1(n618), .C2(n3321), .A(n1785), 
        .ZN(n1782) );
  NOR4_X1 U1025 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .ZN(n1762)
         );
  OAI221_X1 U1026 ( .B1(n969), .B2(n3300), .C1(n937), .C2(n3297), .A(n1770), 
        .ZN(n1763) );
  OAI221_X1 U1027 ( .B1(n841), .B2(n3312), .C1(n809), .C2(n3309), .A(n1769), 
        .ZN(n1764) );
  OAI221_X1 U1028 ( .B1(n649), .B2(n3324), .C1(n617), .C2(n3321), .A(n1768), 
        .ZN(n1765) );
  NOR4_X1 U1029 ( .A1(n1746), .A2(n1747), .A3(n1748), .A4(n1749), .ZN(n1745)
         );
  OAI221_X1 U1030 ( .B1(n968), .B2(n3300), .C1(n936), .C2(n3297), .A(n1753), 
        .ZN(n1746) );
  OAI221_X1 U1031 ( .B1(n840), .B2(n3312), .C1(n808), .C2(n3309), .A(n1752), 
        .ZN(n1747) );
  OAI221_X1 U1032 ( .B1(n648), .B2(n3324), .C1(n616), .C2(n3321), .A(n1751), 
        .ZN(n1748) );
  NOR4_X1 U1033 ( .A1(n1729), .A2(n1730), .A3(n1731), .A4(n1732), .ZN(n1728)
         );
  OAI221_X1 U1035 ( .B1(n967), .B2(n3300), .C1(n935), .C2(n3297), .A(n1736), 
        .ZN(n1729) );
  OAI221_X1 U1038 ( .B1(n839), .B2(n3312), .C1(n807), .C2(n3309), .A(n1735), 
        .ZN(n1730) );
  OAI221_X1 U1039 ( .B1(n647), .B2(n3324), .C1(n615), .C2(n3321), .A(n1734), 
        .ZN(n1731) );
  NOR4_X1 U1040 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711)
         );
  OAI221_X1 U1041 ( .B1(n966), .B2(n3300), .C1(n934), .C2(n3297), .A(n1719), 
        .ZN(n1712) );
  OAI221_X1 U1042 ( .B1(n838), .B2(n3312), .C1(n806), .C2(n3309), .A(n1718), 
        .ZN(n1713) );
  OAI221_X1 U1043 ( .B1(n646), .B2(n3324), .C1(n614), .C2(n3321), .A(n1717), 
        .ZN(n1714) );
  NOR4_X1 U1044 ( .A1(n1695), .A2(n1696), .A3(n1697), .A4(n1698), .ZN(n1694)
         );
  OAI221_X1 U1045 ( .B1(n965), .B2(n3300), .C1(n933), .C2(n3297), .A(n1702), 
        .ZN(n1695) );
  OAI221_X1 U1046 ( .B1(n837), .B2(n3312), .C1(n805), .C2(n3309), .A(n1701), 
        .ZN(n1696) );
  OAI221_X1 U1047 ( .B1(n645), .B2(n3324), .C1(n613), .C2(n3321), .A(n1700), 
        .ZN(n1697) );
  NOR4_X1 U1048 ( .A1(n1678), .A2(n1679), .A3(n1680), .A4(n1681), .ZN(n1677)
         );
  OAI221_X1 U1049 ( .B1(n964), .B2(n3300), .C1(n932), .C2(n3297), .A(n1685), 
        .ZN(n1678) );
  OAI221_X1 U1050 ( .B1(n836), .B2(n3312), .C1(n804), .C2(n3309), .A(n1684), 
        .ZN(n1679) );
  OAI221_X1 U1051 ( .B1(n644), .B2(n3324), .C1(n612), .C2(n3321), .A(n1683), 
        .ZN(n1680) );
  NOR4_X1 U1052 ( .A1(n1661), .A2(n1662), .A3(n1663), .A4(n1664), .ZN(n1660)
         );
  OAI221_X1 U1053 ( .B1(n963), .B2(n3300), .C1(n931), .C2(n3297), .A(n1668), 
        .ZN(n1661) );
  OAI221_X1 U1054 ( .B1(n835), .B2(n3312), .C1(n803), .C2(n3309), .A(n1667), 
        .ZN(n1662) );
  OAI221_X1 U1055 ( .B1(n643), .B2(n3324), .C1(n611), .C2(n3321), .A(n1666), 
        .ZN(n1663) );
  NOR4_X1 U1056 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .ZN(n1643)
         );
  OAI221_X1 U1057 ( .B1(n962), .B2(n3300), .C1(n930), .C2(n3297), .A(n1651), 
        .ZN(n1644) );
  OAI221_X1 U1058 ( .B1(n834), .B2(n3312), .C1(n802), .C2(n3309), .A(n1650), 
        .ZN(n1645) );
  OAI221_X1 U1059 ( .B1(n642), .B2(n3324), .C1(n610), .C2(n3321), .A(n1649), 
        .ZN(n1646) );
  NOR4_X1 U1060 ( .A1(n1596), .A2(n1597), .A3(n1598), .A4(n1599), .ZN(n1595)
         );
  OAI221_X1 U1061 ( .B1(n961), .B2(n3300), .C1(n929), .C2(n3297), .A(n1617), 
        .ZN(n1596) );
  OAI221_X1 U1062 ( .B1(n833), .B2(n3312), .C1(n801), .C2(n3309), .A(n1612), 
        .ZN(n1597) );
  OAI221_X1 U1063 ( .B1(n641), .B2(n3324), .C1(n609), .C2(n3321), .A(n1607), 
        .ZN(n1598) );
  NOR4_X1 U1064 ( .A1(n2371), .A2(n2372), .A3(n2373), .A4(n2374), .ZN(n2370)
         );
  OAI221_X1 U1065 ( .B1(n970), .B2(n1026), .C1(n938), .C2(n1023), .A(n2378), 
        .ZN(n2371) );
  OAI221_X1 U1066 ( .B1(n842), .B2(n1038), .C1(n810), .C2(n1035), .A(n2377), 
        .ZN(n2372) );
  OAI221_X1 U1067 ( .B1(n650), .B2(n1050), .C1(n618), .C2(n1047), .A(n2376), 
        .ZN(n2373) );
  NOR4_X1 U1068 ( .A1(n2354), .A2(n2355), .A3(n2356), .A4(n2357), .ZN(n2353)
         );
  OAI221_X1 U1069 ( .B1(n969), .B2(n1026), .C1(n937), .C2(n1023), .A(n2361), 
        .ZN(n2354) );
  OAI221_X1 U1070 ( .B1(n841), .B2(n1038), .C1(n809), .C2(n1035), .A(n2360), 
        .ZN(n2355) );
  OAI221_X1 U1071 ( .B1(n649), .B2(n1050), .C1(n617), .C2(n1047), .A(n2359), 
        .ZN(n2356) );
  NOR4_X1 U1072 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n2336)
         );
  OAI221_X1 U1073 ( .B1(n968), .B2(n1026), .C1(n936), .C2(n1023), .A(n2344), 
        .ZN(n2337) );
  OAI221_X1 U1074 ( .B1(n840), .B2(n1038), .C1(n808), .C2(n1035), .A(n2343), 
        .ZN(n2338) );
  OAI221_X1 U1075 ( .B1(n648), .B2(n1050), .C1(n616), .C2(n1047), .A(n2342), 
        .ZN(n2339) );
  NOR4_X1 U1076 ( .A1(n2320), .A2(n2321), .A3(n2322), .A4(n2323), .ZN(n2319)
         );
  OAI221_X1 U1077 ( .B1(n967), .B2(n1026), .C1(n935), .C2(n1023), .A(n2327), 
        .ZN(n2320) );
  OAI221_X1 U1078 ( .B1(n839), .B2(n1038), .C1(n807), .C2(n1035), .A(n2326), 
        .ZN(n2321) );
  OAI221_X1 U1079 ( .B1(n647), .B2(n1050), .C1(n615), .C2(n1047), .A(n2325), 
        .ZN(n2322) );
  NOR4_X1 U1080 ( .A1(n2303), .A2(n2304), .A3(n2305), .A4(n2306), .ZN(n2302)
         );
  OAI221_X1 U1081 ( .B1(n966), .B2(n1026), .C1(n934), .C2(n1023), .A(n2310), 
        .ZN(n2303) );
  OAI221_X1 U1082 ( .B1(n838), .B2(n1038), .C1(n806), .C2(n1035), .A(n2309), 
        .ZN(n2304) );
  OAI221_X1 U1083 ( .B1(n646), .B2(n1050), .C1(n614), .C2(n1047), .A(n2308), 
        .ZN(n2305) );
  NOR4_X1 U1084 ( .A1(n2286), .A2(n2287), .A3(n2288), .A4(n2289), .ZN(n2285)
         );
  OAI221_X1 U1085 ( .B1(n965), .B2(n1026), .C1(n933), .C2(n1023), .A(n2293), 
        .ZN(n2286) );
  OAI221_X1 U1086 ( .B1(n837), .B2(n1038), .C1(n805), .C2(n1035), .A(n2292), 
        .ZN(n2287) );
  OAI221_X1 U1087 ( .B1(n645), .B2(n1050), .C1(n613), .C2(n1047), .A(n2291), 
        .ZN(n2288) );
  NOR4_X1 U1088 ( .A1(n2269), .A2(n2270), .A3(n2271), .A4(n2272), .ZN(n2268)
         );
  OAI221_X1 U1089 ( .B1(n964), .B2(n1026), .C1(n932), .C2(n1023), .A(n2276), 
        .ZN(n2269) );
  OAI221_X1 U1090 ( .B1(n836), .B2(n1038), .C1(n804), .C2(n1035), .A(n2275), 
        .ZN(n2270) );
  OAI221_X1 U1091 ( .B1(n644), .B2(n1050), .C1(n612), .C2(n1047), .A(n2274), 
        .ZN(n2271) );
  NOR4_X1 U1092 ( .A1(n2252), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2251)
         );
  OAI221_X1 U1093 ( .B1(n963), .B2(n1026), .C1(n931), .C2(n1023), .A(n2259), 
        .ZN(n2252) );
  OAI221_X1 U1094 ( .B1(n835), .B2(n1038), .C1(n803), .C2(n1035), .A(n2258), 
        .ZN(n2253) );
  OAI221_X1 U1095 ( .B1(n643), .B2(n1050), .C1(n611), .C2(n1047), .A(n2257), 
        .ZN(n2254) );
  NOR4_X1 U1096 ( .A1(n2235), .A2(n2236), .A3(n2237), .A4(n2238), .ZN(n2234)
         );
  OAI221_X1 U1097 ( .B1(n962), .B2(n1026), .C1(n930), .C2(n1023), .A(n2242), 
        .ZN(n2235) );
  OAI221_X1 U1098 ( .B1(n834), .B2(n1038), .C1(n802), .C2(n1035), .A(n2241), 
        .ZN(n2236) );
  OAI221_X1 U1099 ( .B1(n642), .B2(n1050), .C1(n610), .C2(n1047), .A(n2240), 
        .ZN(n2237) );
  NOR4_X1 U1100 ( .A1(n2187), .A2(n2188), .A3(n2189), .A4(n2190), .ZN(n2186)
         );
  OAI221_X1 U1101 ( .B1(n961), .B2(n1026), .C1(n929), .C2(n1023), .A(n2208), 
        .ZN(n2187) );
  OAI221_X1 U1102 ( .B1(n833), .B2(n1038), .C1(n801), .C2(n1035), .A(n2203), 
        .ZN(n2188) );
  OAI221_X1 U1103 ( .B1(n641), .B2(n1050), .C1(n609), .C2(n1047), .A(n2198), 
        .ZN(n2189) );
  NOR4_X1 U1104 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2153)
         );
  OAI221_X1 U1105 ( .B1(n992), .B2(n3298), .C1(n960), .C2(n3295), .A(n2170), 
        .ZN(n2154) );
  OAI221_X1 U1106 ( .B1(n864), .B2(n3310), .C1(n832), .C2(n3307), .A(n2167), 
        .ZN(n2155) );
  OAI221_X1 U1107 ( .B1(n672), .B2(n3322), .C1(n640), .C2(n3319), .A(n2163), 
        .ZN(n2156) );
  NOR4_X1 U1108 ( .A1(n2137), .A2(n2138), .A3(n2139), .A4(n2140), .ZN(n2136)
         );
  OAI221_X1 U1109 ( .B1(n991), .B2(n3298), .C1(n959), .C2(n3295), .A(n2144), 
        .ZN(n2137) );
  OAI221_X1 U1110 ( .B1(n863), .B2(n3310), .C1(n831), .C2(n3307), .A(n2143), 
        .ZN(n2138) );
  OAI221_X1 U1111 ( .B1(n671), .B2(n3322), .C1(n639), .C2(n3319), .A(n2142), 
        .ZN(n2139) );
  NOR4_X1 U1112 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2119)
         );
  OAI221_X1 U1113 ( .B1(n990), .B2(n3298), .C1(n958), .C2(n3295), .A(n2127), 
        .ZN(n2120) );
  OAI221_X1 U1114 ( .B1(n862), .B2(n3310), .C1(n830), .C2(n3307), .A(n2126), 
        .ZN(n2121) );
  OAI221_X1 U1115 ( .B1(n670), .B2(n3322), .C1(n638), .C2(n3319), .A(n2125), 
        .ZN(n2122) );
  NOR4_X1 U1116 ( .A1(n2103), .A2(n2104), .A3(n2105), .A4(n2106), .ZN(n2102)
         );
  OAI221_X1 U1117 ( .B1(n989), .B2(n3298), .C1(n957), .C2(n3295), .A(n2110), 
        .ZN(n2103) );
  OAI221_X1 U1118 ( .B1(n861), .B2(n3310), .C1(n829), .C2(n3307), .A(n2109), 
        .ZN(n2104) );
  OAI221_X1 U1119 ( .B1(n669), .B2(n3322), .C1(n637), .C2(n3319), .A(n2108), 
        .ZN(n2105) );
  NOR4_X1 U1120 ( .A1(n2086), .A2(n2087), .A3(n2088), .A4(n2089), .ZN(n2085)
         );
  OAI221_X1 U1121 ( .B1(n988), .B2(n3298), .C1(n956), .C2(n3295), .A(n2093), 
        .ZN(n2086) );
  OAI221_X1 U1122 ( .B1(n860), .B2(n3310), .C1(n828), .C2(n3307), .A(n2092), 
        .ZN(n2087) );
  OAI221_X1 U1123 ( .B1(n668), .B2(n3322), .C1(n636), .C2(n3319), .A(n2091), 
        .ZN(n2088) );
  NOR4_X1 U1124 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2068)
         );
  OAI221_X1 U1125 ( .B1(n987), .B2(n3298), .C1(n955), .C2(n3295), .A(n2076), 
        .ZN(n2069) );
  OAI221_X1 U1126 ( .B1(n859), .B2(n3310), .C1(n827), .C2(n3307), .A(n2075), 
        .ZN(n2070) );
  OAI221_X1 U1127 ( .B1(n667), .B2(n3322), .C1(n635), .C2(n3319), .A(n2074), 
        .ZN(n2071) );
  NOR4_X1 U1128 ( .A1(n2052), .A2(n2053), .A3(n2054), .A4(n2055), .ZN(n2051)
         );
  OAI221_X1 U1129 ( .B1(n986), .B2(n3298), .C1(n954), .C2(n3295), .A(n2059), 
        .ZN(n2052) );
  OAI221_X1 U1130 ( .B1(n858), .B2(n3310), .C1(n826), .C2(n3307), .A(n2058), 
        .ZN(n2053) );
  OAI221_X1 U1131 ( .B1(n666), .B2(n3322), .C1(n634), .C2(n3319), .A(n2057), 
        .ZN(n2054) );
  NOR4_X1 U1132 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .ZN(n2034)
         );
  OAI221_X1 U1133 ( .B1(n985), .B2(n3298), .C1(n953), .C2(n3295), .A(n2042), 
        .ZN(n2035) );
  OAI221_X1 U1134 ( .B1(n857), .B2(n3310), .C1(n825), .C2(n3307), .A(n2041), 
        .ZN(n2036) );
  OAI221_X1 U1135 ( .B1(n665), .B2(n3322), .C1(n633), .C2(n3319), .A(n2040), 
        .ZN(n2037) );
  NOR4_X1 U1136 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2017)
         );
  OAI221_X1 U1137 ( .B1(n984), .B2(n3298), .C1(n952), .C2(n3295), .A(n2025), 
        .ZN(n2018) );
  OAI221_X1 U1138 ( .B1(n856), .B2(n3310), .C1(n824), .C2(n3307), .A(n2024), 
        .ZN(n2019) );
  OAI221_X1 U1139 ( .B1(n664), .B2(n3322), .C1(n632), .C2(n3319), .A(n2023), 
        .ZN(n2020) );
  NOR4_X1 U1140 ( .A1(n2001), .A2(n2002), .A3(n2003), .A4(n2004), .ZN(n2000)
         );
  OAI221_X1 U1141 ( .B1(n983), .B2(n3298), .C1(n951), .C2(n3295), .A(n2008), 
        .ZN(n2001) );
  OAI221_X1 U1142 ( .B1(n855), .B2(n3310), .C1(n823), .C2(n3307), .A(n2007), 
        .ZN(n2002) );
  OAI221_X1 U1143 ( .B1(n663), .B2(n3322), .C1(n631), .C2(n3319), .A(n2006), 
        .ZN(n2003) );
  NOR4_X1 U1144 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(n1983)
         );
  OAI221_X1 U1145 ( .B1(n982), .B2(n3298), .C1(n950), .C2(n3295), .A(n1991), 
        .ZN(n1984) );
  OAI221_X1 U1146 ( .B1(n854), .B2(n3310), .C1(n822), .C2(n3307), .A(n1990), 
        .ZN(n1985) );
  OAI221_X1 U1147 ( .B1(n662), .B2(n3322), .C1(n630), .C2(n3319), .A(n1989), 
        .ZN(n1986) );
  NOR4_X1 U1148 ( .A1(n1967), .A2(n1968), .A3(n1969), .A4(n1970), .ZN(n1966)
         );
  OAI221_X1 U1149 ( .B1(n981), .B2(n3299), .C1(n949), .C2(n3296), .A(n1974), 
        .ZN(n1967) );
  OAI221_X1 U1150 ( .B1(n853), .B2(n3311), .C1(n821), .C2(n3308), .A(n1973), 
        .ZN(n1968) );
  OAI221_X1 U1151 ( .B1(n661), .B2(n3323), .C1(n629), .C2(n3320), .A(n1972), 
        .ZN(n1969) );
  NOR4_X1 U1152 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1949)
         );
  OAI221_X1 U1153 ( .B1(n980), .B2(n3299), .C1(n948), .C2(n3296), .A(n1957), 
        .ZN(n1950) );
  OAI221_X1 U1154 ( .B1(n852), .B2(n3311), .C1(n820), .C2(n3308), .A(n1956), 
        .ZN(n1951) );
  OAI221_X1 U1155 ( .B1(n660), .B2(n3323), .C1(n628), .C2(n3320), .A(n1955), 
        .ZN(n1952) );
  NOR4_X1 U1156 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(n1932)
         );
  OAI221_X1 U1157 ( .B1(n979), .B2(n3299), .C1(n947), .C2(n3296), .A(n1940), 
        .ZN(n1933) );
  OAI221_X1 U1158 ( .B1(n851), .B2(n3311), .C1(n819), .C2(n3308), .A(n1939), 
        .ZN(n1934) );
  OAI221_X1 U1159 ( .B1(n659), .B2(n3323), .C1(n627), .C2(n3320), .A(n1938), 
        .ZN(n1935) );
  NOR4_X1 U1160 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(n1915)
         );
  OAI221_X1 U1161 ( .B1(n978), .B2(n3299), .C1(n946), .C2(n3296), .A(n1923), 
        .ZN(n1916) );
  OAI221_X1 U1162 ( .B1(n850), .B2(n3311), .C1(n818), .C2(n3308), .A(n1922), 
        .ZN(n1917) );
  OAI221_X1 U1163 ( .B1(n658), .B2(n3323), .C1(n626), .C2(n3320), .A(n1921), 
        .ZN(n1918) );
  NOR4_X1 U1164 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898)
         );
  OAI221_X1 U1165 ( .B1(n977), .B2(n3299), .C1(n945), .C2(n3296), .A(n1906), 
        .ZN(n1899) );
  OAI221_X1 U1166 ( .B1(n849), .B2(n3311), .C1(n817), .C2(n3308), .A(n1905), 
        .ZN(n1900) );
  OAI221_X1 U1167 ( .B1(n657), .B2(n3323), .C1(n625), .C2(n3320), .A(n1904), 
        .ZN(n1901) );
  NOR4_X1 U1168 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .ZN(n1881)
         );
  OAI221_X1 U1169 ( .B1(n976), .B2(n3299), .C1(n944), .C2(n3296), .A(n1889), 
        .ZN(n1882) );
  OAI221_X1 U1170 ( .B1(n848), .B2(n3311), .C1(n816), .C2(n3308), .A(n1888), 
        .ZN(n1883) );
  OAI221_X1 U1171 ( .B1(n656), .B2(n3323), .C1(n624), .C2(n3320), .A(n1887), 
        .ZN(n1884) );
  NOR4_X1 U1172 ( .A1(n1865), .A2(n1866), .A3(n1867), .A4(n1868), .ZN(n1864)
         );
  OAI221_X1 U1173 ( .B1(n975), .B2(n3299), .C1(n943), .C2(n3296), .A(n1872), 
        .ZN(n1865) );
  OAI221_X1 U1174 ( .B1(n847), .B2(n3311), .C1(n815), .C2(n3308), .A(n1871), 
        .ZN(n1866) );
  OAI221_X1 U1175 ( .B1(n655), .B2(n3323), .C1(n623), .C2(n3320), .A(n1870), 
        .ZN(n1867) );
  NOR4_X1 U1176 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1847)
         );
  OAI221_X1 U1177 ( .B1(n974), .B2(n3299), .C1(n942), .C2(n3296), .A(n1855), 
        .ZN(n1848) );
  OAI221_X1 U1178 ( .B1(n846), .B2(n3311), .C1(n814), .C2(n3308), .A(n1854), 
        .ZN(n1849) );
  OAI221_X1 U1179 ( .B1(n654), .B2(n3323), .C1(n622), .C2(n3320), .A(n1853), 
        .ZN(n1850) );
  NOR4_X1 U1180 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(n1830)
         );
  OAI221_X1 U1181 ( .B1(n973), .B2(n3299), .C1(n941), .C2(n3296), .A(n1838), 
        .ZN(n1831) );
  OAI221_X1 U1182 ( .B1(n845), .B2(n3311), .C1(n813), .C2(n3308), .A(n1837), 
        .ZN(n1832) );
  OAI221_X1 U1183 ( .B1(n653), .B2(n3323), .C1(n621), .C2(n3320), .A(n1836), 
        .ZN(n1833) );
  NOR4_X1 U1184 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .ZN(n1813)
         );
  OAI221_X1 U1185 ( .B1(n972), .B2(n3299), .C1(n940), .C2(n3296), .A(n1821), 
        .ZN(n1814) );
  OAI221_X1 U1186 ( .B1(n844), .B2(n3311), .C1(n812), .C2(n3308), .A(n1820), 
        .ZN(n1815) );
  OAI221_X1 U1187 ( .B1(n652), .B2(n3323), .C1(n620), .C2(n3320), .A(n1819), 
        .ZN(n1816) );
  NOR4_X1 U1188 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1796)
         );
  OAI221_X1 U1189 ( .B1(n971), .B2(n3299), .C1(n939), .C2(n3296), .A(n1804), 
        .ZN(n1797) );
  OAI221_X1 U1190 ( .B1(n843), .B2(n3311), .C1(n811), .C2(n3308), .A(n1803), 
        .ZN(n1798) );
  OAI221_X1 U1191 ( .B1(n651), .B2(n3323), .C1(n619), .C2(n3320), .A(n1802), 
        .ZN(n1799) );
  NOR4_X1 U1192 ( .A1(n2745), .A2(n2746), .A3(n2747), .A4(n2748), .ZN(n2744)
         );
  OAI221_X1 U1193 ( .B1(n992), .B2(n1024), .C1(n960), .C2(n1021), .A(n2761), 
        .ZN(n2745) );
  OAI221_X1 U1194 ( .B1(n864), .B2(n1036), .C1(n832), .C2(n1033), .A(n2758), 
        .ZN(n2746) );
  OAI221_X1 U1195 ( .B1(n672), .B2(n1048), .C1(n640), .C2(n1045), .A(n2754), 
        .ZN(n2747) );
  NOR4_X1 U1196 ( .A1(n2728), .A2(n2729), .A3(n2730), .A4(n2731), .ZN(n2727)
         );
  OAI221_X1 U1197 ( .B1(n991), .B2(n1024), .C1(n959), .C2(n1021), .A(n2735), 
        .ZN(n2728) );
  OAI221_X1 U1198 ( .B1(n863), .B2(n1036), .C1(n831), .C2(n1033), .A(n2734), 
        .ZN(n2729) );
  OAI221_X1 U1199 ( .B1(n671), .B2(n1048), .C1(n639), .C2(n1045), .A(n2733), 
        .ZN(n2730) );
  NOR4_X1 U1200 ( .A1(n2711), .A2(n2712), .A3(n2713), .A4(n2714), .ZN(n2710)
         );
  OAI221_X1 U1201 ( .B1(n990), .B2(n1024), .C1(n958), .C2(n1021), .A(n2718), 
        .ZN(n2711) );
  OAI221_X1 U1202 ( .B1(n862), .B2(n1036), .C1(n830), .C2(n1033), .A(n2717), 
        .ZN(n2712) );
  OAI221_X1 U1203 ( .B1(n670), .B2(n1048), .C1(n638), .C2(n1045), .A(n2716), 
        .ZN(n2713) );
  NOR4_X1 U1204 ( .A1(n2694), .A2(n2695), .A3(n2696), .A4(n2697), .ZN(n2693)
         );
  OAI221_X1 U1205 ( .B1(n989), .B2(n1024), .C1(n957), .C2(n1021), .A(n2701), 
        .ZN(n2694) );
  OAI221_X1 U1206 ( .B1(n861), .B2(n1036), .C1(n829), .C2(n1033), .A(n2700), 
        .ZN(n2695) );
  OAI221_X1 U1207 ( .B1(n669), .B2(n1048), .C1(n637), .C2(n1045), .A(n2699), 
        .ZN(n2696) );
  NOR4_X1 U1208 ( .A1(n2677), .A2(n2678), .A3(n2679), .A4(n2680), .ZN(n2676)
         );
  OAI221_X1 U1209 ( .B1(n988), .B2(n1024), .C1(n956), .C2(n1021), .A(n2684), 
        .ZN(n2677) );
  OAI221_X1 U1210 ( .B1(n860), .B2(n1036), .C1(n828), .C2(n1033), .A(n2683), 
        .ZN(n2678) );
  OAI221_X1 U1211 ( .B1(n668), .B2(n1048), .C1(n636), .C2(n1045), .A(n2682), 
        .ZN(n2679) );
  NOR4_X1 U1212 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(n2659)
         );
  OAI221_X1 U1213 ( .B1(n987), .B2(n1024), .C1(n955), .C2(n1021), .A(n2667), 
        .ZN(n2660) );
  OAI221_X1 U1214 ( .B1(n859), .B2(n1036), .C1(n827), .C2(n1033), .A(n2666), 
        .ZN(n2661) );
  OAI221_X1 U1215 ( .B1(n667), .B2(n1048), .C1(n635), .C2(n1045), .A(n2665), 
        .ZN(n2662) );
  NOR4_X1 U1216 ( .A1(n2643), .A2(n2644), .A3(n2645), .A4(n2646), .ZN(n2642)
         );
  OAI221_X1 U1217 ( .B1(n986), .B2(n1024), .C1(n954), .C2(n1021), .A(n2650), 
        .ZN(n2643) );
  OAI221_X1 U1218 ( .B1(n858), .B2(n1036), .C1(n826), .C2(n1033), .A(n2649), 
        .ZN(n2644) );
  OAI221_X1 U1219 ( .B1(n666), .B2(n1048), .C1(n634), .C2(n1045), .A(n2648), 
        .ZN(n2645) );
  NOR4_X1 U1220 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(n2625)
         );
  OAI221_X1 U1221 ( .B1(n985), .B2(n1024), .C1(n953), .C2(n1021), .A(n2633), 
        .ZN(n2626) );
  OAI221_X1 U1222 ( .B1(n857), .B2(n1036), .C1(n825), .C2(n1033), .A(n2632), 
        .ZN(n2627) );
  OAI221_X1 U1223 ( .B1(n665), .B2(n1048), .C1(n633), .C2(n1045), .A(n2631), 
        .ZN(n2628) );
  NOR4_X1 U1224 ( .A1(n2609), .A2(n2610), .A3(n2611), .A4(n2612), .ZN(n2608)
         );
  OAI221_X1 U1225 ( .B1(n984), .B2(n1024), .C1(n952), .C2(n1021), .A(n2616), 
        .ZN(n2609) );
  OAI221_X1 U1226 ( .B1(n856), .B2(n1036), .C1(n824), .C2(n1033), .A(n2615), 
        .ZN(n2610) );
  OAI221_X1 U1227 ( .B1(n664), .B2(n1048), .C1(n632), .C2(n1045), .A(n2614), 
        .ZN(n2611) );
  NOR4_X1 U1228 ( .A1(n2592), .A2(n2593), .A3(n2594), .A4(n2595), .ZN(n2591)
         );
  OAI221_X1 U1229 ( .B1(n983), .B2(n1024), .C1(n951), .C2(n1021), .A(n2599), 
        .ZN(n2592) );
  OAI221_X1 U1230 ( .B1(n855), .B2(n1036), .C1(n823), .C2(n1033), .A(n2598), 
        .ZN(n2593) );
  OAI221_X1 U1231 ( .B1(n663), .B2(n1048), .C1(n631), .C2(n1045), .A(n2597), 
        .ZN(n2594) );
  NOR4_X1 U1232 ( .A1(n2575), .A2(n2576), .A3(n2577), .A4(n2578), .ZN(n2574)
         );
  OAI221_X1 U1233 ( .B1(n982), .B2(n1024), .C1(n950), .C2(n1021), .A(n2582), 
        .ZN(n2575) );
  OAI221_X1 U1234 ( .B1(n854), .B2(n1036), .C1(n822), .C2(n1033), .A(n2581), 
        .ZN(n2576) );
  OAI221_X1 U1235 ( .B1(n662), .B2(n1048), .C1(n630), .C2(n1045), .A(n2580), 
        .ZN(n2577) );
  NOR4_X1 U1236 ( .A1(n2558), .A2(n2559), .A3(n2560), .A4(n2561), .ZN(n2557)
         );
  OAI221_X1 U1237 ( .B1(n981), .B2(n1025), .C1(n949), .C2(n1022), .A(n2565), 
        .ZN(n2558) );
  OAI221_X1 U1238 ( .B1(n853), .B2(n1037), .C1(n821), .C2(n1034), .A(n2564), 
        .ZN(n2559) );
  OAI221_X1 U1239 ( .B1(n661), .B2(n1049), .C1(n629), .C2(n1046), .A(n2563), 
        .ZN(n2560) );
  NOR4_X1 U1240 ( .A1(n2541), .A2(n2542), .A3(n2543), .A4(n2544), .ZN(n2540)
         );
  OAI221_X1 U1241 ( .B1(n980), .B2(n1025), .C1(n948), .C2(n1022), .A(n2548), 
        .ZN(n2541) );
  OAI221_X1 U1242 ( .B1(n852), .B2(n1037), .C1(n820), .C2(n1034), .A(n2547), 
        .ZN(n2542) );
  OAI221_X1 U1243 ( .B1(n660), .B2(n1049), .C1(n628), .C2(n1046), .A(n2546), 
        .ZN(n2543) );
  NOR4_X1 U1244 ( .A1(n2524), .A2(n2525), .A3(n2526), .A4(n2527), .ZN(n2523)
         );
  OAI221_X1 U1245 ( .B1(n979), .B2(n1025), .C1(n947), .C2(n1022), .A(n2531), 
        .ZN(n2524) );
  OAI221_X1 U1246 ( .B1(n851), .B2(n1037), .C1(n819), .C2(n1034), .A(n2530), 
        .ZN(n2525) );
  OAI221_X1 U1247 ( .B1(n659), .B2(n1049), .C1(n627), .C2(n1046), .A(n2529), 
        .ZN(n2526) );
  NOR4_X1 U1248 ( .A1(n2507), .A2(n2508), .A3(n2509), .A4(n2510), .ZN(n2506)
         );
  OAI221_X1 U1249 ( .B1(n978), .B2(n1025), .C1(n946), .C2(n1022), .A(n2514), 
        .ZN(n2507) );
  OAI221_X1 U1250 ( .B1(n850), .B2(n1037), .C1(n818), .C2(n1034), .A(n2513), 
        .ZN(n2508) );
  OAI221_X1 U1251 ( .B1(n658), .B2(n1049), .C1(n626), .C2(n1046), .A(n2512), 
        .ZN(n2509) );
  NOR4_X1 U1252 ( .A1(n2490), .A2(n2491), .A3(n2492), .A4(n2493), .ZN(n2489)
         );
  OAI221_X1 U1253 ( .B1(n977), .B2(n1025), .C1(n945), .C2(n1022), .A(n2497), 
        .ZN(n2490) );
  OAI221_X1 U1254 ( .B1(n849), .B2(n1037), .C1(n817), .C2(n1034), .A(n2496), 
        .ZN(n2491) );
  OAI221_X1 U1255 ( .B1(n657), .B2(n1049), .C1(n625), .C2(n1046), .A(n2495), 
        .ZN(n2492) );
  NOR4_X1 U1256 ( .A1(n2473), .A2(n2474), .A3(n2475), .A4(n2476), .ZN(n2472)
         );
  OAI221_X1 U1257 ( .B1(n976), .B2(n1025), .C1(n944), .C2(n1022), .A(n2480), 
        .ZN(n2473) );
  OAI221_X1 U1258 ( .B1(n848), .B2(n1037), .C1(n816), .C2(n1034), .A(n2479), 
        .ZN(n2474) );
  OAI221_X1 U1259 ( .B1(n656), .B2(n1049), .C1(n624), .C2(n1046), .A(n2478), 
        .ZN(n2475) );
  NOR4_X1 U1260 ( .A1(n2456), .A2(n2457), .A3(n2458), .A4(n2459), .ZN(n2455)
         );
  OAI221_X1 U1261 ( .B1(n975), .B2(n1025), .C1(n943), .C2(n1022), .A(n2463), 
        .ZN(n2456) );
  OAI221_X1 U1262 ( .B1(n847), .B2(n1037), .C1(n815), .C2(n1034), .A(n2462), 
        .ZN(n2457) );
  OAI221_X1 U1263 ( .B1(n655), .B2(n1049), .C1(n623), .C2(n1046), .A(n2461), 
        .ZN(n2458) );
  NOR4_X1 U1264 ( .A1(n2439), .A2(n2440), .A3(n2441), .A4(n2442), .ZN(n2438)
         );
  OAI221_X1 U1265 ( .B1(n974), .B2(n1025), .C1(n942), .C2(n1022), .A(n2446), 
        .ZN(n2439) );
  OAI221_X1 U1266 ( .B1(n846), .B2(n1037), .C1(n814), .C2(n1034), .A(n2445), 
        .ZN(n2440) );
  OAI221_X1 U1267 ( .B1(n654), .B2(n1049), .C1(n622), .C2(n1046), .A(n2444), 
        .ZN(n2441) );
  NOR4_X1 U1268 ( .A1(n2422), .A2(n2423), .A3(n2424), .A4(n2425), .ZN(n2421)
         );
  OAI221_X1 U1269 ( .B1(n973), .B2(n1025), .C1(n941), .C2(n1022), .A(n2429), 
        .ZN(n2422) );
  OAI221_X1 U1270 ( .B1(n845), .B2(n1037), .C1(n813), .C2(n1034), .A(n2428), 
        .ZN(n2423) );
  OAI221_X1 U1271 ( .B1(n653), .B2(n1049), .C1(n621), .C2(n1046), .A(n2427), 
        .ZN(n2424) );
  NOR4_X1 U1272 ( .A1(n2405), .A2(n2406), .A3(n2407), .A4(n2408), .ZN(n2404)
         );
  OAI221_X1 U1273 ( .B1(n972), .B2(n1025), .C1(n940), .C2(n1022), .A(n2412), 
        .ZN(n2405) );
  OAI221_X1 U1274 ( .B1(n844), .B2(n1037), .C1(n812), .C2(n1034), .A(n2411), 
        .ZN(n2406) );
  OAI221_X1 U1275 ( .B1(n652), .B2(n1049), .C1(n620), .C2(n1046), .A(n2410), 
        .ZN(n2407) );
  NOR4_X1 U1276 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2387)
         );
  OAI221_X1 U1277 ( .B1(n971), .B2(n1025), .C1(n939), .C2(n1022), .A(n2395), 
        .ZN(n2388) );
  OAI221_X1 U1278 ( .B1(n843), .B2(n1037), .C1(n811), .C2(n1034), .A(n2394), 
        .ZN(n2389) );
  OAI221_X1 U1279 ( .B1(n651), .B2(n1049), .C1(n619), .C2(n1046), .A(n2393), 
        .ZN(n2390) );
  OAI221_X1 U1280 ( .B1(n544), .B2(n3334), .C1(n512), .C2(n3331), .A(n2158), 
        .ZN(n2157) );
  AOI22_X1 U1281 ( .A1(n3328), .A2(\registers[19][0] ), .B1(n3325), .B2(
        \registers[18][0] ), .ZN(n2158) );
  OAI221_X1 U1282 ( .B1(n543), .B2(n3334), .C1(n511), .C2(n3331), .A(n2141), 
        .ZN(n2140) );
  AOI22_X1 U1283 ( .A1(n3328), .A2(\registers[19][1] ), .B1(n3325), .B2(
        \registers[18][1] ), .ZN(n2141) );
  OAI221_X1 U1284 ( .B1(n542), .B2(n3334), .C1(n510), .C2(n3331), .A(n2124), 
        .ZN(n2123) );
  AOI22_X1 U1285 ( .A1(n3328), .A2(\registers[19][2] ), .B1(n3325), .B2(
        \registers[18][2] ), .ZN(n2124) );
  OAI221_X1 U1286 ( .B1(n541), .B2(n3334), .C1(n509), .C2(n3331), .A(n2107), 
        .ZN(n2106) );
  AOI22_X1 U1287 ( .A1(n3328), .A2(\registers[19][3] ), .B1(n3325), .B2(
        \registers[18][3] ), .ZN(n2107) );
  OAI221_X1 U1288 ( .B1(n540), .B2(n3334), .C1(n508), .C2(n3331), .A(n2090), 
        .ZN(n2089) );
  AOI22_X1 U1289 ( .A1(n3328), .A2(\registers[19][4] ), .B1(n3325), .B2(
        \registers[18][4] ), .ZN(n2090) );
  OAI221_X1 U1290 ( .B1(n539), .B2(n3334), .C1(n507), .C2(n3331), .A(n2073), 
        .ZN(n2072) );
  AOI22_X1 U1291 ( .A1(n3328), .A2(\registers[19][5] ), .B1(n3325), .B2(
        \registers[18][5] ), .ZN(n2073) );
  OAI221_X1 U1292 ( .B1(n538), .B2(n3334), .C1(n506), .C2(n3331), .A(n2056), 
        .ZN(n2055) );
  AOI22_X1 U1293 ( .A1(n3328), .A2(\registers[19][6] ), .B1(n3325), .B2(
        \registers[18][6] ), .ZN(n2056) );
  OAI221_X1 U1294 ( .B1(n537), .B2(n3334), .C1(n505), .C2(n3331), .A(n2039), 
        .ZN(n2038) );
  AOI22_X1 U1295 ( .A1(n3328), .A2(\registers[19][7] ), .B1(n3325), .B2(
        \registers[18][7] ), .ZN(n2039) );
  OAI221_X1 U1296 ( .B1(n536), .B2(n3334), .C1(n504), .C2(n3331), .A(n2022), 
        .ZN(n2021) );
  AOI22_X1 U1297 ( .A1(n3328), .A2(\registers[19][8] ), .B1(n3325), .B2(
        \registers[18][8] ), .ZN(n2022) );
  OAI221_X1 U1298 ( .B1(n535), .B2(n3334), .C1(n503), .C2(n3331), .A(n2005), 
        .ZN(n2004) );
  AOI22_X1 U1299 ( .A1(n3328), .A2(\registers[19][9] ), .B1(n3325), .B2(
        \registers[18][9] ), .ZN(n2005) );
  OAI221_X1 U1300 ( .B1(n534), .B2(n3334), .C1(n502), .C2(n3331), .A(n1988), 
        .ZN(n1987) );
  AOI22_X1 U1301 ( .A1(n3328), .A2(\registers[19][10] ), .B1(n3325), .B2(
        \registers[18][10] ), .ZN(n1988) );
  OAI221_X1 U1302 ( .B1(n544), .B2(n1060), .C1(n512), .C2(n1057), .A(n2749), 
        .ZN(n2748) );
  AOI22_X1 U1303 ( .A1(n1054), .A2(\registers[19][0] ), .B1(n1051), .B2(
        \registers[18][0] ), .ZN(n2749) );
  OAI221_X1 U1304 ( .B1(n543), .B2(n1060), .C1(n511), .C2(n1057), .A(n2732), 
        .ZN(n2731) );
  AOI22_X1 U1305 ( .A1(n1054), .A2(\registers[19][1] ), .B1(n1051), .B2(
        \registers[18][1] ), .ZN(n2732) );
  OAI221_X1 U1306 ( .B1(n542), .B2(n1060), .C1(n510), .C2(n1057), .A(n2715), 
        .ZN(n2714) );
  AOI22_X1 U1307 ( .A1(n1054), .A2(\registers[19][2] ), .B1(n1051), .B2(
        \registers[18][2] ), .ZN(n2715) );
  OAI221_X1 U1308 ( .B1(n541), .B2(n1060), .C1(n509), .C2(n1057), .A(n2698), 
        .ZN(n2697) );
  AOI22_X1 U1309 ( .A1(n1054), .A2(\registers[19][3] ), .B1(n1051), .B2(
        \registers[18][3] ), .ZN(n2698) );
  OAI221_X1 U1310 ( .B1(n540), .B2(n1060), .C1(n508), .C2(n1057), .A(n2681), 
        .ZN(n2680) );
  AOI22_X1 U1311 ( .A1(n1054), .A2(\registers[19][4] ), .B1(n1051), .B2(
        \registers[18][4] ), .ZN(n2681) );
  OAI221_X1 U1312 ( .B1(n539), .B2(n1060), .C1(n507), .C2(n1057), .A(n2664), 
        .ZN(n2663) );
  AOI22_X1 U1313 ( .A1(n1054), .A2(\registers[19][5] ), .B1(n1051), .B2(
        \registers[18][5] ), .ZN(n2664) );
  OAI221_X1 U1314 ( .B1(n538), .B2(n1060), .C1(n506), .C2(n1057), .A(n2647), 
        .ZN(n2646) );
  AOI22_X1 U1315 ( .A1(n1054), .A2(\registers[19][6] ), .B1(n1051), .B2(
        \registers[18][6] ), .ZN(n2647) );
  OAI221_X1 U1316 ( .B1(n537), .B2(n1060), .C1(n505), .C2(n1057), .A(n2630), 
        .ZN(n2629) );
  AOI22_X1 U1317 ( .A1(n1054), .A2(\registers[19][7] ), .B1(n1051), .B2(
        \registers[18][7] ), .ZN(n2630) );
  OAI221_X1 U1318 ( .B1(n536), .B2(n1060), .C1(n504), .C2(n1057), .A(n2613), 
        .ZN(n2612) );
  AOI22_X1 U1319 ( .A1(n1054), .A2(\registers[19][8] ), .B1(n1051), .B2(
        \registers[18][8] ), .ZN(n2613) );
  OAI221_X1 U1320 ( .B1(n535), .B2(n1060), .C1(n503), .C2(n1057), .A(n2596), 
        .ZN(n2595) );
  AOI22_X1 U1321 ( .A1(n1054), .A2(\registers[19][9] ), .B1(n1051), .B2(
        \registers[18][9] ), .ZN(n2596) );
  OAI221_X1 U1322 ( .B1(n534), .B2(n1060), .C1(n502), .C2(n1057), .A(n2579), 
        .ZN(n2578) );
  AOI22_X1 U1323 ( .A1(n1054), .A2(\registers[19][10] ), .B1(n1051), .B2(
        \registers[18][10] ), .ZN(n2579) );
  OAI221_X1 U1324 ( .B1(n522), .B2(n3336), .C1(n490), .C2(n3333), .A(n1784), 
        .ZN(n1783) );
  AOI22_X1 U1325 ( .A1(n3330), .A2(\registers[19][22] ), .B1(n3327), .B2(
        \registers[18][22] ), .ZN(n1784) );
  OAI221_X1 U1326 ( .B1(n521), .B2(n3336), .C1(n489), .C2(n3333), .A(n1767), 
        .ZN(n1766) );
  AOI22_X1 U1327 ( .A1(n3330), .A2(\registers[19][23] ), .B1(n3327), .B2(
        \registers[18][23] ), .ZN(n1767) );
  OAI221_X1 U1328 ( .B1(n520), .B2(n3336), .C1(n488), .C2(n3333), .A(n1750), 
        .ZN(n1749) );
  AOI22_X1 U1329 ( .A1(n3330), .A2(\registers[19][24] ), .B1(n3327), .B2(
        \registers[18][24] ), .ZN(n1750) );
  OAI221_X1 U1330 ( .B1(n519), .B2(n3336), .C1(n487), .C2(n3333), .A(n1733), 
        .ZN(n1732) );
  AOI22_X1 U1331 ( .A1(n3330), .A2(\registers[19][25] ), .B1(n3327), .B2(
        \registers[18][25] ), .ZN(n1733) );
  OAI221_X1 U1332 ( .B1(n518), .B2(n3336), .C1(n486), .C2(n3333), .A(n1716), 
        .ZN(n1715) );
  AOI22_X1 U1333 ( .A1(n3330), .A2(\registers[19][26] ), .B1(n3327), .B2(
        \registers[18][26] ), .ZN(n1716) );
  OAI221_X1 U1334 ( .B1(n517), .B2(n3336), .C1(n485), .C2(n3333), .A(n1699), 
        .ZN(n1698) );
  AOI22_X1 U1335 ( .A1(n3330), .A2(\registers[19][27] ), .B1(n3327), .B2(
        \registers[18][27] ), .ZN(n1699) );
  OAI221_X1 U1336 ( .B1(n516), .B2(n3336), .C1(n484), .C2(n3333), .A(n1682), 
        .ZN(n1681) );
  AOI22_X1 U1337 ( .A1(n3330), .A2(\registers[19][28] ), .B1(n3327), .B2(
        \registers[18][28] ), .ZN(n1682) );
  OAI221_X1 U1338 ( .B1(n515), .B2(n3336), .C1(n483), .C2(n3333), .A(n1665), 
        .ZN(n1664) );
  AOI22_X1 U1339 ( .A1(n3330), .A2(\registers[19][29] ), .B1(n3327), .B2(
        \registers[18][29] ), .ZN(n1665) );
  OAI221_X1 U1340 ( .B1(n514), .B2(n3336), .C1(n482), .C2(n3333), .A(n1648), 
        .ZN(n1647) );
  AOI22_X1 U1341 ( .A1(n3330), .A2(\registers[19][30] ), .B1(n3327), .B2(
        \registers[18][30] ), .ZN(n1648) );
  OAI221_X1 U1342 ( .B1(n513), .B2(n3336), .C1(n481), .C2(n3333), .A(n1602), 
        .ZN(n1599) );
  AOI22_X1 U1343 ( .A1(n3330), .A2(\registers[19][31] ), .B1(n3327), .B2(
        \registers[18][31] ), .ZN(n1602) );
  OAI221_X1 U1344 ( .B1(n522), .B2(n1062), .C1(n490), .C2(n1059), .A(n2375), 
        .ZN(n2374) );
  AOI22_X1 U1345 ( .A1(n1056), .A2(\registers[19][22] ), .B1(n1053), .B2(
        \registers[18][22] ), .ZN(n2375) );
  OAI221_X1 U1346 ( .B1(n521), .B2(n1062), .C1(n489), .C2(n1059), .A(n2358), 
        .ZN(n2357) );
  AOI22_X1 U1347 ( .A1(n1056), .A2(\registers[19][23] ), .B1(n1053), .B2(
        \registers[18][23] ), .ZN(n2358) );
  OAI221_X1 U1348 ( .B1(n520), .B2(n1062), .C1(n488), .C2(n1059), .A(n2341), 
        .ZN(n2340) );
  AOI22_X1 U1349 ( .A1(n1056), .A2(\registers[19][24] ), .B1(n1053), .B2(
        \registers[18][24] ), .ZN(n2341) );
  OAI221_X1 U1350 ( .B1(n519), .B2(n1062), .C1(n487), .C2(n1059), .A(n2324), 
        .ZN(n2323) );
  AOI22_X1 U1351 ( .A1(n1056), .A2(\registers[19][25] ), .B1(n1053), .B2(
        \registers[18][25] ), .ZN(n2324) );
  OAI221_X1 U1352 ( .B1(n518), .B2(n1062), .C1(n486), .C2(n1059), .A(n2307), 
        .ZN(n2306) );
  AOI22_X1 U1353 ( .A1(n1056), .A2(\registers[19][26] ), .B1(n1053), .B2(
        \registers[18][26] ), .ZN(n2307) );
  OAI221_X1 U1354 ( .B1(n517), .B2(n1062), .C1(n485), .C2(n1059), .A(n2290), 
        .ZN(n2289) );
  AOI22_X1 U1355 ( .A1(n1056), .A2(\registers[19][27] ), .B1(n1053), .B2(
        \registers[18][27] ), .ZN(n2290) );
  OAI221_X1 U1356 ( .B1(n516), .B2(n1062), .C1(n484), .C2(n1059), .A(n2273), 
        .ZN(n2272) );
  AOI22_X1 U1357 ( .A1(n1056), .A2(\registers[19][28] ), .B1(n1053), .B2(
        \registers[18][28] ), .ZN(n2273) );
  OAI221_X1 U1358 ( .B1(n515), .B2(n1062), .C1(n483), .C2(n1059), .A(n2256), 
        .ZN(n2255) );
  AOI22_X1 U1359 ( .A1(n1056), .A2(\registers[19][29] ), .B1(n1053), .B2(
        \registers[18][29] ), .ZN(n2256) );
  OAI221_X1 U1360 ( .B1(n514), .B2(n1062), .C1(n482), .C2(n1059), .A(n2239), 
        .ZN(n2238) );
  AOI22_X1 U1361 ( .A1(n1056), .A2(\registers[19][30] ), .B1(n1053), .B2(
        \registers[18][30] ), .ZN(n2239) );
  OAI221_X1 U1362 ( .B1(n513), .B2(n1062), .C1(n481), .C2(n1059), .A(n2193), 
        .ZN(n2190) );
  AOI22_X1 U1363 ( .A1(n1056), .A2(\registers[19][31] ), .B1(n1053), .B2(
        \registers[18][31] ), .ZN(n2193) );
  OAI221_X1 U1364 ( .B1(n533), .B2(n3335), .C1(n501), .C2(n3332), .A(n1971), 
        .ZN(n1970) );
  AOI22_X1 U1365 ( .A1(n3329), .A2(\registers[19][11] ), .B1(n3326), .B2(
        \registers[18][11] ), .ZN(n1971) );
  OAI221_X1 U1366 ( .B1(n532), .B2(n3335), .C1(n500), .C2(n3332), .A(n1954), 
        .ZN(n1953) );
  AOI22_X1 U1367 ( .A1(n3329), .A2(\registers[19][12] ), .B1(n3326), .B2(
        \registers[18][12] ), .ZN(n1954) );
  OAI221_X1 U1368 ( .B1(n531), .B2(n3335), .C1(n499), .C2(n3332), .A(n1937), 
        .ZN(n1936) );
  AOI22_X1 U1369 ( .A1(n3329), .A2(\registers[19][13] ), .B1(n3326), .B2(
        \registers[18][13] ), .ZN(n1937) );
  OAI221_X1 U1370 ( .B1(n530), .B2(n3335), .C1(n498), .C2(n3332), .A(n1920), 
        .ZN(n1919) );
  AOI22_X1 U1371 ( .A1(n3329), .A2(\registers[19][14] ), .B1(n3326), .B2(
        \registers[18][14] ), .ZN(n1920) );
  OAI221_X1 U1372 ( .B1(n529), .B2(n3335), .C1(n497), .C2(n3332), .A(n1903), 
        .ZN(n1902) );
  AOI22_X1 U1373 ( .A1(n3329), .A2(\registers[19][15] ), .B1(n3326), .B2(
        \registers[18][15] ), .ZN(n1903) );
  OAI221_X1 U1374 ( .B1(n528), .B2(n3335), .C1(n496), .C2(n3332), .A(n1886), 
        .ZN(n1885) );
  AOI22_X1 U1375 ( .A1(n3329), .A2(\registers[19][16] ), .B1(n3326), .B2(
        \registers[18][16] ), .ZN(n1886) );
  OAI221_X1 U1376 ( .B1(n527), .B2(n3335), .C1(n495), .C2(n3332), .A(n1869), 
        .ZN(n1868) );
  AOI22_X1 U1377 ( .A1(n3329), .A2(\registers[19][17] ), .B1(n3326), .B2(
        \registers[18][17] ), .ZN(n1869) );
  OAI221_X1 U1378 ( .B1(n526), .B2(n3335), .C1(n494), .C2(n3332), .A(n1852), 
        .ZN(n1851) );
  AOI22_X1 U1379 ( .A1(n3329), .A2(\registers[19][18] ), .B1(n3326), .B2(
        \registers[18][18] ), .ZN(n1852) );
  OAI221_X1 U1380 ( .B1(n525), .B2(n3335), .C1(n493), .C2(n3332), .A(n1835), 
        .ZN(n1834) );
  AOI22_X1 U1381 ( .A1(n3329), .A2(\registers[19][19] ), .B1(n3326), .B2(
        \registers[18][19] ), .ZN(n1835) );
  OAI221_X1 U1382 ( .B1(n524), .B2(n3335), .C1(n492), .C2(n3332), .A(n1818), 
        .ZN(n1817) );
  AOI22_X1 U1383 ( .A1(n3329), .A2(\registers[19][20] ), .B1(n3326), .B2(
        \registers[18][20] ), .ZN(n1818) );
  OAI221_X1 U1384 ( .B1(n523), .B2(n3335), .C1(n491), .C2(n3332), .A(n1801), 
        .ZN(n1800) );
  AOI22_X1 U1385 ( .A1(n3329), .A2(\registers[19][21] ), .B1(n3326), .B2(
        \registers[18][21] ), .ZN(n1801) );
  OAI221_X1 U1386 ( .B1(n533), .B2(n1061), .C1(n501), .C2(n1058), .A(n2562), 
        .ZN(n2561) );
  AOI22_X1 U1387 ( .A1(n1055), .A2(\registers[19][11] ), .B1(n1052), .B2(
        \registers[18][11] ), .ZN(n2562) );
  OAI221_X1 U1388 ( .B1(n532), .B2(n1061), .C1(n500), .C2(n1058), .A(n2545), 
        .ZN(n2544) );
  AOI22_X1 U1389 ( .A1(n1055), .A2(\registers[19][12] ), .B1(n1052), .B2(
        \registers[18][12] ), .ZN(n2545) );
  OAI221_X1 U1390 ( .B1(n531), .B2(n1061), .C1(n499), .C2(n1058), .A(n2528), 
        .ZN(n2527) );
  AOI22_X1 U1391 ( .A1(n1055), .A2(\registers[19][13] ), .B1(n1052), .B2(
        \registers[18][13] ), .ZN(n2528) );
  OAI221_X1 U1392 ( .B1(n530), .B2(n1061), .C1(n498), .C2(n1058), .A(n2511), 
        .ZN(n2510) );
  AOI22_X1 U1393 ( .A1(n1055), .A2(\registers[19][14] ), .B1(n1052), .B2(
        \registers[18][14] ), .ZN(n2511) );
  OAI221_X1 U1394 ( .B1(n529), .B2(n1061), .C1(n497), .C2(n1058), .A(n2494), 
        .ZN(n2493) );
  AOI22_X1 U1395 ( .A1(n1055), .A2(\registers[19][15] ), .B1(n1052), .B2(
        \registers[18][15] ), .ZN(n2494) );
  OAI221_X1 U1396 ( .B1(n528), .B2(n1061), .C1(n496), .C2(n1058), .A(n2477), 
        .ZN(n2476) );
  AOI22_X1 U1397 ( .A1(n1055), .A2(\registers[19][16] ), .B1(n1052), .B2(
        \registers[18][16] ), .ZN(n2477) );
  OAI221_X1 U1398 ( .B1(n527), .B2(n1061), .C1(n495), .C2(n1058), .A(n2460), 
        .ZN(n2459) );
  AOI22_X1 U1399 ( .A1(n1055), .A2(\registers[19][17] ), .B1(n1052), .B2(
        \registers[18][17] ), .ZN(n2460) );
  OAI221_X1 U1400 ( .B1(n526), .B2(n1061), .C1(n494), .C2(n1058), .A(n2443), 
        .ZN(n2442) );
  AOI22_X1 U1401 ( .A1(n1055), .A2(\registers[19][18] ), .B1(n1052), .B2(
        \registers[18][18] ), .ZN(n2443) );
  OAI221_X1 U1402 ( .B1(n525), .B2(n1061), .C1(n493), .C2(n1058), .A(n2426), 
        .ZN(n2425) );
  AOI22_X1 U1403 ( .A1(n1055), .A2(\registers[19][19] ), .B1(n1052), .B2(
        \registers[18][19] ), .ZN(n2426) );
  OAI221_X1 U1404 ( .B1(n524), .B2(n1061), .C1(n492), .C2(n1058), .A(n2409), 
        .ZN(n2408) );
  AOI22_X1 U1405 ( .A1(n1055), .A2(\registers[19][20] ), .B1(n1052), .B2(
        \registers[18][20] ), .ZN(n2409) );
  OAI221_X1 U1406 ( .B1(n523), .B2(n1061), .C1(n491), .C2(n1058), .A(n2392), 
        .ZN(n2391) );
  AOI22_X1 U1407 ( .A1(n1055), .A2(\registers[19][21] ), .B1(n1052), .B2(
        \registers[18][21] ), .ZN(n2392) );
  OAI221_X1 U1408 ( .B1(n160), .B2(n1424), .C1(n128), .C2(n1420), .A(n2176), 
        .ZN(n2172) );
  AOI22_X1 U1409 ( .A1(n1399), .A2(\registers[7][0] ), .B1(n1357), .B2(
        \registers[6][0] ), .ZN(n2176) );
  OAI221_X1 U1410 ( .B1(n159), .B2(n1424), .C1(n127), .C2(n1420), .A(n2147), 
        .ZN(n2145) );
  AOI22_X1 U1411 ( .A1(n1399), .A2(\registers[7][1] ), .B1(n1357), .B2(
        \registers[6][1] ), .ZN(n2147) );
  OAI221_X1 U1412 ( .B1(n158), .B2(n1424), .C1(n126), .C2(n1420), .A(n2130), 
        .ZN(n2128) );
  AOI22_X1 U1413 ( .A1(n1399), .A2(\registers[7][2] ), .B1(n1357), .B2(
        \registers[6][2] ), .ZN(n2130) );
  OAI221_X1 U1414 ( .B1(n157), .B2(n1424), .C1(n125), .C2(n1420), .A(n2113), 
        .ZN(n2111) );
  AOI22_X1 U1415 ( .A1(n1399), .A2(\registers[7][3] ), .B1(n1357), .B2(
        \registers[6][3] ), .ZN(n2113) );
  OAI221_X1 U1416 ( .B1(n156), .B2(n1424), .C1(n124), .C2(n1420), .A(n2096), 
        .ZN(n2094) );
  AOI22_X1 U1417 ( .A1(n1399), .A2(\registers[7][4] ), .B1(n1357), .B2(
        \registers[6][4] ), .ZN(n2096) );
  OAI221_X1 U1418 ( .B1(n155), .B2(n1424), .C1(n123), .C2(n1420), .A(n2079), 
        .ZN(n2077) );
  AOI22_X1 U1419 ( .A1(n1399), .A2(\registers[7][5] ), .B1(n1357), .B2(
        \registers[6][5] ), .ZN(n2079) );
  OAI221_X1 U1420 ( .B1(n154), .B2(n1424), .C1(n122), .C2(n1420), .A(n2062), 
        .ZN(n2060) );
  AOI22_X1 U1421 ( .A1(n1399), .A2(\registers[7][6] ), .B1(n1357), .B2(
        \registers[6][6] ), .ZN(n2062) );
  OAI221_X1 U1422 ( .B1(n153), .B2(n1424), .C1(n121), .C2(n1420), .A(n2045), 
        .ZN(n2043) );
  AOI22_X1 U1423 ( .A1(n1399), .A2(\registers[7][7] ), .B1(n1357), .B2(
        \registers[6][7] ), .ZN(n2045) );
  OAI221_X1 U1424 ( .B1(n152), .B2(n1424), .C1(n120), .C2(n1420), .A(n2028), 
        .ZN(n2026) );
  AOI22_X1 U1425 ( .A1(n1399), .A2(\registers[7][8] ), .B1(n1357), .B2(
        \registers[6][8] ), .ZN(n2028) );
  OAI221_X1 U1426 ( .B1(n151), .B2(n1424), .C1(n119), .C2(n1420), .A(n2011), 
        .ZN(n2009) );
  AOI22_X1 U1427 ( .A1(n1399), .A2(\registers[7][9] ), .B1(n1357), .B2(
        \registers[6][9] ), .ZN(n2011) );
  OAI221_X1 U1428 ( .B1(n150), .B2(n1424), .C1(n118), .C2(n1420), .A(n1994), 
        .ZN(n1992) );
  AOI22_X1 U1429 ( .A1(n1399), .A2(\registers[7][10] ), .B1(n1357), .B2(
        \registers[6][10] ), .ZN(n1994) );
  OAI221_X1 U1430 ( .B1(n160), .B2(n1003), .C1(n128), .C2(n1000), .A(n2767), 
        .ZN(n2763) );
  AOI22_X1 U1431 ( .A1(n997), .A2(\registers[7][0] ), .B1(n994), .B2(
        \registers[6][0] ), .ZN(n2767) );
  OAI221_X1 U1432 ( .B1(n159), .B2(n1003), .C1(n127), .C2(n1000), .A(n2738), 
        .ZN(n2736) );
  AOI22_X1 U1433 ( .A1(n997), .A2(\registers[7][1] ), .B1(n994), .B2(
        \registers[6][1] ), .ZN(n2738) );
  OAI221_X1 U1434 ( .B1(n158), .B2(n1003), .C1(n126), .C2(n1000), .A(n2721), 
        .ZN(n2719) );
  AOI22_X1 U1435 ( .A1(n997), .A2(\registers[7][2] ), .B1(n994), .B2(
        \registers[6][2] ), .ZN(n2721) );
  OAI221_X1 U1436 ( .B1(n157), .B2(n1003), .C1(n125), .C2(n1000), .A(n2704), 
        .ZN(n2702) );
  AOI22_X1 U1437 ( .A1(n997), .A2(\registers[7][3] ), .B1(n994), .B2(
        \registers[6][3] ), .ZN(n2704) );
  OAI221_X1 U1438 ( .B1(n156), .B2(n1003), .C1(n124), .C2(n1000), .A(n2687), 
        .ZN(n2685) );
  AOI22_X1 U1439 ( .A1(n997), .A2(\registers[7][4] ), .B1(n994), .B2(
        \registers[6][4] ), .ZN(n2687) );
  OAI221_X1 U1440 ( .B1(n155), .B2(n1003), .C1(n123), .C2(n1000), .A(n2670), 
        .ZN(n2668) );
  AOI22_X1 U1441 ( .A1(n997), .A2(\registers[7][5] ), .B1(n994), .B2(
        \registers[6][5] ), .ZN(n2670) );
  OAI221_X1 U1442 ( .B1(n154), .B2(n1003), .C1(n122), .C2(n1000), .A(n2653), 
        .ZN(n2651) );
  AOI22_X1 U1443 ( .A1(n997), .A2(\registers[7][6] ), .B1(n994), .B2(
        \registers[6][6] ), .ZN(n2653) );
  OAI221_X1 U1444 ( .B1(n153), .B2(n1003), .C1(n121), .C2(n1000), .A(n2636), 
        .ZN(n2634) );
  AOI22_X1 U1445 ( .A1(n997), .A2(\registers[7][7] ), .B1(n994), .B2(
        \registers[6][7] ), .ZN(n2636) );
  OAI221_X1 U1446 ( .B1(n152), .B2(n1003), .C1(n120), .C2(n1000), .A(n2619), 
        .ZN(n2617) );
  AOI22_X1 U1447 ( .A1(n997), .A2(\registers[7][8] ), .B1(n994), .B2(
        \registers[6][8] ), .ZN(n2619) );
  OAI221_X1 U1448 ( .B1(n151), .B2(n1003), .C1(n119), .C2(n1000), .A(n2602), 
        .ZN(n2600) );
  AOI22_X1 U1449 ( .A1(n997), .A2(\registers[7][9] ), .B1(n994), .B2(
        \registers[6][9] ), .ZN(n2602) );
  OAI221_X1 U1450 ( .B1(n150), .B2(n1003), .C1(n118), .C2(n1000), .A(n2585), 
        .ZN(n2583) );
  AOI22_X1 U1451 ( .A1(n997), .A2(\registers[7][10] ), .B1(n994), .B2(
        \registers[6][10] ), .ZN(n2585) );
  OAI221_X1 U1452 ( .B1(n138), .B2(n1429), .C1(n106), .C2(n1422), .A(n1790), 
        .ZN(n1788) );
  AOI22_X1 U1453 ( .A1(n1404), .A2(\registers[7][22] ), .B1(n1387), .B2(
        \registers[6][22] ), .ZN(n1790) );
  OAI221_X1 U1454 ( .B1(n137), .B2(n1429), .C1(n105), .C2(n1422), .A(n1773), 
        .ZN(n1771) );
  AOI22_X1 U1455 ( .A1(n1404), .A2(\registers[7][23] ), .B1(n1387), .B2(
        \registers[6][23] ), .ZN(n1773) );
  OAI221_X1 U1456 ( .B1(n136), .B2(n1429), .C1(n104), .C2(n1422), .A(n1756), 
        .ZN(n1754) );
  AOI22_X1 U1457 ( .A1(n1404), .A2(\registers[7][24] ), .B1(n1387), .B2(
        \registers[6][24] ), .ZN(n1756) );
  OAI221_X1 U1458 ( .B1(n135), .B2(n1429), .C1(n103), .C2(n1422), .A(n1739), 
        .ZN(n1737) );
  AOI22_X1 U1459 ( .A1(n1404), .A2(\registers[7][25] ), .B1(n1387), .B2(
        \registers[6][25] ), .ZN(n1739) );
  OAI221_X1 U1460 ( .B1(n134), .B2(n1429), .C1(n102), .C2(n1422), .A(n1722), 
        .ZN(n1720) );
  AOI22_X1 U1461 ( .A1(n1404), .A2(\registers[7][26] ), .B1(n1387), .B2(
        \registers[6][26] ), .ZN(n1722) );
  OAI221_X1 U1462 ( .B1(n133), .B2(n1429), .C1(n101), .C2(n1422), .A(n1705), 
        .ZN(n1703) );
  AOI22_X1 U1463 ( .A1(n1404), .A2(\registers[7][27] ), .B1(n1387), .B2(
        \registers[6][27] ), .ZN(n1705) );
  OAI221_X1 U1464 ( .B1(n132), .B2(n1429), .C1(n100), .C2(n1422), .A(n1688), 
        .ZN(n1686) );
  AOI22_X1 U1465 ( .A1(n1404), .A2(\registers[7][28] ), .B1(n1387), .B2(
        \registers[6][28] ), .ZN(n1688) );
  OAI221_X1 U1466 ( .B1(n131), .B2(n1429), .C1(n99), .C2(n1422), .A(n1671), 
        .ZN(n1669) );
  AOI22_X1 U1467 ( .A1(n1404), .A2(\registers[7][29] ), .B1(n1387), .B2(
        \registers[6][29] ), .ZN(n1671) );
  OAI221_X1 U1468 ( .B1(n130), .B2(n1429), .C1(n98), .C2(n1422), .A(n1654), 
        .ZN(n1652) );
  AOI22_X1 U1469 ( .A1(n1404), .A2(\registers[7][30] ), .B1(n1387), .B2(
        \registers[6][30] ), .ZN(n1654) );
  OAI221_X1 U1470 ( .B1(n129), .B2(n1429), .C1(n97), .C2(n1422), .A(n1627), 
        .ZN(n1621) );
  AOI22_X1 U1471 ( .A1(n1404), .A2(\registers[7][31] ), .B1(n1387), .B2(
        \registers[6][31] ), .ZN(n1627) );
  OAI221_X1 U1472 ( .B1(n138), .B2(n1005), .C1(n106), .C2(n1002), .A(n2381), 
        .ZN(n2379) );
  AOI22_X1 U1473 ( .A1(n999), .A2(\registers[7][22] ), .B1(n996), .B2(
        \registers[6][22] ), .ZN(n2381) );
  OAI221_X1 U1474 ( .B1(n137), .B2(n1005), .C1(n105), .C2(n1002), .A(n2364), 
        .ZN(n2362) );
  AOI22_X1 U1475 ( .A1(n999), .A2(\registers[7][23] ), .B1(n996), .B2(
        \registers[6][23] ), .ZN(n2364) );
  OAI221_X1 U1476 ( .B1(n136), .B2(n1005), .C1(n104), .C2(n1002), .A(n2347), 
        .ZN(n2345) );
  AOI22_X1 U1477 ( .A1(n999), .A2(\registers[7][24] ), .B1(n996), .B2(
        \registers[6][24] ), .ZN(n2347) );
  OAI221_X1 U1478 ( .B1(n135), .B2(n1005), .C1(n103), .C2(n1002), .A(n2330), 
        .ZN(n2328) );
  AOI22_X1 U1479 ( .A1(n999), .A2(\registers[7][25] ), .B1(n996), .B2(
        \registers[6][25] ), .ZN(n2330) );
  OAI221_X1 U1480 ( .B1(n134), .B2(n1005), .C1(n102), .C2(n1002), .A(n2313), 
        .ZN(n2311) );
  AOI22_X1 U1481 ( .A1(n999), .A2(\registers[7][26] ), .B1(n996), .B2(
        \registers[6][26] ), .ZN(n2313) );
  OAI221_X1 U1482 ( .B1(n133), .B2(n1005), .C1(n101), .C2(n1002), .A(n2296), 
        .ZN(n2294) );
  AOI22_X1 U1483 ( .A1(n999), .A2(\registers[7][27] ), .B1(n996), .B2(
        \registers[6][27] ), .ZN(n2296) );
  OAI221_X1 U1484 ( .B1(n132), .B2(n1005), .C1(n100), .C2(n1002), .A(n2279), 
        .ZN(n2277) );
  AOI22_X1 U1485 ( .A1(n999), .A2(\registers[7][28] ), .B1(n996), .B2(
        \registers[6][28] ), .ZN(n2279) );
  OAI221_X1 U1486 ( .B1(n131), .B2(n1005), .C1(n99), .C2(n1002), .A(n2262), 
        .ZN(n2260) );
  AOI22_X1 U1487 ( .A1(n999), .A2(\registers[7][29] ), .B1(n996), .B2(
        \registers[6][29] ), .ZN(n2262) );
  OAI221_X1 U1488 ( .B1(n130), .B2(n1005), .C1(n98), .C2(n1002), .A(n2245), 
        .ZN(n2243) );
  AOI22_X1 U1489 ( .A1(n999), .A2(\registers[7][30] ), .B1(n996), .B2(
        \registers[6][30] ), .ZN(n2245) );
  OAI221_X1 U1490 ( .B1(n129), .B2(n1005), .C1(n97), .C2(n1002), .A(n2218), 
        .ZN(n2212) );
  AOI22_X1 U1491 ( .A1(n999), .A2(\registers[7][31] ), .B1(n996), .B2(
        \registers[6][31] ), .ZN(n2218) );
  OAI221_X1 U1492 ( .B1(n149), .B2(n1427), .C1(n117), .C2(n1421), .A(n1977), 
        .ZN(n1975) );
  AOI22_X1 U1493 ( .A1(n1403), .A2(\registers[7][11] ), .B1(n1367), .B2(
        \registers[6][11] ), .ZN(n1977) );
  OAI221_X1 U1494 ( .B1(n148), .B2(n1427), .C1(n116), .C2(n1421), .A(n1960), 
        .ZN(n1958) );
  AOI22_X1 U1495 ( .A1(n1403), .A2(\registers[7][12] ), .B1(n1367), .B2(
        \registers[6][12] ), .ZN(n1960) );
  OAI221_X1 U1496 ( .B1(n147), .B2(n1427), .C1(n115), .C2(n1421), .A(n1943), 
        .ZN(n1941) );
  AOI22_X1 U1497 ( .A1(n1403), .A2(\registers[7][13] ), .B1(n1367), .B2(
        \registers[6][13] ), .ZN(n1943) );
  OAI221_X1 U1498 ( .B1(n146), .B2(n1427), .C1(n114), .C2(n1421), .A(n1926), 
        .ZN(n1924) );
  AOI22_X1 U1499 ( .A1(n1403), .A2(\registers[7][14] ), .B1(n1367), .B2(
        \registers[6][14] ), .ZN(n1926) );
  OAI221_X1 U1500 ( .B1(n145), .B2(n1427), .C1(n113), .C2(n1421), .A(n1909), 
        .ZN(n1907) );
  AOI22_X1 U1501 ( .A1(n1403), .A2(\registers[7][15] ), .B1(n1367), .B2(
        \registers[6][15] ), .ZN(n1909) );
  OAI221_X1 U1502 ( .B1(n144), .B2(n1427), .C1(n112), .C2(n1421), .A(n1892), 
        .ZN(n1890) );
  AOI22_X1 U1503 ( .A1(n1403), .A2(\registers[7][16] ), .B1(n1367), .B2(
        \registers[6][16] ), .ZN(n1892) );
  OAI221_X1 U1504 ( .B1(n143), .B2(n1427), .C1(n111), .C2(n1421), .A(n1875), 
        .ZN(n1873) );
  AOI22_X1 U1505 ( .A1(n1403), .A2(\registers[7][17] ), .B1(n1367), .B2(
        \registers[6][17] ), .ZN(n1875) );
  OAI221_X1 U1506 ( .B1(n142), .B2(n1427), .C1(n110), .C2(n1421), .A(n1858), 
        .ZN(n1856) );
  AOI22_X1 U1507 ( .A1(n1403), .A2(\registers[7][18] ), .B1(n1367), .B2(
        \registers[6][18] ), .ZN(n1858) );
  OAI221_X1 U1508 ( .B1(n141), .B2(n1427), .C1(n109), .C2(n1421), .A(n1841), 
        .ZN(n1839) );
  AOI22_X1 U1509 ( .A1(n1403), .A2(\registers[7][19] ), .B1(n1367), .B2(
        \registers[6][19] ), .ZN(n1841) );
  OAI221_X1 U1510 ( .B1(n140), .B2(n1427), .C1(n108), .C2(n1421), .A(n1824), 
        .ZN(n1822) );
  AOI22_X1 U1511 ( .A1(n1403), .A2(\registers[7][20] ), .B1(n1367), .B2(
        \registers[6][20] ), .ZN(n1824) );
  OAI221_X1 U1512 ( .B1(n139), .B2(n1427), .C1(n107), .C2(n1421), .A(n1807), 
        .ZN(n1805) );
  AOI22_X1 U1513 ( .A1(n1403), .A2(\registers[7][21] ), .B1(n1367), .B2(
        \registers[6][21] ), .ZN(n1807) );
  OAI221_X1 U1514 ( .B1(n149), .B2(n1004), .C1(n117), .C2(n1001), .A(n2568), 
        .ZN(n2566) );
  AOI22_X1 U1515 ( .A1(n998), .A2(\registers[7][11] ), .B1(n995), .B2(
        \registers[6][11] ), .ZN(n2568) );
  OAI221_X1 U1516 ( .B1(n148), .B2(n1004), .C1(n116), .C2(n1001), .A(n2551), 
        .ZN(n2549) );
  AOI22_X1 U1517 ( .A1(n998), .A2(\registers[7][12] ), .B1(n995), .B2(
        \registers[6][12] ), .ZN(n2551) );
  OAI221_X1 U1518 ( .B1(n147), .B2(n1004), .C1(n115), .C2(n1001), .A(n2534), 
        .ZN(n2532) );
  AOI22_X1 U1519 ( .A1(n998), .A2(\registers[7][13] ), .B1(n995), .B2(
        \registers[6][13] ), .ZN(n2534) );
  OAI221_X1 U1520 ( .B1(n146), .B2(n1004), .C1(n114), .C2(n1001), .A(n2517), 
        .ZN(n2515) );
  AOI22_X1 U1521 ( .A1(n998), .A2(\registers[7][14] ), .B1(n995), .B2(
        \registers[6][14] ), .ZN(n2517) );
  OAI221_X1 U1522 ( .B1(n145), .B2(n1004), .C1(n113), .C2(n1001), .A(n2500), 
        .ZN(n2498) );
  AOI22_X1 U1523 ( .A1(n998), .A2(\registers[7][15] ), .B1(n995), .B2(
        \registers[6][15] ), .ZN(n2500) );
  OAI221_X1 U1524 ( .B1(n144), .B2(n1004), .C1(n112), .C2(n1001), .A(n2483), 
        .ZN(n2481) );
  AOI22_X1 U1525 ( .A1(n998), .A2(\registers[7][16] ), .B1(n995), .B2(
        \registers[6][16] ), .ZN(n2483) );
  OAI221_X1 U1526 ( .B1(n143), .B2(n1004), .C1(n111), .C2(n1001), .A(n2466), 
        .ZN(n2464) );
  AOI22_X1 U1527 ( .A1(n998), .A2(\registers[7][17] ), .B1(n995), .B2(
        \registers[6][17] ), .ZN(n2466) );
  OAI221_X1 U1528 ( .B1(n142), .B2(n1004), .C1(n110), .C2(n1001), .A(n2449), 
        .ZN(n2447) );
  AOI22_X1 U1529 ( .A1(n998), .A2(\registers[7][18] ), .B1(n995), .B2(
        \registers[6][18] ), .ZN(n2449) );
  OAI221_X1 U1530 ( .B1(n141), .B2(n1004), .C1(n109), .C2(n1001), .A(n2432), 
        .ZN(n2430) );
  AOI22_X1 U1531 ( .A1(n998), .A2(\registers[7][19] ), .B1(n995), .B2(
        \registers[6][19] ), .ZN(n2432) );
  OAI221_X1 U1532 ( .B1(n140), .B2(n1004), .C1(n108), .C2(n1001), .A(n2415), 
        .ZN(n2413) );
  AOI22_X1 U1533 ( .A1(n998), .A2(\registers[7][20] ), .B1(n995), .B2(
        \registers[6][20] ), .ZN(n2415) );
  OAI221_X1 U1534 ( .B1(n139), .B2(n1004), .C1(n107), .C2(n1001), .A(n2398), 
        .ZN(n2396) );
  AOI22_X1 U1535 ( .A1(n998), .A2(\registers[7][21] ), .B1(n995), .B2(
        \registers[6][21] ), .ZN(n2398) );
  AND2_X1 U1536 ( .A1(ADD_RD2[2]), .A2(n4178), .ZN(n2165) );
  AND2_X1 U1537 ( .A1(ADD_RD1[2]), .A2(n4175), .ZN(n2756) );
  AND2_X1 U1538 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n2164) );
  AND2_X1 U1539 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n2755) );
  OAI22_X1 U1540 ( .A1(n296), .A2(n1071), .B1(n328), .B2(n1065), .ZN(n1758) );
  OAI22_X1 U1541 ( .A1(n295), .A2(n1071), .B1(n327), .B2(n1065), .ZN(n1741) );
  OAI22_X1 U1542 ( .A1(n294), .A2(n1071), .B1(n326), .B2(n1065), .ZN(n1724) );
  OAI22_X1 U1543 ( .A1(n293), .A2(n1071), .B1(n325), .B2(n1065), .ZN(n1707) );
  OAI22_X1 U1544 ( .A1(n292), .A2(n1071), .B1(n324), .B2(n1065), .ZN(n1690) );
  OAI22_X1 U1545 ( .A1(n291), .A2(n1071), .B1(n323), .B2(n1065), .ZN(n1673) );
  OAI22_X1 U1546 ( .A1(n290), .A2(n1071), .B1(n322), .B2(n1065), .ZN(n1656) );
  OAI22_X1 U1547 ( .A1(n289), .A2(n1071), .B1(n321), .B2(n1065), .ZN(n1637) );
  OAI22_X1 U1548 ( .A1(n296), .A2(n911), .B1(n328), .B2(n908), .ZN(n2349) );
  OAI22_X1 U1549 ( .A1(n295), .A2(n911), .B1(n327), .B2(n908), .ZN(n2332) );
  OAI22_X1 U1550 ( .A1(n294), .A2(n911), .B1(n326), .B2(n908), .ZN(n2315) );
  OAI22_X1 U1551 ( .A1(n293), .A2(n911), .B1(n325), .B2(n908), .ZN(n2298) );
  OAI22_X1 U1552 ( .A1(n292), .A2(n911), .B1(n324), .B2(n908), .ZN(n2281) );
  OAI22_X1 U1553 ( .A1(n291), .A2(n911), .B1(n323), .B2(n908), .ZN(n2264) );
  OAI22_X1 U1554 ( .A1(n290), .A2(n911), .B1(n322), .B2(n908), .ZN(n2247) );
  OAI22_X1 U1555 ( .A1(n289), .A2(n911), .B1(n321), .B2(n908), .ZN(n2228) );
  OAI22_X1 U1556 ( .A1(n424), .A2(n1282), .B1(n456), .B2(n1266), .ZN(n1757) );
  OAI22_X1 U1557 ( .A1(n423), .A2(n1282), .B1(n455), .B2(n1266), .ZN(n1740) );
  OAI22_X1 U1558 ( .A1(n422), .A2(n1282), .B1(n454), .B2(n1266), .ZN(n1723) );
  OAI22_X1 U1559 ( .A1(n421), .A2(n1282), .B1(n453), .B2(n1266), .ZN(n1706) );
  OAI22_X1 U1560 ( .A1(n420), .A2(n1282), .B1(n452), .B2(n1266), .ZN(n1689) );
  OAI22_X1 U1561 ( .A1(n419), .A2(n1282), .B1(n451), .B2(n1266), .ZN(n1672) );
  OAI22_X1 U1562 ( .A1(n418), .A2(n1282), .B1(n450), .B2(n1266), .ZN(n1655) );
  OAI22_X1 U1563 ( .A1(n417), .A2(n1282), .B1(n449), .B2(n1266), .ZN(n1632) );
  OAI22_X1 U1564 ( .A1(n424), .A2(n923), .B1(n456), .B2(n920), .ZN(n2348) );
  OAI22_X1 U1565 ( .A1(n423), .A2(n923), .B1(n455), .B2(n920), .ZN(n2331) );
  OAI22_X1 U1566 ( .A1(n422), .A2(n923), .B1(n454), .B2(n920), .ZN(n2314) );
  OAI22_X1 U1567 ( .A1(n421), .A2(n923), .B1(n453), .B2(n920), .ZN(n2297) );
  OAI22_X1 U1568 ( .A1(n420), .A2(n923), .B1(n452), .B2(n920), .ZN(n2280) );
  OAI22_X1 U1569 ( .A1(n419), .A2(n923), .B1(n451), .B2(n920), .ZN(n2263) );
  OAI22_X1 U1570 ( .A1(n418), .A2(n923), .B1(n450), .B2(n920), .ZN(n2246) );
  OAI22_X1 U1571 ( .A1(n417), .A2(n923), .B1(n449), .B2(n920), .ZN(n2223) );
  OAI22_X1 U1572 ( .A1(n448), .A2(n1280), .B1(n480), .B2(n1254), .ZN(n2178) );
  OAI22_X1 U1573 ( .A1(n320), .A2(n1066), .B1(n352), .B2(n1063), .ZN(n2181) );
  OAI22_X1 U1574 ( .A1(n447), .A2(n1280), .B1(n479), .B2(n1254), .ZN(n2148) );
  OAI22_X1 U1575 ( .A1(n319), .A2(n1066), .B1(n351), .B2(n1063), .ZN(n2149) );
  OAI22_X1 U1576 ( .A1(n446), .A2(n1280), .B1(n478), .B2(n1254), .ZN(n2131) );
  OAI22_X1 U1577 ( .A1(n318), .A2(n1066), .B1(n350), .B2(n1063), .ZN(n2132) );
  OAI22_X1 U1578 ( .A1(n445), .A2(n1280), .B1(n477), .B2(n1254), .ZN(n2114) );
  OAI22_X1 U1579 ( .A1(n317), .A2(n1066), .B1(n349), .B2(n1063), .ZN(n2115) );
  OAI22_X1 U1580 ( .A1(n444), .A2(n1280), .B1(n476), .B2(n1254), .ZN(n2097) );
  OAI22_X1 U1581 ( .A1(n316), .A2(n1066), .B1(n348), .B2(n1063), .ZN(n2098) );
  OAI22_X1 U1582 ( .A1(n443), .A2(n1280), .B1(n475), .B2(n1254), .ZN(n2080) );
  OAI22_X1 U1583 ( .A1(n315), .A2(n1066), .B1(n347), .B2(n1063), .ZN(n2081) );
  OAI22_X1 U1584 ( .A1(n442), .A2(n1280), .B1(n474), .B2(n1254), .ZN(n2063) );
  OAI22_X1 U1585 ( .A1(n314), .A2(n1066), .B1(n346), .B2(n1063), .ZN(n2064) );
  OAI22_X1 U1586 ( .A1(n441), .A2(n1280), .B1(n473), .B2(n1254), .ZN(n2046) );
  OAI22_X1 U1587 ( .A1(n313), .A2(n1066), .B1(n345), .B2(n1063), .ZN(n2047) );
  OAI22_X1 U1588 ( .A1(n440), .A2(n1280), .B1(n472), .B2(n1254), .ZN(n2029) );
  OAI22_X1 U1589 ( .A1(n312), .A2(n1066), .B1(n344), .B2(n1063), .ZN(n2030) );
  OAI22_X1 U1590 ( .A1(n439), .A2(n1280), .B1(n471), .B2(n1254), .ZN(n2012) );
  OAI22_X1 U1591 ( .A1(n311), .A2(n1066), .B1(n343), .B2(n1063), .ZN(n2013) );
  OAI22_X1 U1592 ( .A1(n438), .A2(n1280), .B1(n470), .B2(n1254), .ZN(n1995) );
  OAI22_X1 U1593 ( .A1(n310), .A2(n1066), .B1(n342), .B2(n1063), .ZN(n1996) );
  OAI22_X1 U1594 ( .A1(n437), .A2(n1280), .B1(n469), .B2(n1254), .ZN(n1978) );
  OAI22_X1 U1595 ( .A1(n309), .A2(n1066), .B1(n341), .B2(n1063), .ZN(n1979) );
  OAI22_X1 U1596 ( .A1(n436), .A2(n1281), .B1(n468), .B2(n1258), .ZN(n1961) );
  OAI22_X1 U1597 ( .A1(n308), .A2(n1067), .B1(n340), .B2(n1064), .ZN(n1962) );
  OAI22_X1 U1598 ( .A1(n435), .A2(n1281), .B1(n467), .B2(n1258), .ZN(n1944) );
  OAI22_X1 U1599 ( .A1(n307), .A2(n1067), .B1(n339), .B2(n1064), .ZN(n1945) );
  OAI22_X1 U1600 ( .A1(n434), .A2(n1281), .B1(n466), .B2(n1258), .ZN(n1927) );
  OAI22_X1 U1601 ( .A1(n306), .A2(n1067), .B1(n338), .B2(n1064), .ZN(n1928) );
  OAI22_X1 U1602 ( .A1(n433), .A2(n1281), .B1(n465), .B2(n1258), .ZN(n1910) );
  OAI22_X1 U1603 ( .A1(n305), .A2(n1067), .B1(n337), .B2(n1064), .ZN(n1911) );
  OAI22_X1 U1604 ( .A1(n432), .A2(n1281), .B1(n464), .B2(n1258), .ZN(n1893) );
  OAI22_X1 U1605 ( .A1(n304), .A2(n1067), .B1(n336), .B2(n1064), .ZN(n1894) );
  OAI22_X1 U1606 ( .A1(n431), .A2(n1281), .B1(n463), .B2(n1258), .ZN(n1876) );
  OAI22_X1 U1607 ( .A1(n303), .A2(n1067), .B1(n335), .B2(n1064), .ZN(n1877) );
  OAI22_X1 U1608 ( .A1(n430), .A2(n1281), .B1(n462), .B2(n1258), .ZN(n1859) );
  OAI22_X1 U1609 ( .A1(n302), .A2(n1067), .B1(n334), .B2(n1064), .ZN(n1860) );
  OAI22_X1 U1610 ( .A1(n429), .A2(n1281), .B1(n461), .B2(n1258), .ZN(n1842) );
  OAI22_X1 U1611 ( .A1(n301), .A2(n1067), .B1(n333), .B2(n1064), .ZN(n1843) );
  OAI22_X1 U1612 ( .A1(n428), .A2(n1281), .B1(n460), .B2(n1258), .ZN(n1825) );
  OAI22_X1 U1613 ( .A1(n300), .A2(n1067), .B1(n332), .B2(n1064), .ZN(n1826) );
  OAI22_X1 U1614 ( .A1(n427), .A2(n1281), .B1(n459), .B2(n1258), .ZN(n1808) );
  OAI22_X1 U1615 ( .A1(n299), .A2(n1067), .B1(n331), .B2(n1064), .ZN(n1809) );
  OAI22_X1 U1616 ( .A1(n426), .A2(n1281), .B1(n458), .B2(n1258), .ZN(n1791) );
  OAI22_X1 U1617 ( .A1(n298), .A2(n1067), .B1(n330), .B2(n1064), .ZN(n1792) );
  OAI22_X1 U1618 ( .A1(n425), .A2(n1281), .B1(n457), .B2(n1258), .ZN(n1774) );
  OAI22_X1 U1619 ( .A1(n297), .A2(n1067), .B1(n329), .B2(n1064), .ZN(n1775) );
  OAI22_X1 U1620 ( .A1(n448), .A2(n921), .B1(n480), .B2(n918), .ZN(n2769) );
  OAI22_X1 U1621 ( .A1(n320), .A2(n909), .B1(n352), .B2(n906), .ZN(n2772) );
  OAI22_X1 U1622 ( .A1(n447), .A2(n921), .B1(n479), .B2(n918), .ZN(n2739) );
  OAI22_X1 U1623 ( .A1(n319), .A2(n909), .B1(n351), .B2(n906), .ZN(n2740) );
  OAI22_X1 U1624 ( .A1(n446), .A2(n921), .B1(n478), .B2(n918), .ZN(n2722) );
  OAI22_X1 U1625 ( .A1(n318), .A2(n909), .B1(n350), .B2(n906), .ZN(n2723) );
  OAI22_X1 U1626 ( .A1(n445), .A2(n921), .B1(n477), .B2(n918), .ZN(n2705) );
  OAI22_X1 U1627 ( .A1(n317), .A2(n909), .B1(n349), .B2(n906), .ZN(n2706) );
  OAI22_X1 U1628 ( .A1(n444), .A2(n921), .B1(n476), .B2(n918), .ZN(n2688) );
  OAI22_X1 U1629 ( .A1(n316), .A2(n909), .B1(n348), .B2(n906), .ZN(n2689) );
  OAI22_X1 U1630 ( .A1(n443), .A2(n921), .B1(n475), .B2(n918), .ZN(n2671) );
  OAI22_X1 U1631 ( .A1(n315), .A2(n909), .B1(n347), .B2(n906), .ZN(n2672) );
  OAI22_X1 U1632 ( .A1(n442), .A2(n921), .B1(n474), .B2(n918), .ZN(n2654) );
  OAI22_X1 U1633 ( .A1(n314), .A2(n909), .B1(n346), .B2(n906), .ZN(n2655) );
  OAI22_X1 U1634 ( .A1(n441), .A2(n921), .B1(n473), .B2(n918), .ZN(n2637) );
  OAI22_X1 U1635 ( .A1(n313), .A2(n909), .B1(n345), .B2(n906), .ZN(n2638) );
  OAI22_X1 U1636 ( .A1(n440), .A2(n921), .B1(n472), .B2(n918), .ZN(n2620) );
  OAI22_X1 U1637 ( .A1(n312), .A2(n909), .B1(n344), .B2(n906), .ZN(n2621) );
  OAI22_X1 U1638 ( .A1(n439), .A2(n921), .B1(n471), .B2(n918), .ZN(n2603) );
  OAI22_X1 U1639 ( .A1(n311), .A2(n909), .B1(n343), .B2(n906), .ZN(n2604) );
  OAI22_X1 U1640 ( .A1(n438), .A2(n921), .B1(n470), .B2(n918), .ZN(n2586) );
  OAI22_X1 U1641 ( .A1(n310), .A2(n909), .B1(n342), .B2(n906), .ZN(n2587) );
  OAI22_X1 U1642 ( .A1(n437), .A2(n921), .B1(n469), .B2(n918), .ZN(n2569) );
  OAI22_X1 U1643 ( .A1(n309), .A2(n909), .B1(n341), .B2(n906), .ZN(n2570) );
  OAI22_X1 U1644 ( .A1(n436), .A2(n922), .B1(n468), .B2(n919), .ZN(n2552) );
  OAI22_X1 U1645 ( .A1(n308), .A2(n910), .B1(n340), .B2(n907), .ZN(n2553) );
  OAI22_X1 U1646 ( .A1(n435), .A2(n922), .B1(n467), .B2(n919), .ZN(n2535) );
  OAI22_X1 U1647 ( .A1(n307), .A2(n910), .B1(n339), .B2(n907), .ZN(n2536) );
  OAI22_X1 U1648 ( .A1(n434), .A2(n922), .B1(n466), .B2(n919), .ZN(n2518) );
  OAI22_X1 U1649 ( .A1(n306), .A2(n910), .B1(n338), .B2(n907), .ZN(n2519) );
  OAI22_X1 U1650 ( .A1(n433), .A2(n922), .B1(n465), .B2(n919), .ZN(n2501) );
  OAI22_X1 U1651 ( .A1(n305), .A2(n910), .B1(n337), .B2(n907), .ZN(n2502) );
  OAI22_X1 U1652 ( .A1(n432), .A2(n922), .B1(n464), .B2(n919), .ZN(n2484) );
  OAI22_X1 U1653 ( .A1(n304), .A2(n910), .B1(n336), .B2(n907), .ZN(n2485) );
  OAI22_X1 U1654 ( .A1(n431), .A2(n922), .B1(n463), .B2(n919), .ZN(n2467) );
  OAI22_X1 U1655 ( .A1(n303), .A2(n910), .B1(n335), .B2(n907), .ZN(n2468) );
  OAI22_X1 U1656 ( .A1(n430), .A2(n922), .B1(n462), .B2(n919), .ZN(n2450) );
  OAI22_X1 U1657 ( .A1(n302), .A2(n910), .B1(n334), .B2(n907), .ZN(n2451) );
  OAI22_X1 U1658 ( .A1(n429), .A2(n922), .B1(n461), .B2(n919), .ZN(n2433) );
  OAI22_X1 U1659 ( .A1(n301), .A2(n910), .B1(n333), .B2(n907), .ZN(n2434) );
  OAI22_X1 U1660 ( .A1(n428), .A2(n922), .B1(n460), .B2(n919), .ZN(n2416) );
  OAI22_X1 U1661 ( .A1(n300), .A2(n910), .B1(n332), .B2(n907), .ZN(n2417) );
  OAI22_X1 U1662 ( .A1(n427), .A2(n922), .B1(n459), .B2(n919), .ZN(n2399) );
  OAI22_X1 U1663 ( .A1(n299), .A2(n910), .B1(n331), .B2(n907), .ZN(n2400) );
  OAI22_X1 U1664 ( .A1(n426), .A2(n922), .B1(n458), .B2(n919), .ZN(n2382) );
  OAI22_X1 U1665 ( .A1(n298), .A2(n910), .B1(n330), .B2(n907), .ZN(n2383) );
  OAI22_X1 U1666 ( .A1(n425), .A2(n922), .B1(n457), .B2(n919), .ZN(n2365) );
  OAI22_X1 U1667 ( .A1(n297), .A2(n910), .B1(n329), .B2(n907), .ZN(n2366) );
  OAI22_X1 U1668 ( .A1(n40), .A2(n1558), .B1(n72), .B2(n1555), .ZN(n1755) );
  OAI22_X1 U1669 ( .A1(n39), .A2(n1558), .B1(n71), .B2(n1555), .ZN(n1738) );
  OAI22_X1 U1670 ( .A1(n38), .A2(n1558), .B1(n70), .B2(n1555), .ZN(n1721) );
  OAI22_X1 U1671 ( .A1(n37), .A2(n1558), .B1(n69), .B2(n1555), .ZN(n1704) );
  OAI22_X1 U1672 ( .A1(n36), .A2(n1558), .B1(n68), .B2(n1555), .ZN(n1687) );
  OAI22_X1 U1673 ( .A1(n35), .A2(n1558), .B1(n67), .B2(n1555), .ZN(n1670) );
  OAI22_X1 U1674 ( .A1(n34), .A2(n1558), .B1(n66), .B2(n1555), .ZN(n1653) );
  OAI22_X1 U1675 ( .A1(n33), .A2(n1558), .B1(n65), .B2(n1555), .ZN(n1622) );
  OAI22_X1 U1676 ( .A1(n40), .A2(n1011), .B1(n72), .B2(n1008), .ZN(n2346) );
  OAI22_X1 U1677 ( .A1(n39), .A2(n1011), .B1(n71), .B2(n1008), .ZN(n2329) );
  OAI22_X1 U1678 ( .A1(n38), .A2(n1011), .B1(n70), .B2(n1008), .ZN(n2312) );
  OAI22_X1 U1679 ( .A1(n37), .A2(n1011), .B1(n69), .B2(n1008), .ZN(n2295) );
  OAI22_X1 U1680 ( .A1(n36), .A2(n1011), .B1(n68), .B2(n1008), .ZN(n2278) );
  OAI22_X1 U1681 ( .A1(n35), .A2(n1011), .B1(n67), .B2(n1008), .ZN(n2261) );
  OAI22_X1 U1682 ( .A1(n34), .A2(n1011), .B1(n66), .B2(n1008), .ZN(n2244) );
  OAI22_X1 U1683 ( .A1(n33), .A2(n1011), .B1(n65), .B2(n1008), .ZN(n2213) );
  OAI22_X1 U1684 ( .A1(n64), .A2(n1556), .B1(n96), .B2(n1432), .ZN(n2173) );
  OAI22_X1 U1685 ( .A1(n63), .A2(n1556), .B1(n95), .B2(n1432), .ZN(n2146) );
  OAI22_X1 U1686 ( .A1(n62), .A2(n1556), .B1(n94), .B2(n1432), .ZN(n2129) );
  OAI22_X1 U1687 ( .A1(n61), .A2(n1556), .B1(n93), .B2(n1432), .ZN(n2112) );
  OAI22_X1 U1688 ( .A1(n60), .A2(n1556), .B1(n92), .B2(n1432), .ZN(n2095) );
  OAI22_X1 U1689 ( .A1(n59), .A2(n1556), .B1(n91), .B2(n1432), .ZN(n2078) );
  OAI22_X1 U1690 ( .A1(n58), .A2(n1556), .B1(n90), .B2(n1432), .ZN(n2061) );
  OAI22_X1 U1691 ( .A1(n57), .A2(n1556), .B1(n89), .B2(n1432), .ZN(n2044) );
  OAI22_X1 U1692 ( .A1(n56), .A2(n1556), .B1(n88), .B2(n1432), .ZN(n2027) );
  OAI22_X1 U1693 ( .A1(n55), .A2(n1556), .B1(n87), .B2(n1432), .ZN(n2010) );
  OAI22_X1 U1694 ( .A1(n54), .A2(n1556), .B1(n86), .B2(n1432), .ZN(n1993) );
  OAI22_X1 U1695 ( .A1(n53), .A2(n1556), .B1(n85), .B2(n1432), .ZN(n1976) );
  OAI22_X1 U1696 ( .A1(n52), .A2(n1557), .B1(n84), .B2(n1445), .ZN(n1959) );
  OAI22_X1 U1697 ( .A1(n51), .A2(n1557), .B1(n83), .B2(n1445), .ZN(n1942) );
  OAI22_X1 U1698 ( .A1(n50), .A2(n1557), .B1(n82), .B2(n1445), .ZN(n1925) );
  OAI22_X1 U1699 ( .A1(n49), .A2(n1557), .B1(n81), .B2(n1445), .ZN(n1908) );
  OAI22_X1 U1700 ( .A1(n48), .A2(n1557), .B1(n80), .B2(n1445), .ZN(n1891) );
  OAI22_X1 U1701 ( .A1(n47), .A2(n1557), .B1(n79), .B2(n1445), .ZN(n1874) );
  OAI22_X1 U1702 ( .A1(n46), .A2(n1557), .B1(n78), .B2(n1445), .ZN(n1857) );
  OAI22_X1 U1703 ( .A1(n45), .A2(n1557), .B1(n77), .B2(n1445), .ZN(n1840) );
  OAI22_X1 U1704 ( .A1(n44), .A2(n1557), .B1(n76), .B2(n1445), .ZN(n1823) );
  OAI22_X1 U1705 ( .A1(n43), .A2(n1557), .B1(n75), .B2(n1445), .ZN(n1806) );
  OAI22_X1 U1706 ( .A1(n42), .A2(n1557), .B1(n74), .B2(n1445), .ZN(n1789) );
  OAI22_X1 U1707 ( .A1(n41), .A2(n1557), .B1(n73), .B2(n1445), .ZN(n1772) );
  OAI22_X1 U1708 ( .A1(n64), .A2(n1009), .B1(n96), .B2(n1006), .ZN(n2764) );
  OAI22_X1 U1709 ( .A1(n63), .A2(n1009), .B1(n95), .B2(n1006), .ZN(n2737) );
  OAI22_X1 U1710 ( .A1(n62), .A2(n1009), .B1(n94), .B2(n1006), .ZN(n2720) );
  OAI22_X1 U1711 ( .A1(n61), .A2(n1009), .B1(n93), .B2(n1006), .ZN(n2703) );
  OAI22_X1 U1712 ( .A1(n60), .A2(n1009), .B1(n92), .B2(n1006), .ZN(n2686) );
  OAI22_X1 U1713 ( .A1(n59), .A2(n1009), .B1(n91), .B2(n1006), .ZN(n2669) );
  OAI22_X1 U1714 ( .A1(n58), .A2(n1009), .B1(n90), .B2(n1006), .ZN(n2652) );
  OAI22_X1 U1715 ( .A1(n57), .A2(n1009), .B1(n89), .B2(n1006), .ZN(n2635) );
  OAI22_X1 U1716 ( .A1(n56), .A2(n1009), .B1(n88), .B2(n1006), .ZN(n2618) );
  OAI22_X1 U1717 ( .A1(n55), .A2(n1009), .B1(n87), .B2(n1006), .ZN(n2601) );
  OAI22_X1 U1718 ( .A1(n54), .A2(n1009), .B1(n86), .B2(n1006), .ZN(n2584) );
  OAI22_X1 U1719 ( .A1(n53), .A2(n1009), .B1(n85), .B2(n1006), .ZN(n2567) );
  OAI22_X1 U1720 ( .A1(n52), .A2(n1010), .B1(n84), .B2(n1007), .ZN(n2550) );
  OAI22_X1 U1721 ( .A1(n51), .A2(n1010), .B1(n83), .B2(n1007), .ZN(n2533) );
  OAI22_X1 U1722 ( .A1(n50), .A2(n1010), .B1(n82), .B2(n1007), .ZN(n2516) );
  OAI22_X1 U1723 ( .A1(n49), .A2(n1010), .B1(n81), .B2(n1007), .ZN(n2499) );
  OAI22_X1 U1724 ( .A1(n48), .A2(n1010), .B1(n80), .B2(n1007), .ZN(n2482) );
  OAI22_X1 U1725 ( .A1(n47), .A2(n1010), .B1(n79), .B2(n1007), .ZN(n2465) );
  OAI22_X1 U1726 ( .A1(n46), .A2(n1010), .B1(n78), .B2(n1007), .ZN(n2448) );
  OAI22_X1 U1727 ( .A1(n45), .A2(n1010), .B1(n77), .B2(n1007), .ZN(n2431) );
  OAI22_X1 U1728 ( .A1(n44), .A2(n1010), .B1(n76), .B2(n1007), .ZN(n2414) );
  OAI22_X1 U1729 ( .A1(n43), .A2(n1010), .B1(n75), .B2(n1007), .ZN(n2397) );
  OAI22_X1 U1730 ( .A1(n42), .A2(n1010), .B1(n74), .B2(n1007), .ZN(n2380) );
  OAI22_X1 U1731 ( .A1(n41), .A2(n1010), .B1(n73), .B2(n1007), .ZN(n2363) );
  OAI22_X1 U1732 ( .A1(n253), .A2(n674), .B1(n29), .B2(n952), .ZN(n2814) );
  OAI22_X1 U1733 ( .A1(n370), .A2(n673), .B1(n241), .B2(n951), .ZN(n2815) );
  OAI22_X1 U1734 ( .A1(n4201), .A2(n3573), .B1(n29), .B2(n950), .ZN(n2816) );
  OAI22_X1 U1735 ( .A1(n4200), .A2(n674), .B1(n29), .B2(n949), .ZN(n2817) );
  OAI22_X1 U1736 ( .A1(n786), .A2(n3573), .B1(n240), .B2(n948), .ZN(n2818) );
  OAI22_X1 U1737 ( .A1(n784), .A2(n3575), .B1(n29), .B2(n947), .ZN(n2819) );
  OAI22_X1 U1738 ( .A1(n781), .A2(n3575), .B1(n29), .B2(n946), .ZN(n2820) );
  OAI22_X1 U1739 ( .A1(n778), .A2(n3573), .B1(n29), .B2(n945), .ZN(n2821) );
  OAI22_X1 U1740 ( .A1(n775), .A2(n3574), .B1(n29), .B2(n944), .ZN(n2822) );
  OAI22_X1 U1741 ( .A1(n772), .A2(n560), .B1(n29), .B2(n943), .ZN(n2823) );
  OAI22_X1 U1742 ( .A1(n769), .A2(n3574), .B1(n29), .B2(n942), .ZN(n2824) );
  OAI22_X1 U1743 ( .A1(n677), .A2(n673), .B1(n29), .B2(n941), .ZN(n2825) );
  OAI22_X1 U1744 ( .A1(n4191), .A2(n3575), .B1(n239), .B2(n940), .ZN(n2826) );
  OAI22_X1 U1745 ( .A1(n4190), .A2(n3575), .B1(n239), .B2(n939), .ZN(n2827) );
  OAI22_X1 U1746 ( .A1(n4189), .A2(n3574), .B1(n29), .B2(n938), .ZN(n2828) );
  OAI22_X1 U1747 ( .A1(n287), .A2(n560), .B1(n239), .B2(n937), .ZN(n2829) );
  OAI22_X1 U1748 ( .A1(n4187), .A2(n673), .B1(n239), .B2(n936), .ZN(n2830) );
  OAI22_X1 U1749 ( .A1(n283), .A2(n674), .B1(n240), .B2(n935), .ZN(n2831) );
  OAI22_X1 U1750 ( .A1(n4185), .A2(n238), .B1(n241), .B2(n934), .ZN(n2832) );
  OAI22_X1 U1751 ( .A1(n4184), .A2(n674), .B1(n240), .B2(n933), .ZN(n2833) );
  OAI22_X1 U1752 ( .A1(n683), .A2(n3573), .B1(n241), .B2(n932), .ZN(n2834) );
  OAI22_X1 U1753 ( .A1(n376), .A2(n673), .B1(n240), .B2(n931), .ZN(n2835) );
  OAI22_X1 U1754 ( .A1(n4181), .A2(n410), .B1(n3578), .B2(n930), .ZN(n2836) );
  OAI22_X1 U1755 ( .A1(n4180), .A2(n673), .B1(n3578), .B2(n929), .ZN(n2837) );
  OAI22_X1 U1756 ( .A1(n254), .A2(n3549), .B1(n3552), .B2(n856), .ZN(n2846) );
  OAI22_X1 U1757 ( .A1(n370), .A2(n3549), .B1(n3552), .B2(n855), .ZN(n2847) );
  OAI22_X1 U1758 ( .A1(n4201), .A2(n3549), .B1(n3553), .B2(n854), .ZN(n2848)
         );
  OAI22_X1 U1759 ( .A1(n789), .A2(n3549), .B1(n3553), .B2(n853), .ZN(n2849) );
  OAI22_X1 U1760 ( .A1(n4199), .A2(n3549), .B1(n3553), .B2(n852), .ZN(n2850)
         );
  OAI22_X1 U1761 ( .A1(n4198), .A2(n3549), .B1(n3553), .B2(n851), .ZN(n2851)
         );
  OAI22_X1 U1762 ( .A1(n4197), .A2(n3549), .B1(n3553), .B2(n850), .ZN(n2852)
         );
  OAI22_X1 U1763 ( .A1(n4196), .A2(n3548), .B1(n3554), .B2(n849), .ZN(n2853)
         );
  OAI22_X1 U1764 ( .A1(n4195), .A2(n728), .B1(n3554), .B2(n848), .ZN(n2854) );
  OAI22_X1 U1765 ( .A1(n4194), .A2(n727), .B1(n3554), .B2(n847), .ZN(n2855) );
  OAI22_X1 U1766 ( .A1(n4193), .A2(n3550), .B1(n3554), .B2(n846), .ZN(n2856)
         );
  OAI22_X1 U1767 ( .A1(n4192), .A2(n3548), .B1(n3554), .B2(n845), .ZN(n2857)
         );
  OAI22_X1 U1768 ( .A1(n687), .A2(n728), .B1(n3555), .B2(n844), .ZN(n2858) );
  OAI22_X1 U1769 ( .A1(n4190), .A2(n727), .B1(n3555), .B2(n843), .ZN(n2859) );
  OAI22_X1 U1770 ( .A1(n4189), .A2(n3550), .B1(n3555), .B2(n842), .ZN(n2860)
         );
  OAI22_X1 U1771 ( .A1(n286), .A2(n3548), .B1(n3555), .B2(n841), .ZN(n2861) );
  OAI22_X1 U1772 ( .A1(n4187), .A2(n728), .B1(n3555), .B2(n840), .ZN(n2862) );
  OAI22_X1 U1773 ( .A1(n284), .A2(n727), .B1(n3556), .B2(n839), .ZN(n2863) );
  OAI22_X1 U1774 ( .A1(n684), .A2(n3550), .B1(n3556), .B2(n838), .ZN(n2864) );
  OAI22_X1 U1775 ( .A1(n271), .A2(n3548), .B1(n3556), .B2(n837), .ZN(n2865) );
  OAI22_X1 U1776 ( .A1(n4183), .A2(n728), .B1(n3556), .B2(n836), .ZN(n2866) );
  OAI22_X1 U1777 ( .A1(n377), .A2(n727), .B1(n3556), .B2(n835), .ZN(n2867) );
  OAI22_X1 U1778 ( .A1(n247), .A2(n3550), .B1(n3557), .B2(n834), .ZN(n2868) );
  OAI22_X1 U1779 ( .A1(n4180), .A2(n3548), .B1(n3556), .B2(n833), .ZN(n2869)
         );
  OAI22_X1 U1780 ( .A1(n4203), .A2(n732), .B1(n3546), .B2(n824), .ZN(n2878) );
  OAI22_X1 U1781 ( .A1(n369), .A2(n731), .B1(n3543), .B2(n823), .ZN(n2879) );
  OAI22_X1 U1782 ( .A1(n4201), .A2(n732), .B1(n3545), .B2(n822), .ZN(n2880) );
  OAI22_X1 U1783 ( .A1(n168), .A2(n3539), .B1(n3542), .B2(n821), .ZN(n2881) );
  OAI22_X1 U1784 ( .A1(n4199), .A2(n3538), .B1(n3546), .B2(n820), .ZN(n2882)
         );
  OAI22_X1 U1785 ( .A1(n4198), .A2(n3539), .B1(n3545), .B2(n819), .ZN(n2883)
         );
  OAI22_X1 U1786 ( .A1(n4197), .A2(n732), .B1(n3544), .B2(n818), .ZN(n2884) );
  OAI22_X1 U1787 ( .A1(n4196), .A2(n572), .B1(n3546), .B2(n817), .ZN(n2885) );
  OAI22_X1 U1788 ( .A1(n4195), .A2(n3540), .B1(n3545), .B2(n816), .ZN(n2886)
         );
  OAI22_X1 U1789 ( .A1(n4194), .A2(n732), .B1(n3541), .B2(n815), .ZN(n2887) );
  OAI22_X1 U1790 ( .A1(n4193), .A2(n731), .B1(n3541), .B2(n814), .ZN(n2888) );
  OAI22_X1 U1791 ( .A1(n192), .A2(n731), .B1(n3542), .B2(n813), .ZN(n2889) );
  OAI22_X1 U1792 ( .A1(n172), .A2(n732), .B1(n3543), .B2(n812), .ZN(n2890) );
  OAI22_X1 U1793 ( .A1(n257), .A2(n3538), .B1(n3546), .B2(n811), .ZN(n2891) );
  OAI22_X1 U1794 ( .A1(n4189), .A2(n3538), .B1(n3541), .B2(n810), .ZN(n2892)
         );
  OAI22_X1 U1795 ( .A1(n287), .A2(n3540), .B1(n3541), .B2(n809), .ZN(n2893) );
  OAI22_X1 U1796 ( .A1(n686), .A2(n3538), .B1(n3542), .B2(n808), .ZN(n2894) );
  OAI22_X1 U1797 ( .A1(n283), .A2(n3539), .B1(n3543), .B2(n807), .ZN(n2895) );
  OAI22_X1 U1798 ( .A1(n171), .A2(n732), .B1(n3544), .B2(n806), .ZN(n2896) );
  OAI22_X1 U1799 ( .A1(n716), .A2(n572), .B1(n3543), .B2(n805), .ZN(n2897) );
  OAI22_X1 U1800 ( .A1(n683), .A2(n572), .B1(n3541), .B2(n804), .ZN(n2898) );
  OAI22_X1 U1801 ( .A1(n378), .A2(n3540), .B1(n3542), .B2(n803), .ZN(n2899) );
  OAI22_X1 U1802 ( .A1(n680), .A2(n3539), .B1(n3547), .B2(n802), .ZN(n2900) );
  OAI22_X1 U1803 ( .A1(n5), .A2(n572), .B1(n178), .B2(n801), .ZN(n2901) );
  OAI22_X1 U1804 ( .A1(n254), .A2(n577), .B1(n3506), .B2(n664), .ZN(n2910) );
  OAI22_X1 U1805 ( .A1(n369), .A2(n3502), .B1(n3510), .B2(n663), .ZN(n2911) );
  OAI22_X1 U1806 ( .A1(n3503), .A2(n4201), .B1(n3510), .B2(n662), .ZN(n2912)
         );
  OAI22_X1 U1807 ( .A1(n789), .A2(n3504), .B1(n3510), .B2(n661), .ZN(n2913) );
  OAI22_X1 U1808 ( .A1(n4199), .A2(n738), .B1(n3505), .B2(n660), .ZN(n2914) );
  OAI22_X1 U1809 ( .A1(n4198), .A2(n3504), .B1(n3505), .B2(n659), .ZN(n2915)
         );
  OAI22_X1 U1810 ( .A1(n4197), .A2(n577), .B1(n3505), .B2(n658), .ZN(n2916) );
  OAI22_X1 U1811 ( .A1(n4196), .A2(n738), .B1(n3509), .B2(n657), .ZN(n2917) );
  OAI22_X1 U1812 ( .A1(n4195), .A2(n3503), .B1(n3507), .B2(n656), .ZN(n2918)
         );
  OAI22_X1 U1813 ( .A1(n4194), .A2(n738), .B1(n3506), .B2(n655), .ZN(n2919) );
  OAI22_X1 U1814 ( .A1(n3502), .A2(n4193), .B1(n3509), .B2(n654), .ZN(n2920)
         );
  OAI22_X1 U1815 ( .A1(n3502), .A2(n192), .B1(n3509), .B2(n653), .ZN(n2921) );
  OAI22_X1 U1816 ( .A1(n3503), .A2(n688), .B1(n3508), .B2(n652), .ZN(n2922) );
  OAI22_X1 U1817 ( .A1(n10), .A2(n3502), .B1(n3509), .B2(n651), .ZN(n2923) );
  OAI22_X1 U1818 ( .A1(n4189), .A2(n577), .B1(n3506), .B2(n650), .ZN(n2924) );
  OAI22_X1 U1819 ( .A1(n287), .A2(n3504), .B1(n3507), .B2(n649), .ZN(n2925) );
  OAI22_X1 U1820 ( .A1(n167), .A2(n3504), .B1(n3510), .B2(n648), .ZN(n2926) );
  OAI22_X1 U1821 ( .A1(n3503), .A2(n284), .B1(n3505), .B2(n647), .ZN(n2927) );
  OAI22_X1 U1822 ( .A1(n685), .A2(n3503), .B1(n3508), .B2(n646), .ZN(n2928) );
  OAI22_X1 U1823 ( .A1(n4184), .A2(n577), .B1(n3508), .B2(n645), .ZN(n2929) );
  OAI22_X1 U1824 ( .A1(n3502), .A2(n4183), .B1(n3507), .B2(n644), .ZN(n2930)
         );
  OAI22_X1 U1825 ( .A1(n377), .A2(n577), .B1(n3508), .B2(n643), .ZN(n2931) );
  OAI22_X1 U1826 ( .A1(n738), .A2(n681), .B1(n281), .B2(n642), .ZN(n2932) );
  OAI22_X1 U1827 ( .A1(n713), .A2(n3504), .B1(n281), .B2(n641), .ZN(n2933) );
  OAI22_X1 U1828 ( .A1(n254), .A2(n579), .B1(n3497), .B2(n632), .ZN(n2942) );
  OAI22_X1 U1829 ( .A1(n370), .A2(n579), .B1(n3498), .B2(n631), .ZN(n2943) );
  OAI22_X1 U1830 ( .A1(n579), .A2(n758), .B1(n3496), .B2(n630), .ZN(n2944) );
  OAI22_X1 U1831 ( .A1(n4200), .A2(n3494), .B1(n3500), .B2(n629), .ZN(n2945)
         );
  OAI22_X1 U1832 ( .A1(n4199), .A2(n3492), .B1(n3499), .B2(n628), .ZN(n2946)
         );
  OAI22_X1 U1833 ( .A1(n4198), .A2(n3494), .B1(n3496), .B2(n627), .ZN(n2947)
         );
  OAI22_X1 U1834 ( .A1(n4197), .A2(n3493), .B1(n3497), .B2(n626), .ZN(n2948)
         );
  OAI22_X1 U1835 ( .A1(n4196), .A2(n3493), .B1(n3497), .B2(n625), .ZN(n2949)
         );
  OAI22_X1 U1836 ( .A1(n4195), .A2(n579), .B1(n3498), .B2(n624), .ZN(n2950) );
  OAI22_X1 U1837 ( .A1(n4194), .A2(n735), .B1(n3500), .B2(n623), .ZN(n2951) );
  OAI22_X1 U1838 ( .A1(n4193), .A2(n735), .B1(n3499), .B2(n622), .ZN(n2952) );
  OAI22_X1 U1839 ( .A1(n4192), .A2(n3494), .B1(n3498), .B2(n621), .ZN(n2953)
         );
  OAI22_X1 U1840 ( .A1(n4191), .A2(n3492), .B1(n3495), .B2(n620), .ZN(n2954)
         );
  OAI22_X1 U1841 ( .A1(n257), .A2(n579), .B1(n619), .B2(n3495), .ZN(n2955) );
  OAI22_X1 U1842 ( .A1(n607), .A2(n3492), .B1(n3497), .B2(n618), .ZN(n2956) );
  OAI22_X1 U1843 ( .A1(n286), .A2(n3492), .B1(n3499), .B2(n617), .ZN(n2957) );
  OAI22_X1 U1844 ( .A1(n579), .A2(n166), .B1(n3496), .B2(n616), .ZN(n2958) );
  OAI22_X1 U1845 ( .A1(n3493), .A2(n284), .B1(n3495), .B2(n615), .ZN(n2959) );
  OAI22_X1 U1846 ( .A1(n4185), .A2(n579), .B1(n614), .B2(n3495), .ZN(n2960) );
  OAI22_X1 U1847 ( .A1(n716), .A2(n735), .B1(n3495), .B2(n613), .ZN(n2961) );
  OAI22_X1 U1848 ( .A1(n682), .A2(n3494), .B1(n3498), .B2(n612), .ZN(n2962) );
  OAI22_X1 U1849 ( .A1(n378), .A2(n3492), .B1(n3500), .B2(n611), .ZN(n2963) );
  OAI22_X1 U1850 ( .A1(n4181), .A2(n3492), .B1(n359), .B2(n610), .ZN(n2964) );
  OAI22_X1 U1851 ( .A1(n5), .A2(n3494), .B1(n359), .B2(n609), .ZN(n2965) );
  OAI22_X1 U1852 ( .A1(n4203), .A2(n594), .B1(n3453), .B2(n472), .ZN(n3038) );
  OAI22_X1 U1853 ( .A1(n370), .A2(n3450), .B1(n3453), .B2(n471), .ZN(n3039) );
  OAI22_X1 U1854 ( .A1(n758), .A2(n372), .B1(n3454), .B2(n470), .ZN(n3040) );
  OAI22_X1 U1855 ( .A1(n168), .A2(n372), .B1(n3454), .B2(n469), .ZN(n3041) );
  OAI22_X1 U1856 ( .A1(n786), .A2(n3451), .B1(n3454), .B2(n468), .ZN(n3042) );
  OAI22_X1 U1857 ( .A1(n784), .A2(n593), .B1(n3454), .B2(n467), .ZN(n3043) );
  OAI22_X1 U1858 ( .A1(n781), .A2(n594), .B1(n3454), .B2(n466), .ZN(n3044) );
  OAI22_X1 U1859 ( .A1(n778), .A2(n3450), .B1(n3455), .B2(n465), .ZN(n3045) );
  OAI22_X1 U1860 ( .A1(n775), .A2(n594), .B1(n3455), .B2(n464), .ZN(n3046) );
  OAI22_X1 U1861 ( .A1(n772), .A2(n594), .B1(n3455), .B2(n463), .ZN(n3047) );
  OAI22_X1 U1862 ( .A1(n769), .A2(n3451), .B1(n3455), .B2(n462), .ZN(n3048) );
  OAI22_X1 U1863 ( .A1(n4192), .A2(n594), .B1(n3455), .B2(n461), .ZN(n3049) );
  OAI22_X1 U1864 ( .A1(n4191), .A2(n593), .B1(n3456), .B2(n460), .ZN(n3050) );
  OAI22_X1 U1865 ( .A1(n257), .A2(n593), .B1(n3456), .B2(n459), .ZN(n3051) );
  OAI22_X1 U1866 ( .A1(n607), .A2(n3451), .B1(n3456), .B2(n458), .ZN(n3052) );
  OAI22_X1 U1867 ( .A1(n287), .A2(n594), .B1(n3456), .B2(n457), .ZN(n3053) );
  OAI22_X1 U1868 ( .A1(n167), .A2(n3450), .B1(n3456), .B2(n456), .ZN(n3054) );
  OAI22_X1 U1869 ( .A1(n282), .A2(n3451), .B1(n3457), .B2(n455), .ZN(n3055) );
  OAI22_X1 U1870 ( .A1(n685), .A2(n372), .B1(n3457), .B2(n454), .ZN(n3056) );
  OAI22_X1 U1871 ( .A1(n716), .A2(n593), .B1(n3457), .B2(n453), .ZN(n3057) );
  OAI22_X1 U1872 ( .A1(n4183), .A2(n3451), .B1(n3457), .B2(n452), .ZN(n3058)
         );
  OAI22_X1 U1873 ( .A1(n376), .A2(n3450), .B1(n3457), .B2(n451), .ZN(n3059) );
  OAI22_X1 U1874 ( .A1(n680), .A2(n3450), .B1(n3458), .B2(n450), .ZN(n3060) );
  OAI22_X1 U1875 ( .A1(n713), .A2(n3450), .B1(n3458), .B2(n449), .ZN(n3061) );
  OAI22_X1 U1876 ( .A1(n254), .A2(n559), .B1(n226), .B2(n440), .ZN(n3070) );
  OAI22_X1 U1877 ( .A1(n370), .A2(n3446), .B1(n225), .B2(n439), .ZN(n3071) );
  OAI22_X1 U1878 ( .A1(n759), .A2(n3447), .B1(n225), .B2(n438), .ZN(n3072) );
  OAI22_X1 U1879 ( .A1(n4200), .A2(n698), .B1(n226), .B2(n437), .ZN(n3073) );
  OAI22_X1 U1880 ( .A1(n786), .A2(n697), .B1(n226), .B2(n436), .ZN(n3074) );
  OAI22_X1 U1881 ( .A1(n784), .A2(n559), .B1(n3448), .B2(n435), .ZN(n3075) );
  OAI22_X1 U1882 ( .A1(n781), .A2(n558), .B1(n3448), .B2(n434), .ZN(n3076) );
  OAI22_X1 U1883 ( .A1(n778), .A2(n697), .B1(n3448), .B2(n433), .ZN(n3077) );
  OAI22_X1 U1884 ( .A1(n775), .A2(n698), .B1(n3448), .B2(n432), .ZN(n3078) );
  OAI22_X1 U1885 ( .A1(n772), .A2(n697), .B1(n3448), .B2(n431), .ZN(n3079) );
  OAI22_X1 U1886 ( .A1(n769), .A2(n3446), .B1(n225), .B2(n430), .ZN(n3080) );
  OAI22_X1 U1887 ( .A1(n677), .A2(n698), .B1(n226), .B2(n429), .ZN(n3081) );
  OAI22_X1 U1888 ( .A1(n687), .A2(n3447), .B1(n3448), .B2(n428), .ZN(n3082) );
  OAI22_X1 U1889 ( .A1(n744), .A2(n698), .B1(n226), .B2(n427), .ZN(n3083) );
  OAI22_X1 U1890 ( .A1(n608), .A2(n698), .B1(n225), .B2(n426), .ZN(n3084) );
  OAI22_X1 U1891 ( .A1(n285), .A2(n558), .B1(n225), .B2(n425), .ZN(n3085) );
  OAI22_X1 U1892 ( .A1(n4187), .A2(n559), .B1(n226), .B2(n424), .ZN(n3086) );
  OAI22_X1 U1893 ( .A1(n282), .A2(n3447), .B1(n226), .B2(n423), .ZN(n3087) );
  OAI22_X1 U1894 ( .A1(n171), .A2(n3447), .B1(n225), .B2(n422), .ZN(n3088) );
  OAI22_X1 U1895 ( .A1(n24), .A2(n558), .B1(n226), .B2(n421), .ZN(n3089) );
  OAI22_X1 U1896 ( .A1(n15), .A2(n3446), .B1(n226), .B2(n420), .ZN(n3090) );
  OAI22_X1 U1897 ( .A1(n376), .A2(n558), .B1(n225), .B2(n419), .ZN(n3091) );
  OAI22_X1 U1898 ( .A1(n681), .A2(n697), .B1(n225), .B2(n418), .ZN(n3092) );
  OAI22_X1 U1899 ( .A1(n272), .A2(n559), .B1(n225), .B2(n417), .ZN(n3093) );
  OAI22_X1 U1900 ( .A1(n253), .A2(n737), .B1(n3376), .B2(n152), .ZN(n3166) );
  OAI22_X1 U1901 ( .A1(n369), .A2(n3372), .B1(n3376), .B2(n151), .ZN(n3167) );
  OAI22_X1 U1902 ( .A1(n758), .A2(n3373), .B1(n3377), .B2(n150), .ZN(n3168) );
  OAI22_X1 U1903 ( .A1(n790), .A2(n737), .B1(n3377), .B2(n149), .ZN(n3169) );
  OAI22_X1 U1904 ( .A1(n787), .A2(n736), .B1(n3377), .B2(n148), .ZN(n3170) );
  OAI22_X1 U1905 ( .A1(n785), .A2(n3374), .B1(n3377), .B2(n147), .ZN(n3171) );
  OAI22_X1 U1906 ( .A1(n782), .A2(n3374), .B1(n3377), .B2(n146), .ZN(n3172) );
  OAI22_X1 U1907 ( .A1(n779), .A2(n736), .B1(n3378), .B2(n145), .ZN(n3173) );
  OAI22_X1 U1908 ( .A1(n776), .A2(n737), .B1(n3378), .B2(n144), .ZN(n3174) );
  OAI22_X1 U1909 ( .A1(n773), .A2(n736), .B1(n3378), .B2(n143), .ZN(n3175) );
  OAI22_X1 U1910 ( .A1(n770), .A2(n3372), .B1(n3378), .B2(n142), .ZN(n3176) );
  OAI22_X1 U1911 ( .A1(n192), .A2(n737), .B1(n3378), .B2(n141), .ZN(n3177) );
  OAI22_X1 U1912 ( .A1(n688), .A2(n3373), .B1(n3379), .B2(n140), .ZN(n3178) );
  OAI22_X1 U1913 ( .A1(n10), .A2(n737), .B1(n3379), .B2(n139), .ZN(n3179) );
  OAI22_X1 U1914 ( .A1(n607), .A2(n737), .B1(n3379), .B2(n138), .ZN(n3180) );
  OAI22_X1 U1915 ( .A1(n285), .A2(n3374), .B1(n3379), .B2(n137), .ZN(n3181) );
  OAI22_X1 U1916 ( .A1(n166), .A2(n3374), .B1(n3379), .B2(n136), .ZN(n3182) );
  OAI22_X1 U1917 ( .A1(n283), .A2(n3373), .B1(n3380), .B2(n135), .ZN(n3183) );
  OAI22_X1 U1918 ( .A1(n685), .A2(n3373), .B1(n3380), .B2(n134), .ZN(n3184) );
  OAI22_X1 U1919 ( .A1(n4184), .A2(n737), .B1(n3380), .B2(n133), .ZN(n3185) );
  OAI22_X1 U1920 ( .A1(n682), .A2(n3372), .B1(n3380), .B2(n132), .ZN(n3186) );
  OAI22_X1 U1921 ( .A1(n377), .A2(n3372), .B1(n3380), .B2(n131), .ZN(n3187) );
  OAI22_X1 U1922 ( .A1(n247), .A2(n736), .B1(n3381), .B2(n130), .ZN(n3188) );
  OAI22_X1 U1923 ( .A1(n272), .A2(n3374), .B1(n3381), .B2(n129), .ZN(n3189) );
  OAI22_X1 U1924 ( .A1(n4203), .A2(n578), .B1(n3366), .B2(n120), .ZN(n3198) );
  OAI22_X1 U1925 ( .A1(n369), .A2(n3363), .B1(n3366), .B2(n119), .ZN(n3199) );
  OAI22_X1 U1926 ( .A1(n759), .A2(n734), .B1(n3367), .B2(n118), .ZN(n3200) );
  OAI22_X1 U1927 ( .A1(n789), .A2(n734), .B1(n3367), .B2(n117), .ZN(n3201) );
  OAI22_X1 U1928 ( .A1(n786), .A2(n733), .B1(n3367), .B2(n116), .ZN(n3202) );
  OAI22_X1 U1929 ( .A1(n784), .A2(n3364), .B1(n3367), .B2(n115), .ZN(n3203) );
  OAI22_X1 U1930 ( .A1(n781), .A2(n578), .B1(n3367), .B2(n114), .ZN(n3204) );
  OAI22_X1 U1931 ( .A1(n778), .A2(n733), .B1(n3368), .B2(n113), .ZN(n3205) );
  OAI22_X1 U1932 ( .A1(n775), .A2(n734), .B1(n3368), .B2(n112), .ZN(n3206) );
  OAI22_X1 U1933 ( .A1(n772), .A2(n578), .B1(n3368), .B2(n111), .ZN(n3207) );
  OAI22_X1 U1934 ( .A1(n769), .A2(n3364), .B1(n3368), .B2(n110), .ZN(n3208) );
  OAI22_X1 U1935 ( .A1(n677), .A2(n734), .B1(n3368), .B2(n109), .ZN(n3209) );
  OAI22_X1 U1936 ( .A1(n172), .A2(n578), .B1(n3369), .B2(n108), .ZN(n3210) );
  OAI22_X1 U1937 ( .A1(n744), .A2(n578), .B1(n3369), .B2(n107), .ZN(n3211) );
  OAI22_X1 U1938 ( .A1(n608), .A2(n733), .B1(n3369), .B2(n106), .ZN(n3212) );
  OAI22_X1 U1939 ( .A1(n286), .A2(n3364), .B1(n3369), .B2(n105), .ZN(n3213) );
  OAI22_X1 U1940 ( .A1(n686), .A2(n733), .B1(n3369), .B2(n104), .ZN(n3214) );
  OAI22_X1 U1941 ( .A1(n283), .A2(n3364), .B1(n3370), .B2(n103), .ZN(n3215) );
  OAI22_X1 U1942 ( .A1(n684), .A2(n3363), .B1(n3370), .B2(n102), .ZN(n3216) );
  OAI22_X1 U1943 ( .A1(n25), .A2(n578), .B1(n3370), .B2(n101), .ZN(n3217) );
  OAI22_X1 U1944 ( .A1(n15), .A2(n3364), .B1(n3370), .B2(n100), .ZN(n3218) );
  OAI22_X1 U1945 ( .A1(n378), .A2(n734), .B1(n3370), .B2(n99), .ZN(n3219) );
  OAI22_X1 U1946 ( .A1(n247), .A2(n733), .B1(n3371), .B2(n98), .ZN(n3220) );
  OAI22_X1 U1947 ( .A1(n5), .A2(n3364), .B1(n3371), .B2(n97), .ZN(n3221) );
  OAI22_X1 U1948 ( .A1(n4203), .A2(n555), .B1(n223), .B2(n536), .ZN(n2974) );
  OAI22_X1 U1949 ( .A1(n368), .A2(n723), .B1(n3473), .B2(n535), .ZN(n2975) );
  OAI22_X1 U1950 ( .A1(n758), .A2(n555), .B1(n3473), .B2(n534), .ZN(n2976) );
  OAI22_X1 U1951 ( .A1(n723), .A2(n790), .B1(n205), .B2(n533), .ZN(n2977) );
  OAI22_X1 U1952 ( .A1(n787), .A2(n722), .B1(n3470), .B2(n532), .ZN(n2978) );
  OAI22_X1 U1953 ( .A1(n785), .A2(n3469), .B1(n3475), .B2(n531), .ZN(n2979) );
  OAI22_X1 U1954 ( .A1(n782), .A2(n3468), .B1(n212), .B2(n530), .ZN(n2980) );
  OAI22_X1 U1955 ( .A1(n556), .A2(n779), .B1(n224), .B2(n529), .ZN(n2981) );
  OAI22_X1 U1956 ( .A1(n776), .A2(n555), .B1(n3473), .B2(n528), .ZN(n2982) );
  OAI22_X1 U1957 ( .A1(n773), .A2(n3469), .B1(n223), .B2(n527), .ZN(n2983) );
  OAI22_X1 U1958 ( .A1(n770), .A2(n412), .B1(n3475), .B2(n526), .ZN(n2984) );
  OAI22_X1 U1959 ( .A1(n4192), .A2(n556), .B1(n3470), .B2(n525), .ZN(n2985) );
  OAI22_X1 U1960 ( .A1(n687), .A2(n3469), .B1(n223), .B2(n524), .ZN(n2986) );
  OAI22_X1 U1961 ( .A1(n4190), .A2(n722), .B1(n3473), .B2(n523), .ZN(n2987) );
  OAI22_X1 U1962 ( .A1(n3468), .A2(n607), .B1(n179), .B2(n522), .ZN(n2988) );
  OAI22_X1 U1963 ( .A1(n286), .A2(n555), .B1(n3473), .B2(n521), .ZN(n2989) );
  OAI22_X1 U1964 ( .A1(n686), .A2(n722), .B1(n3470), .B2(n520), .ZN(n2990) );
  OAI22_X1 U1965 ( .A1(n284), .A2(n3468), .B1(n224), .B2(n519), .ZN(n2991) );
  OAI22_X1 U1966 ( .A1(n171), .A2(n412), .B1(n3475), .B2(n518), .ZN(n2992) );
  OAI22_X1 U1967 ( .A1(n24), .A2(n722), .B1(n212), .B2(n517), .ZN(n2993) );
  OAI22_X1 U1968 ( .A1(n16), .A2(n3468), .B1(n224), .B2(n516), .ZN(n2994) );
  OAI22_X1 U1969 ( .A1(n377), .A2(n3468), .B1(n3473), .B2(n515), .ZN(n2995) );
  OAI22_X1 U1970 ( .A1(n680), .A2(n723), .B1(n3475), .B2(n514), .ZN(n2996) );
  OAI22_X1 U1971 ( .A1(n272), .A2(n412), .B1(n3475), .B2(n513), .ZN(n2997) );
  OAI22_X1 U1972 ( .A1(n689), .A2(n3425), .B1(n3428), .B2(n344), .ZN(n3102) );
  OAI22_X1 U1973 ( .A1(n368), .A2(n3423), .B1(n3427), .B2(n343), .ZN(n3103) );
  OAI22_X1 U1974 ( .A1(n759), .A2(n570), .B1(n3427), .B2(n342), .ZN(n3104) );
  OAI22_X1 U1975 ( .A1(n169), .A2(n726), .B1(n3429), .B2(n341), .ZN(n3105) );
  OAI22_X1 U1976 ( .A1(n571), .A2(n786), .B1(n3431), .B2(n340), .ZN(n3106) );
  OAI22_X1 U1977 ( .A1(n784), .A2(n3425), .B1(n174), .B2(n339), .ZN(n3107) );
  OAI22_X1 U1978 ( .A1(n781), .A2(n570), .B1(n3430), .B2(n338), .ZN(n3108) );
  OAI22_X1 U1979 ( .A1(n778), .A2(n3423), .B1(n3429), .B2(n337), .ZN(n3109) );
  OAI22_X1 U1980 ( .A1(n775), .A2(n726), .B1(n3431), .B2(n336), .ZN(n3110) );
  OAI22_X1 U1981 ( .A1(n772), .A2(n571), .B1(n3430), .B2(n335), .ZN(n3111) );
  OAI22_X1 U1982 ( .A1(n769), .A2(n3423), .B1(n3427), .B2(n334), .ZN(n3112) );
  OAI22_X1 U1983 ( .A1(n677), .A2(n726), .B1(n174), .B2(n333), .ZN(n3113) );
  OAI22_X1 U1984 ( .A1(n688), .A2(n571), .B1(n174), .B2(n332), .ZN(n3114) );
  OAI22_X1 U1985 ( .A1(n10), .A2(n726), .B1(n3428), .B2(n331), .ZN(n3115) );
  OAI22_X1 U1986 ( .A1(n608), .A2(n726), .B1(n3429), .B2(n330), .ZN(n3116) );
  OAI22_X1 U1987 ( .A1(n3424), .A2(n286), .B1(n3431), .B2(n329), .ZN(n3117) );
  OAI22_X1 U1988 ( .A1(n686), .A2(n3424), .B1(n3430), .B2(n328), .ZN(n3118) );
  OAI22_X1 U1989 ( .A1(n284), .A2(n571), .B1(n3428), .B2(n327), .ZN(n3119) );
  OAI22_X1 U1990 ( .A1(n4185), .A2(n571), .B1(n326), .B2(n3429), .ZN(n3120) );
  OAI22_X1 U1991 ( .A1(n4184), .A2(n570), .B1(n270), .B2(n325), .ZN(n3121) );
  OAI22_X1 U1992 ( .A1(n16), .A2(n3423), .B1(n324), .B2(n174), .ZN(n3122) );
  OAI22_X1 U1993 ( .A1(n378), .A2(n570), .B1(n3430), .B2(n323), .ZN(n3123) );
  OAI22_X1 U1994 ( .A1(n4181), .A2(n3425), .B1(n270), .B2(n322), .ZN(n3124) );
  OAI22_X1 U1995 ( .A1(n713), .A2(n3424), .B1(n270), .B2(n321), .ZN(n3125) );
  OAI22_X1 U1996 ( .A1(n689), .A2(n3413), .B1(n3417), .B2(n312), .ZN(n3134) );
  OAI22_X1 U1997 ( .A1(n368), .A2(n569), .B1(n3419), .B2(n311), .ZN(n3135) );
  OAI22_X1 U1998 ( .A1(n758), .A2(n569), .B1(n3419), .B2(n310), .ZN(n3136) );
  OAI22_X1 U1999 ( .A1(n169), .A2(n3415), .B1(n3421), .B2(n309), .ZN(n3137) );
  OAI22_X1 U2000 ( .A1(n787), .A2(n3413), .B1(n3418), .B2(n308), .ZN(n3138) );
  OAI22_X1 U2001 ( .A1(n785), .A2(n3415), .B1(n3420), .B2(n307), .ZN(n3139) );
  OAI22_X1 U2002 ( .A1(n782), .A2(n176), .B1(n3420), .B2(n306), .ZN(n3140) );
  OAI22_X1 U2003 ( .A1(n779), .A2(n3414), .B1(n3419), .B2(n305), .ZN(n3141) );
  OAI22_X1 U2004 ( .A1(n776), .A2(n742), .B1(n3421), .B2(n304), .ZN(n3142) );
  OAI22_X1 U2005 ( .A1(n773), .A2(n568), .B1(n3418), .B2(n303), .ZN(n3143) );
  OAI22_X1 U2006 ( .A1(n770), .A2(n568), .B1(n3420), .B2(n302), .ZN(n3144) );
  OAI22_X1 U2007 ( .A1(n4192), .A2(n743), .B1(n3417), .B2(n301), .ZN(n3145) );
  OAI22_X1 U2008 ( .A1(n172), .A2(n742), .B1(n3417), .B2(n300), .ZN(n3146) );
  OAI22_X1 U2009 ( .A1(n744), .A2(n569), .B1(n3419), .B2(n299), .ZN(n3147) );
  OAI22_X1 U2010 ( .A1(n607), .A2(n3413), .B1(n3421), .B2(n298), .ZN(n3148) );
  OAI22_X1 U2011 ( .A1(n286), .A2(n569), .B1(n3418), .B2(n297), .ZN(n3149) );
  OAI22_X1 U2012 ( .A1(n167), .A2(n743), .B1(n3420), .B2(n296), .ZN(n3150) );
  OAI22_X1 U2013 ( .A1(n283), .A2(n176), .B1(n3419), .B2(n295), .ZN(n3151) );
  OAI22_X1 U2014 ( .A1(n685), .A2(n743), .B1(n3421), .B2(n294), .ZN(n3152) );
  OAI22_X1 U2015 ( .A1(n25), .A2(n568), .B1(n3418), .B2(n293), .ZN(n3153) );
  OAI22_X1 U2016 ( .A1(n16), .A2(n743), .B1(n3420), .B2(n292), .ZN(n3154) );
  OAI22_X1 U2017 ( .A1(n377), .A2(n3414), .B1(n3417), .B2(n291), .ZN(n3155) );
  OAI22_X1 U2018 ( .A1(n3415), .A2(n681), .B1(n3422), .B2(n290), .ZN(n3156) );
  OAI22_X1 U2019 ( .A1(n568), .A2(n4180), .B1(n3422), .B2(n289), .ZN(n3157) );
  OAI22_X1 U2020 ( .A1(n689), .A2(n567), .B1(n3357), .B2(n88), .ZN(n3230) );
  OAI22_X1 U2021 ( .A1(n369), .A2(n566), .B1(n3357), .B2(n87), .ZN(n3231) );
  OAI22_X1 U2022 ( .A1(n759), .A2(n739), .B1(n3359), .B2(n86), .ZN(n3232) );
  OAI22_X1 U2023 ( .A1(n790), .A2(n739), .B1(n269), .B2(n85), .ZN(n3233) );
  OAI22_X1 U2024 ( .A1(n786), .A2(n3355), .B1(n3358), .B2(n84), .ZN(n3234) );
  OAI22_X1 U2025 ( .A1(n784), .A2(n3355), .B1(n22), .B2(n83), .ZN(n3235) );
  OAI22_X1 U2026 ( .A1(n781), .A2(n3353), .B1(n3360), .B2(n82), .ZN(n3236) );
  OAI22_X1 U2027 ( .A1(n778), .A2(n566), .B1(n175), .B2(n81), .ZN(n3237) );
  OAI22_X1 U2028 ( .A1(n775), .A2(n3353), .B1(n3358), .B2(n80), .ZN(n3238) );
  OAI22_X1 U2029 ( .A1(n772), .A2(n3354), .B1(n22), .B2(n79), .ZN(n3239) );
  OAI22_X1 U2030 ( .A1(n769), .A2(n739), .B1(n3359), .B2(n78), .ZN(n3240) );
  OAI22_X1 U2031 ( .A1(n192), .A2(n566), .B1(n22), .B2(n77), .ZN(n3241) );
  OAI22_X1 U2032 ( .A1(n4191), .A2(n3354), .B1(n175), .B2(n76), .ZN(n3242) );
  OAI22_X1 U2033 ( .A1(n744), .A2(n566), .B1(n269), .B2(n75), .ZN(n3243) );
  OAI22_X1 U2034 ( .A1(n608), .A2(n3353), .B1(n269), .B2(n74), .ZN(n3244) );
  OAI22_X1 U2035 ( .A1(n3355), .A2(n287), .B1(n3358), .B2(n73), .ZN(n3245) );
  OAI22_X1 U2036 ( .A1(n166), .A2(n3355), .B1(n3360), .B2(n72), .ZN(n3246) );
  OAI22_X1 U2037 ( .A1(n283), .A2(n3354), .B1(n3359), .B2(n71), .ZN(n3247) );
  OAI22_X1 U2038 ( .A1(n684), .A2(n3354), .B1(n70), .B2(n3361), .ZN(n3248) );
  OAI22_X1 U2039 ( .A1(n25), .A2(n739), .B1(n3358), .B2(n69), .ZN(n3249) );
  OAI22_X1 U2040 ( .A1(n683), .A2(n3353), .B1(n175), .B2(n68), .ZN(n3250) );
  OAI22_X1 U2041 ( .A1(n378), .A2(n566), .B1(n3360), .B2(n67), .ZN(n3251) );
  OAI22_X1 U2042 ( .A1(n680), .A2(n567), .B1(n269), .B2(n66), .ZN(n3252) );
  OAI22_X1 U2043 ( .A1(n6), .A2(n567), .B1(n3361), .B2(n65), .ZN(n3253) );
  OAI22_X1 U2044 ( .A1(n253), .A2(n565), .B1(n3349), .B2(n56), .ZN(n3262) );
  OAI22_X1 U2045 ( .A1(n369), .A2(n3343), .B1(n3348), .B2(n55), .ZN(n3263) );
  OAI22_X1 U2046 ( .A1(n758), .A2(n3344), .B1(n3349), .B2(n54), .ZN(n3264) );
  OAI22_X1 U2047 ( .A1(n169), .A2(n741), .B1(n3349), .B2(n53), .ZN(n3265) );
  OAI22_X1 U2048 ( .A1(n787), .A2(n740), .B1(n3349), .B2(n52), .ZN(n3266) );
  OAI22_X1 U2049 ( .A1(n785), .A2(n3345), .B1(n3349), .B2(n51), .ZN(n3267) );
  OAI22_X1 U2050 ( .A1(n782), .A2(n564), .B1(n3349), .B2(n50), .ZN(n3268) );
  OAI22_X1 U2051 ( .A1(n779), .A2(n740), .B1(n3347), .B2(n49), .ZN(n3269) );
  OAI22_X1 U2052 ( .A1(n776), .A2(n741), .B1(n3348), .B2(n48), .ZN(n3270) );
  OAI22_X1 U2053 ( .A1(n773), .A2(n740), .B1(n3351), .B2(n47), .ZN(n3271) );
  OAI22_X1 U2054 ( .A1(n770), .A2(n3343), .B1(n3347), .B2(n46), .ZN(n3272) );
  OAI22_X1 U2055 ( .A1(n192), .A2(n741), .B1(n3347), .B2(n45), .ZN(n3273) );
  OAI22_X1 U2056 ( .A1(n172), .A2(n3344), .B1(n3350), .B2(n44), .ZN(n3274) );
  OAI22_X1 U2057 ( .A1(n4190), .A2(n741), .B1(n3350), .B2(n43), .ZN(n3275) );
  OAI22_X1 U2058 ( .A1(n607), .A2(n741), .B1(n3350), .B2(n42), .ZN(n3276) );
  OAI22_X1 U2059 ( .A1(n286), .A2(n3345), .B1(n3350), .B2(n41), .ZN(n3277) );
  OAI22_X1 U2060 ( .A1(n167), .A2(n3345), .B1(n3350), .B2(n40), .ZN(n3278) );
  OAI22_X1 U2061 ( .A1(n283), .A2(n3344), .B1(n3348), .B2(n39), .ZN(n3279) );
  OAI22_X1 U2062 ( .A1(n4185), .A2(n3344), .B1(n3351), .B2(n38), .ZN(n3280) );
  OAI22_X1 U2063 ( .A1(n271), .A2(n564), .B1(n3348), .B2(n37), .ZN(n3281) );
  OAI22_X1 U2064 ( .A1(n15), .A2(n3343), .B1(n3351), .B2(n36), .ZN(n3282) );
  OAI22_X1 U2065 ( .A1(n378), .A2(n564), .B1(n3351), .B2(n35), .ZN(n3283) );
  OAI22_X1 U2066 ( .A1(n247), .A2(n740), .B1(n3352), .B2(n34), .ZN(n3284) );
  OAI22_X1 U2067 ( .A1(n713), .A2(n565), .B1(n3351), .B2(n33), .ZN(n3285) );
  OAI22_X1 U2068 ( .A1(n693), .A2(n674), .B1(n29), .B2(n959), .ZN(n2807) );
  OAI22_X1 U2069 ( .A1(n4209), .A2(n560), .B1(n241), .B2(n958), .ZN(n2808) );
  OAI22_X1 U2070 ( .A1(n691), .A2(n3573), .B1(n240), .B2(n957), .ZN(n2809) );
  OAI22_X1 U2071 ( .A1(n355), .A2(n560), .B1(n241), .B2(n956), .ZN(n2810) );
  OAI22_X1 U2072 ( .A1(n4206), .A2(n410), .B1(n29), .B2(n955), .ZN(n2811) );
  OAI22_X1 U2073 ( .A1(n170), .A2(n560), .B1(n239), .B2(n954), .ZN(n2812) );
  OAI22_X1 U2074 ( .A1(n4204), .A2(n3574), .B1(n29), .B2(n953), .ZN(n2813) );
  OAI22_X1 U2075 ( .A1(n4211), .A2(n728), .B1(n3551), .B2(n864), .ZN(n2838) );
  OAI22_X1 U2076 ( .A1(n4210), .A2(n727), .B1(n3551), .B2(n863), .ZN(n2839) );
  OAI22_X1 U2077 ( .A1(n4209), .A2(n3550), .B1(n3551), .B2(n862), .ZN(n2840)
         );
  OAI22_X1 U2078 ( .A1(n4208), .A2(n3548), .B1(n3551), .B2(n861), .ZN(n2841)
         );
  OAI22_X1 U2079 ( .A1(n355), .A2(n728), .B1(n3551), .B2(n860), .ZN(n2842) );
  OAI22_X1 U2080 ( .A1(n4206), .A2(n727), .B1(n3552), .B2(n859), .ZN(n2843) );
  OAI22_X1 U2081 ( .A1(n4205), .A2(n3550), .B1(n3552), .B2(n858), .ZN(n2844)
         );
  OAI22_X1 U2082 ( .A1(n248), .A2(n3548), .B1(n3552), .B2(n857), .ZN(n2845) );
  OAI22_X1 U2083 ( .A1(n4211), .A2(n731), .B1(n3542), .B2(n832), .ZN(n2870) );
  OAI22_X1 U2084 ( .A1(n694), .A2(n572), .B1(n3545), .B2(n831), .ZN(n2871) );
  OAI22_X1 U2085 ( .A1(n4209), .A2(n3539), .B1(n3544), .B2(n830), .ZN(n2872)
         );
  OAI22_X1 U2086 ( .A1(n279), .A2(n731), .B1(n3543), .B2(n829), .ZN(n2873) );
  OAI22_X1 U2087 ( .A1(n357), .A2(n3538), .B1(n3544), .B2(n828), .ZN(n2874) );
  OAI22_X1 U2088 ( .A1(n678), .A2(n3540), .B1(n3541), .B2(n827), .ZN(n2875) );
  OAI22_X1 U2089 ( .A1(n715), .A2(n3540), .B1(n3545), .B2(n826), .ZN(n2876) );
  OAI22_X1 U2090 ( .A1(n690), .A2(n572), .B1(n3546), .B2(n825), .ZN(n2877) );
  OAI22_X1 U2091 ( .A1(n4211), .A2(n738), .B1(n3508), .B2(n672), .ZN(n2902) );
  OAI22_X1 U2092 ( .A1(n693), .A2(n3502), .B1(n3510), .B2(n671), .ZN(n2903) );
  OAI22_X1 U2093 ( .A1(n4209), .A2(n738), .B1(n3506), .B2(n670), .ZN(n2904) );
  OAI22_X1 U2094 ( .A1(n279), .A2(n3502), .B1(n3507), .B2(n669), .ZN(n2905) );
  OAI22_X1 U2095 ( .A1(n356), .A2(n577), .B1(n3505), .B2(n668), .ZN(n2906) );
  OAI22_X1 U2096 ( .A1(n3503), .A2(n679), .B1(n3509), .B2(n667), .ZN(n2907) );
  OAI22_X1 U2097 ( .A1(n8), .A2(n3504), .B1(n3507), .B2(n666), .ZN(n2908) );
  OAI22_X1 U2098 ( .A1(n248), .A2(n3503), .B1(n3505), .B2(n665), .ZN(n2909) );
  OAI22_X1 U2099 ( .A1(n766), .A2(n735), .B1(n3499), .B2(n640), .ZN(n2934) );
  OAI22_X1 U2100 ( .A1(n4210), .A2(n3493), .B1(n3498), .B2(n639), .ZN(n2935)
         );
  OAI22_X1 U2101 ( .A1(n4209), .A2(n3493), .B1(n3497), .B2(n638), .ZN(n2936)
         );
  OAI22_X1 U2102 ( .A1(n280), .A2(n735), .B1(n359), .B2(n637), .ZN(n2937) );
  OAI22_X1 U2103 ( .A1(n356), .A2(n3494), .B1(n3500), .B2(n636), .ZN(n2938) );
  OAI22_X1 U2104 ( .A1(n3493), .A2(n678), .B1(n3500), .B2(n635), .ZN(n2939) );
  OAI22_X1 U2105 ( .A1(n8), .A2(n3493), .B1(n3499), .B2(n634), .ZN(n2940) );
  OAI22_X1 U2106 ( .A1(n249), .A2(n735), .B1(n3496), .B2(n633), .ZN(n2941) );
  OAI22_X1 U2107 ( .A1(n766), .A2(n372), .B1(n3452), .B2(n480), .ZN(n3030) );
  OAI22_X1 U2108 ( .A1(n187), .A2(n372), .B1(n3452), .B2(n479), .ZN(n3031) );
  OAI22_X1 U2109 ( .A1(n4209), .A2(n593), .B1(n3452), .B2(n478), .ZN(n3032) );
  OAI22_X1 U2110 ( .A1(n4208), .A2(n593), .B1(n3452), .B2(n477), .ZN(n3033) );
  OAI22_X1 U2111 ( .A1(n356), .A2(n372), .B1(n3452), .B2(n476), .ZN(n3034) );
  OAI22_X1 U2112 ( .A1(n678), .A2(n3451), .B1(n3453), .B2(n475), .ZN(n3035) );
  OAI22_X1 U2113 ( .A1(n715), .A2(n594), .B1(n3453), .B2(n474), .ZN(n3036) );
  OAI22_X1 U2114 ( .A1(n249), .A2(n593), .B1(n3453), .B2(n473), .ZN(n3037) );
  OAI22_X1 U2115 ( .A1(n767), .A2(n559), .B1(n226), .B2(n448), .ZN(n3062) );
  OAI22_X1 U2116 ( .A1(n4209), .A2(n697), .B1(n3448), .B2(n446), .ZN(n3064) );
  OAI22_X1 U2117 ( .A1(n280), .A2(n3446), .B1(n226), .B2(n445), .ZN(n3065) );
  OAI22_X1 U2118 ( .A1(n356), .A2(n558), .B1(n225), .B2(n444), .ZN(n3066) );
  OAI22_X1 U2119 ( .A1(n4206), .A2(n559), .B1(n226), .B2(n443), .ZN(n3067) );
  OAI22_X1 U2120 ( .A1(n9), .A2(n3446), .B1(n225), .B2(n442), .ZN(n3068) );
  OAI22_X1 U2121 ( .A1(n249), .A2(n3447), .B1(n225), .B2(n441), .ZN(n3069) );
  OAI22_X1 U2122 ( .A1(n766), .A2(n736), .B1(n3375), .B2(n160), .ZN(n3158) );
  OAI22_X1 U2123 ( .A1(n188), .A2(n3372), .B1(n3375), .B2(n159), .ZN(n3159) );
  OAI22_X1 U2124 ( .A1(n4209), .A2(n736), .B1(n3375), .B2(n158), .ZN(n3160) );
  OAI22_X1 U2125 ( .A1(n4208), .A2(n3372), .B1(n3375), .B2(n157), .ZN(n3161)
         );
  OAI22_X1 U2126 ( .A1(n356), .A2(n3373), .B1(n3375), .B2(n156), .ZN(n3162) );
  OAI22_X1 U2127 ( .A1(n679), .A2(n3374), .B1(n3376), .B2(n155), .ZN(n3163) );
  OAI22_X1 U2128 ( .A1(n714), .A2(n3374), .B1(n3376), .B2(n154), .ZN(n3164) );
  OAI22_X1 U2129 ( .A1(n690), .A2(n3373), .B1(n3376), .B2(n153), .ZN(n3165) );
  OAI22_X1 U2130 ( .A1(n767), .A2(n3363), .B1(n3365), .B2(n128), .ZN(n3190) );
  OAI22_X1 U2131 ( .A1(n188), .A2(n733), .B1(n3365), .B2(n127), .ZN(n3191) );
  OAI22_X1 U2132 ( .A1(n4209), .A2(n3363), .B1(n3365), .B2(n126), .ZN(n3192)
         );
  OAI22_X1 U2133 ( .A1(n280), .A2(n3363), .B1(n3365), .B2(n125), .ZN(n3193) );
  OAI22_X1 U2134 ( .A1(n357), .A2(n3363), .B1(n3365), .B2(n124), .ZN(n3194) );
  OAI22_X1 U2135 ( .A1(n4206), .A2(n734), .B1(n3366), .B2(n123), .ZN(n3195) );
  OAI22_X1 U2136 ( .A1(n9), .A2(n734), .B1(n3366), .B2(n122), .ZN(n3196) );
  OAI22_X1 U2137 ( .A1(n4204), .A2(n3363), .B1(n3366), .B2(n121), .ZN(n3197)
         );
  OAI22_X1 U2138 ( .A1(n766), .A2(n412), .B1(n3470), .B2(n544), .ZN(n2966) );
  OAI22_X1 U2139 ( .A1(n694), .A2(n556), .B1(n205), .B2(n543), .ZN(n2967) );
  OAI22_X1 U2140 ( .A1(n4209), .A2(n556), .B1(n3470), .B2(n542), .ZN(n2968) );
  OAI22_X1 U2141 ( .A1(n280), .A2(n3468), .B1(n3475), .B2(n541), .ZN(n2969) );
  OAI22_X1 U2142 ( .A1(n357), .A2(n722), .B1(n212), .B2(n540), .ZN(n2970) );
  OAI22_X1 U2143 ( .A1(n679), .A2(n3469), .B1(n179), .B2(n539), .ZN(n2971) );
  OAI22_X1 U2144 ( .A1(n170), .A2(n412), .B1(n3470), .B2(n538), .ZN(n2972) );
  OAI22_X1 U2145 ( .A1(n249), .A2(n723), .B1(n205), .B2(n537), .ZN(n2973) );
  OAI22_X1 U2146 ( .A1(n767), .A2(n3425), .B1(n3426), .B2(n352), .ZN(n3094) );
  OAI22_X1 U2147 ( .A1(n188), .A2(n3423), .B1(n3426), .B2(n351), .ZN(n3095) );
  OAI22_X1 U2148 ( .A1(n4209), .A2(n570), .B1(n3426), .B2(n350), .ZN(n3096) );
  OAI22_X1 U2149 ( .A1(n279), .A2(n3423), .B1(n3426), .B2(n349), .ZN(n3097) );
  OAI22_X1 U2150 ( .A1(n357), .A2(n570), .B1(n270), .B2(n348), .ZN(n3098) );
  OAI22_X1 U2151 ( .A1(n678), .A2(n3424), .B1(n3427), .B2(n347), .ZN(n3099) );
  OAI22_X1 U2152 ( .A1(n3425), .A2(n4205), .B1(n3428), .B2(n346), .ZN(n3100)
         );
  OAI22_X1 U2153 ( .A1(n3424), .A2(n4204), .B1(n3427), .B2(n345), .ZN(n3101)
         );
  OAI22_X1 U2154 ( .A1(n766), .A2(n3413), .B1(n3416), .B2(n320), .ZN(n3126) );
  OAI22_X1 U2155 ( .A1(n693), .A2(n742), .B1(n3416), .B2(n319), .ZN(n3127) );
  OAI22_X1 U2156 ( .A1(n4209), .A2(n176), .B1(n3416), .B2(n318), .ZN(n3128) );
  OAI22_X1 U2157 ( .A1(n4208), .A2(n3414), .B1(n3416), .B2(n317), .ZN(n3129)
         );
  OAI22_X1 U2158 ( .A1(n355), .A2(n3414), .B1(n3416), .B2(n316), .ZN(n3130) );
  OAI22_X1 U2159 ( .A1(n679), .A2(n742), .B1(n3421), .B2(n315), .ZN(n3131) );
  OAI22_X1 U2160 ( .A1(n4205), .A2(n3415), .B1(n3418), .B2(n314), .ZN(n3132)
         );
  OAI22_X1 U2161 ( .A1(n690), .A2(n176), .B1(n3420), .B2(n313), .ZN(n3133) );
  OAI22_X1 U2162 ( .A1(n767), .A2(n567), .B1(n3357), .B2(n96), .ZN(n3222) );
  OAI22_X1 U2163 ( .A1(n187), .A2(n739), .B1(n3356), .B2(n95), .ZN(n3223) );
  OAI22_X1 U2164 ( .A1(n4209), .A2(n3353), .B1(n3356), .B2(n94), .ZN(n3224) );
  OAI22_X1 U2165 ( .A1(n280), .A2(n3353), .B1(n3356), .B2(n93), .ZN(n3225) );
  OAI22_X1 U2166 ( .A1(n357), .A2(n566), .B1(n3361), .B2(n92), .ZN(n3226) );
  OAI22_X1 U2167 ( .A1(n678), .A2(n567), .B1(n3357), .B2(n91), .ZN(n3227) );
  OAI22_X1 U2168 ( .A1(n170), .A2(n3355), .B1(n3357), .B2(n90), .ZN(n3228) );
  OAI22_X1 U2169 ( .A1(n690), .A2(n3354), .B1(n3357), .B2(n89), .ZN(n3229) );
  OAI22_X1 U2170 ( .A1(n766), .A2(n565), .B1(n3346), .B2(n64), .ZN(n3254) );
  OAI22_X1 U2171 ( .A1(n694), .A2(n3343), .B1(n3346), .B2(n63), .ZN(n3255) );
  OAI22_X1 U2172 ( .A1(n4209), .A2(n740), .B1(n3346), .B2(n62), .ZN(n3256) );
  OAI22_X1 U2173 ( .A1(n279), .A2(n3343), .B1(n3346), .B2(n61), .ZN(n3257) );
  OAI22_X1 U2174 ( .A1(n356), .A2(n564), .B1(n3346), .B2(n60), .ZN(n3258) );
  OAI22_X1 U2175 ( .A1(n678), .A2(n565), .B1(n3351), .B2(n59), .ZN(n3259) );
  OAI22_X1 U2176 ( .A1(n9), .A2(n3345), .B1(n3347), .B2(n58), .ZN(n3260) );
  OAI22_X1 U2177 ( .A1(n248), .A2(n3344), .B1(n3351), .B2(n57), .ZN(n3261) );
  OAI22_X1 U2178 ( .A1(n253), .A2(n3459), .B1(n3462), .B2(n504), .ZN(n3006) );
  OAI22_X1 U2179 ( .A1(n370), .A2(n383), .B1(n3462), .B2(n503), .ZN(n3007) );
  OAI22_X1 U2180 ( .A1(n759), .A2(n3460), .B1(n3463), .B2(n502), .ZN(n3008) );
  OAI22_X1 U2181 ( .A1(n789), .A2(n605), .B1(n3463), .B2(n501), .ZN(n3009) );
  OAI22_X1 U2182 ( .A1(n787), .A2(n606), .B1(n3463), .B2(n500), .ZN(n3010) );
  OAI22_X1 U2183 ( .A1(n785), .A2(n3459), .B1(n3463), .B2(n499), .ZN(n3011) );
  OAI22_X1 U2184 ( .A1(n782), .A2(n383), .B1(n3463), .B2(n498), .ZN(n3012) );
  OAI22_X1 U2185 ( .A1(n779), .A2(n383), .B1(n3464), .B2(n497), .ZN(n3013) );
  OAI22_X1 U2186 ( .A1(n776), .A2(n606), .B1(n3464), .B2(n496), .ZN(n3014) );
  OAI22_X1 U2187 ( .A1(n773), .A2(n605), .B1(n3464), .B2(n495), .ZN(n3015) );
  OAI22_X1 U2188 ( .A1(n770), .A2(n605), .B1(n3464), .B2(n494), .ZN(n3016) );
  OAI22_X1 U2189 ( .A1(n192), .A2(n273), .B1(n3464), .B2(n493), .ZN(n3017) );
  OAI22_X1 U2190 ( .A1(n688), .A2(n605), .B1(n3465), .B2(n492), .ZN(n3018) );
  OAI22_X1 U2191 ( .A1(n10), .A2(n3460), .B1(n3465), .B2(n491), .ZN(n3019) );
  OAI22_X1 U2192 ( .A1(n608), .A2(n3459), .B1(n3465), .B2(n490), .ZN(n3020) );
  OAI22_X1 U2193 ( .A1(n285), .A2(n605), .B1(n3465), .B2(n489), .ZN(n3021) );
  OAI22_X1 U2194 ( .A1(n166), .A2(n606), .B1(n3465), .B2(n488), .ZN(n3022) );
  OAI22_X1 U2195 ( .A1(n282), .A2(n383), .B1(n3466), .B2(n487), .ZN(n3023) );
  OAI22_X1 U2196 ( .A1(n171), .A2(n606), .B1(n3466), .B2(n486), .ZN(n3024) );
  OAI22_X1 U2197 ( .A1(n24), .A2(n606), .B1(n3466), .B2(n485), .ZN(n3025) );
  OAI22_X1 U2198 ( .A1(n682), .A2(n3460), .B1(n3466), .B2(n484), .ZN(n3026) );
  OAI22_X1 U2199 ( .A1(n376), .A2(n605), .B1(n3466), .B2(n483), .ZN(n3027) );
  OAI22_X1 U2200 ( .A1(n4181), .A2(n3459), .B1(n3463), .B2(n482), .ZN(n3028)
         );
  OAI22_X1 U2201 ( .A1(n713), .A2(n3460), .B1(n3467), .B2(n481), .ZN(n3029) );
  OAI22_X1 U2202 ( .A1(n767), .A2(n383), .B1(n3461), .B2(n512), .ZN(n2998) );
  OAI22_X1 U2203 ( .A1(n187), .A2(n3459), .B1(n3461), .B2(n511), .ZN(n2999) );
  OAI22_X1 U2204 ( .A1(n4209), .A2(n383), .B1(n3461), .B2(n510), .ZN(n3000) );
  OAI22_X1 U2205 ( .A1(n4208), .A2(n273), .B1(n3461), .B2(n509), .ZN(n3001) );
  OAI22_X1 U2206 ( .A1(n355), .A2(n3459), .B1(n3461), .B2(n508), .ZN(n3002) );
  OAI22_X1 U2207 ( .A1(n4206), .A2(n606), .B1(n3462), .B2(n507), .ZN(n3003) );
  OAI22_X1 U2208 ( .A1(n714), .A2(n3460), .B1(n3462), .B2(n506), .ZN(n3004) );
  OAI22_X1 U2209 ( .A1(n248), .A2(n3460), .B1(n3462), .B2(n505), .ZN(n3005) );
  AOI22_X1 U2210 ( .A1(n3318), .A2(\registers[23][22] ), .B1(n3315), .B2(
        \registers[22][22] ), .ZN(n1785) );
  AOI22_X1 U2211 ( .A1(n3318), .A2(\registers[23][23] ), .B1(n3315), .B2(
        \registers[22][23] ), .ZN(n1768) );
  AOI22_X1 U2212 ( .A1(n3318), .A2(\registers[23][24] ), .B1(n3315), .B2(
        \registers[22][24] ), .ZN(n1751) );
  AOI22_X1 U2213 ( .A1(n3318), .A2(\registers[23][25] ), .B1(n3315), .B2(
        \registers[22][25] ), .ZN(n1734) );
  AOI22_X1 U2214 ( .A1(n3318), .A2(\registers[23][26] ), .B1(n3315), .B2(
        \registers[22][26] ), .ZN(n1717) );
  AOI22_X1 U2215 ( .A1(n3318), .A2(\registers[23][27] ), .B1(n3315), .B2(
        \registers[22][27] ), .ZN(n1700) );
  AOI22_X1 U2216 ( .A1(n3318), .A2(\registers[23][28] ), .B1(n3315), .B2(
        \registers[22][28] ), .ZN(n1683) );
  AOI22_X1 U2217 ( .A1(n3318), .A2(\registers[23][29] ), .B1(n3315), .B2(
        \registers[22][29] ), .ZN(n1666) );
  AOI22_X1 U2218 ( .A1(n3318), .A2(\registers[23][30] ), .B1(n3315), .B2(
        \registers[22][30] ), .ZN(n1649) );
  AOI22_X1 U2219 ( .A1(n3318), .A2(\registers[23][31] ), .B1(n3315), .B2(
        \registers[22][31] ), .ZN(n1607) );
  AOI22_X1 U2220 ( .A1(n1044), .A2(\registers[23][22] ), .B1(n1041), .B2(
        \registers[22][22] ), .ZN(n2376) );
  AOI22_X1 U2221 ( .A1(n1044), .A2(\registers[23][23] ), .B1(n1041), .B2(
        \registers[22][23] ), .ZN(n2359) );
  AOI22_X1 U2222 ( .A1(n1044), .A2(\registers[23][24] ), .B1(n1041), .B2(
        \registers[22][24] ), .ZN(n2342) );
  AOI22_X1 U2223 ( .A1(n1044), .A2(\registers[23][25] ), .B1(n1041), .B2(
        \registers[22][25] ), .ZN(n2325) );
  AOI22_X1 U2224 ( .A1(n1044), .A2(\registers[23][26] ), .B1(n1041), .B2(
        \registers[22][26] ), .ZN(n2308) );
  AOI22_X1 U2225 ( .A1(n1044), .A2(\registers[23][27] ), .B1(n1041), .B2(
        \registers[22][27] ), .ZN(n2291) );
  AOI22_X1 U2226 ( .A1(n1044), .A2(\registers[23][28] ), .B1(n1041), .B2(
        \registers[22][28] ), .ZN(n2274) );
  AOI22_X1 U2227 ( .A1(n1044), .A2(\registers[23][29] ), .B1(n1041), .B2(
        \registers[22][29] ), .ZN(n2257) );
  AOI22_X1 U2228 ( .A1(n1044), .A2(\registers[23][30] ), .B1(n1041), .B2(
        \registers[22][30] ), .ZN(n2240) );
  AOI22_X1 U2229 ( .A1(n1044), .A2(\registers[23][31] ), .B1(n1041), .B2(
        \registers[22][31] ), .ZN(n2198) );
  AOI22_X1 U2230 ( .A1(n3316), .A2(\registers[23][0] ), .B1(n3313), .B2(
        \registers[22][0] ), .ZN(n2163) );
  AOI22_X1 U2231 ( .A1(n3316), .A2(\registers[23][1] ), .B1(n3313), .B2(
        \registers[22][1] ), .ZN(n2142) );
  AOI22_X1 U2232 ( .A1(n3316), .A2(\registers[23][2] ), .B1(n3313), .B2(
        \registers[22][2] ), .ZN(n2125) );
  AOI22_X1 U2233 ( .A1(n3316), .A2(\registers[23][3] ), .B1(n3313), .B2(
        \registers[22][3] ), .ZN(n2108) );
  AOI22_X1 U2234 ( .A1(n3316), .A2(\registers[23][4] ), .B1(n3313), .B2(
        \registers[22][4] ), .ZN(n2091) );
  AOI22_X1 U2235 ( .A1(n3316), .A2(\registers[23][5] ), .B1(n3313), .B2(
        \registers[22][5] ), .ZN(n2074) );
  AOI22_X1 U2236 ( .A1(n3316), .A2(\registers[23][6] ), .B1(n3313), .B2(
        \registers[22][6] ), .ZN(n2057) );
  AOI22_X1 U2237 ( .A1(n3316), .A2(\registers[23][7] ), .B1(n3313), .B2(
        \registers[22][7] ), .ZN(n2040) );
  AOI22_X1 U2238 ( .A1(n3316), .A2(\registers[23][8] ), .B1(n3313), .B2(
        \registers[22][8] ), .ZN(n2023) );
  AOI22_X1 U2239 ( .A1(n3316), .A2(\registers[23][9] ), .B1(n3313), .B2(
        \registers[22][9] ), .ZN(n2006) );
  AOI22_X1 U2240 ( .A1(n3316), .A2(\registers[23][10] ), .B1(n3313), .B2(
        \registers[22][10] ), .ZN(n1989) );
  AOI22_X1 U2241 ( .A1(n3317), .A2(\registers[23][11] ), .B1(n3314), .B2(
        \registers[22][11] ), .ZN(n1972) );
  AOI22_X1 U2242 ( .A1(n3317), .A2(\registers[23][12] ), .B1(n3314), .B2(
        \registers[22][12] ), .ZN(n1955) );
  AOI22_X1 U2243 ( .A1(n3317), .A2(\registers[23][13] ), .B1(n3314), .B2(
        \registers[22][13] ), .ZN(n1938) );
  AOI22_X1 U2244 ( .A1(n3317), .A2(\registers[23][14] ), .B1(n3314), .B2(
        \registers[22][14] ), .ZN(n1921) );
  AOI22_X1 U2245 ( .A1(n3317), .A2(\registers[23][15] ), .B1(n3314), .B2(
        \registers[22][15] ), .ZN(n1904) );
  AOI22_X1 U2246 ( .A1(n3317), .A2(\registers[23][16] ), .B1(n3314), .B2(
        \registers[22][16] ), .ZN(n1887) );
  AOI22_X1 U2247 ( .A1(n3317), .A2(\registers[23][17] ), .B1(n3314), .B2(
        \registers[22][17] ), .ZN(n1870) );
  AOI22_X1 U2248 ( .A1(n3317), .A2(\registers[23][18] ), .B1(n3314), .B2(
        \registers[22][18] ), .ZN(n1853) );
  AOI22_X1 U2249 ( .A1(n3317), .A2(\registers[23][19] ), .B1(n3314), .B2(
        \registers[22][19] ), .ZN(n1836) );
  AOI22_X1 U2250 ( .A1(n3317), .A2(\registers[23][20] ), .B1(n3314), .B2(
        \registers[22][20] ), .ZN(n1819) );
  AOI22_X1 U2251 ( .A1(n3317), .A2(\registers[23][21] ), .B1(n3314), .B2(
        \registers[22][21] ), .ZN(n1802) );
  AOI22_X1 U2252 ( .A1(n1042), .A2(\registers[23][0] ), .B1(n1039), .B2(
        \registers[22][0] ), .ZN(n2754) );
  AOI22_X1 U2253 ( .A1(n1042), .A2(\registers[23][1] ), .B1(n1039), .B2(
        \registers[22][1] ), .ZN(n2733) );
  AOI22_X1 U2254 ( .A1(n1042), .A2(\registers[23][2] ), .B1(n1039), .B2(
        \registers[22][2] ), .ZN(n2716) );
  AOI22_X1 U2255 ( .A1(n1042), .A2(\registers[23][3] ), .B1(n1039), .B2(
        \registers[22][3] ), .ZN(n2699) );
  AOI22_X1 U2256 ( .A1(n1042), .A2(\registers[23][4] ), .B1(n1039), .B2(
        \registers[22][4] ), .ZN(n2682) );
  AOI22_X1 U2257 ( .A1(n1042), .A2(\registers[23][5] ), .B1(n1039), .B2(
        \registers[22][5] ), .ZN(n2665) );
  AOI22_X1 U2258 ( .A1(n1042), .A2(\registers[23][6] ), .B1(n1039), .B2(
        \registers[22][6] ), .ZN(n2648) );
  AOI22_X1 U2259 ( .A1(n1042), .A2(\registers[23][7] ), .B1(n1039), .B2(
        \registers[22][7] ), .ZN(n2631) );
  AOI22_X1 U2260 ( .A1(n1042), .A2(\registers[23][8] ), .B1(n1039), .B2(
        \registers[22][8] ), .ZN(n2614) );
  AOI22_X1 U2261 ( .A1(n1042), .A2(\registers[23][9] ), .B1(n1039), .B2(
        \registers[22][9] ), .ZN(n2597) );
  AOI22_X1 U2262 ( .A1(n1042), .A2(\registers[23][10] ), .B1(n1039), .B2(
        \registers[22][10] ), .ZN(n2580) );
  AOI22_X1 U2263 ( .A1(n1043), .A2(\registers[23][11] ), .B1(n1040), .B2(
        \registers[22][11] ), .ZN(n2563) );
  AOI22_X1 U2264 ( .A1(n1043), .A2(\registers[23][12] ), .B1(n1040), .B2(
        \registers[22][12] ), .ZN(n2546) );
  AOI22_X1 U2265 ( .A1(n1043), .A2(\registers[23][13] ), .B1(n1040), .B2(
        \registers[22][13] ), .ZN(n2529) );
  AOI22_X1 U2266 ( .A1(n1043), .A2(\registers[23][14] ), .B1(n1040), .B2(
        \registers[22][14] ), .ZN(n2512) );
  AOI22_X1 U2267 ( .A1(n1043), .A2(\registers[23][15] ), .B1(n1040), .B2(
        \registers[22][15] ), .ZN(n2495) );
  AOI22_X1 U2268 ( .A1(n1043), .A2(\registers[23][16] ), .B1(n1040), .B2(
        \registers[22][16] ), .ZN(n2478) );
  AOI22_X1 U2269 ( .A1(n1043), .A2(\registers[23][17] ), .B1(n1040), .B2(
        \registers[22][17] ), .ZN(n2461) );
  AOI22_X1 U2270 ( .A1(n1043), .A2(\registers[23][18] ), .B1(n1040), .B2(
        \registers[22][18] ), .ZN(n2444) );
  AOI22_X1 U2271 ( .A1(n1043), .A2(\registers[23][19] ), .B1(n1040), .B2(
        \registers[22][19] ), .ZN(n2427) );
  AOI22_X1 U2272 ( .A1(n1043), .A2(\registers[23][20] ), .B1(n1040), .B2(
        \registers[22][20] ), .ZN(n2410) );
  AOI22_X1 U2273 ( .A1(n1043), .A2(\registers[23][21] ), .B1(n1040), .B2(
        \registers[22][21] ), .ZN(n2393) );
  AOI22_X1 U2274 ( .A1(n3306), .A2(\registers[25][22] ), .B1(n3303), .B2(
        \registers[24][22] ), .ZN(n1786) );
  AOI22_X1 U2275 ( .A1(n3306), .A2(\registers[25][23] ), .B1(n3303), .B2(
        \registers[24][23] ), .ZN(n1769) );
  AOI22_X1 U2276 ( .A1(n3306), .A2(\registers[25][24] ), .B1(n3303), .B2(
        \registers[24][24] ), .ZN(n1752) );
  AOI22_X1 U2277 ( .A1(n3306), .A2(\registers[25][25] ), .B1(n3303), .B2(
        \registers[24][25] ), .ZN(n1735) );
  AOI22_X1 U2278 ( .A1(n3306), .A2(\registers[25][26] ), .B1(n3303), .B2(
        \registers[24][26] ), .ZN(n1718) );
  AOI22_X1 U2279 ( .A1(n3306), .A2(\registers[25][27] ), .B1(n3303), .B2(
        \registers[24][27] ), .ZN(n1701) );
  AOI22_X1 U2280 ( .A1(n3306), .A2(\registers[25][28] ), .B1(n3303), .B2(
        \registers[24][28] ), .ZN(n1684) );
  AOI22_X1 U2281 ( .A1(n3306), .A2(\registers[25][29] ), .B1(n3303), .B2(
        \registers[24][29] ), .ZN(n1667) );
  AOI22_X1 U2282 ( .A1(n3306), .A2(\registers[25][30] ), .B1(n3303), .B2(
        \registers[24][30] ), .ZN(n1650) );
  AOI22_X1 U2283 ( .A1(n3306), .A2(\registers[25][31] ), .B1(n3303), .B2(
        \registers[24][31] ), .ZN(n1612) );
  AOI22_X1 U2284 ( .A1(n1032), .A2(\registers[25][22] ), .B1(n1029), .B2(
        \registers[24][22] ), .ZN(n2377) );
  AOI22_X1 U2285 ( .A1(n1032), .A2(\registers[25][23] ), .B1(n1029), .B2(
        \registers[24][23] ), .ZN(n2360) );
  AOI22_X1 U2286 ( .A1(n1032), .A2(\registers[25][24] ), .B1(n1029), .B2(
        \registers[24][24] ), .ZN(n2343) );
  AOI22_X1 U2287 ( .A1(n1032), .A2(\registers[25][25] ), .B1(n1029), .B2(
        \registers[24][25] ), .ZN(n2326) );
  AOI22_X1 U2288 ( .A1(n1032), .A2(\registers[25][26] ), .B1(n1029), .B2(
        \registers[24][26] ), .ZN(n2309) );
  AOI22_X1 U2289 ( .A1(n1032), .A2(\registers[25][27] ), .B1(n1029), .B2(
        \registers[24][27] ), .ZN(n2292) );
  AOI22_X1 U2290 ( .A1(n1032), .A2(\registers[25][28] ), .B1(n1029), .B2(
        \registers[24][28] ), .ZN(n2275) );
  AOI22_X1 U2291 ( .A1(n1032), .A2(\registers[25][29] ), .B1(n1029), .B2(
        \registers[24][29] ), .ZN(n2258) );
  AOI22_X1 U2292 ( .A1(n1032), .A2(\registers[25][30] ), .B1(n1029), .B2(
        \registers[24][30] ), .ZN(n2241) );
  AOI22_X1 U2293 ( .A1(n1032), .A2(\registers[25][31] ), .B1(n1029), .B2(
        \registers[24][31] ), .ZN(n2203) );
  AOI22_X1 U2294 ( .A1(n3304), .A2(\registers[25][0] ), .B1(n3301), .B2(
        \registers[24][0] ), .ZN(n2167) );
  AOI22_X1 U2295 ( .A1(n3304), .A2(\registers[25][1] ), .B1(n3301), .B2(
        \registers[24][1] ), .ZN(n2143) );
  AOI22_X1 U2296 ( .A1(n3304), .A2(\registers[25][2] ), .B1(n3301), .B2(
        \registers[24][2] ), .ZN(n2126) );
  AOI22_X1 U2297 ( .A1(n3304), .A2(\registers[25][3] ), .B1(n3301), .B2(
        \registers[24][3] ), .ZN(n2109) );
  AOI22_X1 U2298 ( .A1(n3304), .A2(\registers[25][4] ), .B1(n3301), .B2(
        \registers[24][4] ), .ZN(n2092) );
  AOI22_X1 U2299 ( .A1(n3304), .A2(\registers[25][5] ), .B1(n3301), .B2(
        \registers[24][5] ), .ZN(n2075) );
  AOI22_X1 U2300 ( .A1(n3304), .A2(\registers[25][6] ), .B1(n3301), .B2(
        \registers[24][6] ), .ZN(n2058) );
  AOI22_X1 U2301 ( .A1(n3304), .A2(\registers[25][7] ), .B1(n3301), .B2(
        \registers[24][7] ), .ZN(n2041) );
  AOI22_X1 U2302 ( .A1(n3304), .A2(\registers[25][8] ), .B1(n3301), .B2(
        \registers[24][8] ), .ZN(n2024) );
  AOI22_X1 U2303 ( .A1(n3304), .A2(\registers[25][9] ), .B1(n3301), .B2(
        \registers[24][9] ), .ZN(n2007) );
  AOI22_X1 U2304 ( .A1(n3304), .A2(\registers[25][10] ), .B1(n3301), .B2(
        \registers[24][10] ), .ZN(n1990) );
  AOI22_X1 U2305 ( .A1(n3305), .A2(\registers[25][11] ), .B1(n3302), .B2(
        \registers[24][11] ), .ZN(n1973) );
  AOI22_X1 U2306 ( .A1(n3305), .A2(\registers[25][12] ), .B1(n3302), .B2(
        \registers[24][12] ), .ZN(n1956) );
  AOI22_X1 U2307 ( .A1(n3305), .A2(\registers[25][13] ), .B1(n3302), .B2(
        \registers[24][13] ), .ZN(n1939) );
  AOI22_X1 U2308 ( .A1(n3305), .A2(\registers[25][14] ), .B1(n3302), .B2(
        \registers[24][14] ), .ZN(n1922) );
  AOI22_X1 U2309 ( .A1(n3305), .A2(\registers[25][15] ), .B1(n3302), .B2(
        \registers[24][15] ), .ZN(n1905) );
  AOI22_X1 U2310 ( .A1(n3305), .A2(\registers[25][16] ), .B1(n3302), .B2(
        \registers[24][16] ), .ZN(n1888) );
  AOI22_X1 U2311 ( .A1(n3305), .A2(\registers[25][17] ), .B1(n3302), .B2(
        \registers[24][17] ), .ZN(n1871) );
  AOI22_X1 U2312 ( .A1(n3305), .A2(\registers[25][18] ), .B1(n3302), .B2(
        \registers[24][18] ), .ZN(n1854) );
  AOI22_X1 U2313 ( .A1(n3305), .A2(\registers[25][19] ), .B1(n3302), .B2(
        \registers[24][19] ), .ZN(n1837) );
  AOI22_X1 U2314 ( .A1(n3305), .A2(\registers[25][20] ), .B1(n3302), .B2(
        \registers[24][20] ), .ZN(n1820) );
  AOI22_X1 U2315 ( .A1(n3305), .A2(\registers[25][21] ), .B1(n3302), .B2(
        \registers[24][21] ), .ZN(n1803) );
  AOI22_X1 U2316 ( .A1(n1030), .A2(\registers[25][0] ), .B1(n1027), .B2(
        \registers[24][0] ), .ZN(n2758) );
  AOI22_X1 U2317 ( .A1(n1030), .A2(\registers[25][1] ), .B1(n1027), .B2(
        \registers[24][1] ), .ZN(n2734) );
  AOI22_X1 U2318 ( .A1(n1030), .A2(\registers[25][2] ), .B1(n1027), .B2(
        \registers[24][2] ), .ZN(n2717) );
  AOI22_X1 U2319 ( .A1(n1030), .A2(\registers[25][3] ), .B1(n1027), .B2(
        \registers[24][3] ), .ZN(n2700) );
  AOI22_X1 U2320 ( .A1(n1030), .A2(\registers[25][4] ), .B1(n1027), .B2(
        \registers[24][4] ), .ZN(n2683) );
  AOI22_X1 U2321 ( .A1(n1030), .A2(\registers[25][5] ), .B1(n1027), .B2(
        \registers[24][5] ), .ZN(n2666) );
  AOI22_X1 U2322 ( .A1(n1030), .A2(\registers[25][6] ), .B1(n1027), .B2(
        \registers[24][6] ), .ZN(n2649) );
  AOI22_X1 U2323 ( .A1(n1030), .A2(\registers[25][7] ), .B1(n1027), .B2(
        \registers[24][7] ), .ZN(n2632) );
  AOI22_X1 U2324 ( .A1(n1030), .A2(\registers[25][8] ), .B1(n1027), .B2(
        \registers[24][8] ), .ZN(n2615) );
  AOI22_X1 U2325 ( .A1(n1030), .A2(\registers[25][9] ), .B1(n1027), .B2(
        \registers[24][9] ), .ZN(n2598) );
  AOI22_X1 U2326 ( .A1(n1030), .A2(\registers[25][10] ), .B1(n1027), .B2(
        \registers[24][10] ), .ZN(n2581) );
  AOI22_X1 U2327 ( .A1(n1031), .A2(\registers[25][11] ), .B1(n1028), .B2(
        \registers[24][11] ), .ZN(n2564) );
  AOI22_X1 U2328 ( .A1(n1031), .A2(\registers[25][12] ), .B1(n1028), .B2(
        \registers[24][12] ), .ZN(n2547) );
  AOI22_X1 U2329 ( .A1(n1031), .A2(\registers[25][13] ), .B1(n1028), .B2(
        \registers[24][13] ), .ZN(n2530) );
  AOI22_X1 U2330 ( .A1(n1031), .A2(\registers[25][14] ), .B1(n1028), .B2(
        \registers[24][14] ), .ZN(n2513) );
  AOI22_X1 U2331 ( .A1(n1031), .A2(\registers[25][15] ), .B1(n1028), .B2(
        \registers[24][15] ), .ZN(n2496) );
  AOI22_X1 U2332 ( .A1(n1031), .A2(\registers[25][16] ), .B1(n1028), .B2(
        \registers[24][16] ), .ZN(n2479) );
  AOI22_X1 U2333 ( .A1(n1031), .A2(\registers[25][17] ), .B1(n1028), .B2(
        \registers[24][17] ), .ZN(n2462) );
  AOI22_X1 U2334 ( .A1(n1031), .A2(\registers[25][18] ), .B1(n1028), .B2(
        \registers[24][18] ), .ZN(n2445) );
  AOI22_X1 U2335 ( .A1(n1031), .A2(\registers[25][19] ), .B1(n1028), .B2(
        \registers[24][19] ), .ZN(n2428) );
  AOI22_X1 U2336 ( .A1(n1031), .A2(\registers[25][20] ), .B1(n1028), .B2(
        \registers[24][20] ), .ZN(n2411) );
  AOI22_X1 U2337 ( .A1(n1031), .A2(\registers[25][21] ), .B1(n1028), .B2(
        \registers[24][21] ), .ZN(n2394) );
  AOI22_X1 U2338 ( .A1(n3294), .A2(\registers[29][22] ), .B1(n3291), .B2(
        \registers[28][22] ), .ZN(n1787) );
  AOI22_X1 U2339 ( .A1(n3294), .A2(\registers[29][23] ), .B1(n3291), .B2(
        \registers[28][23] ), .ZN(n1770) );
  AOI22_X1 U2340 ( .A1(n3294), .A2(\registers[29][24] ), .B1(n3291), .B2(
        \registers[28][24] ), .ZN(n1753) );
  AOI22_X1 U2341 ( .A1(n3294), .A2(\registers[29][25] ), .B1(n3291), .B2(
        \registers[28][25] ), .ZN(n1736) );
  AOI22_X1 U2342 ( .A1(n3294), .A2(\registers[29][26] ), .B1(n3291), .B2(
        \registers[28][26] ), .ZN(n1719) );
  AOI22_X1 U2343 ( .A1(n3294), .A2(\registers[29][27] ), .B1(n3291), .B2(
        \registers[28][27] ), .ZN(n1702) );
  AOI22_X1 U2344 ( .A1(n3294), .A2(\registers[29][28] ), .B1(n3291), .B2(
        \registers[28][28] ), .ZN(n1685) );
  AOI22_X1 U2345 ( .A1(n3294), .A2(\registers[29][29] ), .B1(n3291), .B2(
        \registers[28][29] ), .ZN(n1668) );
  AOI22_X1 U2346 ( .A1(n3294), .A2(\registers[29][30] ), .B1(n3291), .B2(
        \registers[28][30] ), .ZN(n1651) );
  AOI22_X1 U2347 ( .A1(n3294), .A2(\registers[29][31] ), .B1(n3291), .B2(
        \registers[28][31] ), .ZN(n1617) );
  AOI22_X1 U2348 ( .A1(n1020), .A2(\registers[29][22] ), .B1(n1017), .B2(
        \registers[28][22] ), .ZN(n2378) );
  AOI22_X1 U2349 ( .A1(n1020), .A2(\registers[29][23] ), .B1(n1017), .B2(
        \registers[28][23] ), .ZN(n2361) );
  AOI22_X1 U2350 ( .A1(n1020), .A2(\registers[29][24] ), .B1(n1017), .B2(
        \registers[28][24] ), .ZN(n2344) );
  AOI22_X1 U2351 ( .A1(n1020), .A2(\registers[29][25] ), .B1(n1017), .B2(
        \registers[28][25] ), .ZN(n2327) );
  AOI22_X1 U2352 ( .A1(n1020), .A2(\registers[29][26] ), .B1(n1017), .B2(
        \registers[28][26] ), .ZN(n2310) );
  AOI22_X1 U2353 ( .A1(n1020), .A2(\registers[29][27] ), .B1(n1017), .B2(
        \registers[28][27] ), .ZN(n2293) );
  AOI22_X1 U2354 ( .A1(n1020), .A2(\registers[29][28] ), .B1(n1017), .B2(
        \registers[28][28] ), .ZN(n2276) );
  AOI22_X1 U2355 ( .A1(n1020), .A2(\registers[29][29] ), .B1(n1017), .B2(
        \registers[28][29] ), .ZN(n2259) );
  AOI22_X1 U2356 ( .A1(n1020), .A2(\registers[29][30] ), .B1(n1017), .B2(
        \registers[28][30] ), .ZN(n2242) );
  AOI22_X1 U2357 ( .A1(n1020), .A2(\registers[29][31] ), .B1(n1017), .B2(
        \registers[28][31] ), .ZN(n2208) );
  AOI22_X1 U2358 ( .A1(n3292), .A2(\registers[29][0] ), .B1(n3289), .B2(
        \registers[28][0] ), .ZN(n2170) );
  AOI22_X1 U2359 ( .A1(n3292), .A2(\registers[29][1] ), .B1(n3289), .B2(
        \registers[28][1] ), .ZN(n2144) );
  AOI22_X1 U2360 ( .A1(n3292), .A2(\registers[29][2] ), .B1(n3289), .B2(
        \registers[28][2] ), .ZN(n2127) );
  AOI22_X1 U2361 ( .A1(n3292), .A2(\registers[29][3] ), .B1(n3289), .B2(
        \registers[28][3] ), .ZN(n2110) );
  AOI22_X1 U2362 ( .A1(n3292), .A2(\registers[29][4] ), .B1(n3289), .B2(
        \registers[28][4] ), .ZN(n2093) );
  AOI22_X1 U2363 ( .A1(n3292), .A2(\registers[29][5] ), .B1(n3289), .B2(
        \registers[28][5] ), .ZN(n2076) );
  AOI22_X1 U2364 ( .A1(n3292), .A2(\registers[29][6] ), .B1(n3289), .B2(
        \registers[28][6] ), .ZN(n2059) );
  AOI22_X1 U2365 ( .A1(n3292), .A2(\registers[29][7] ), .B1(n3289), .B2(
        \registers[28][7] ), .ZN(n2042) );
  AOI22_X1 U2366 ( .A1(n3292), .A2(\registers[29][8] ), .B1(n3289), .B2(
        \registers[28][8] ), .ZN(n2025) );
  AOI22_X1 U2367 ( .A1(n3292), .A2(\registers[29][9] ), .B1(n3289), .B2(
        \registers[28][9] ), .ZN(n2008) );
  AOI22_X1 U2368 ( .A1(n3292), .A2(\registers[29][10] ), .B1(n3289), .B2(
        \registers[28][10] ), .ZN(n1991) );
  AOI22_X1 U2369 ( .A1(n3293), .A2(\registers[29][11] ), .B1(n3290), .B2(
        \registers[28][11] ), .ZN(n1974) );
  AOI22_X1 U2370 ( .A1(n3293), .A2(\registers[29][12] ), .B1(n3290), .B2(
        \registers[28][12] ), .ZN(n1957) );
  AOI22_X1 U2371 ( .A1(n3293), .A2(\registers[29][13] ), .B1(n3290), .B2(
        \registers[28][13] ), .ZN(n1940) );
  AOI22_X1 U2372 ( .A1(n3293), .A2(\registers[29][14] ), .B1(n3290), .B2(
        \registers[28][14] ), .ZN(n1923) );
  AOI22_X1 U2373 ( .A1(n3293), .A2(\registers[29][15] ), .B1(n3290), .B2(
        \registers[28][15] ), .ZN(n1906) );
  AOI22_X1 U2374 ( .A1(n3293), .A2(\registers[29][16] ), .B1(n3290), .B2(
        \registers[28][16] ), .ZN(n1889) );
  AOI22_X1 U2375 ( .A1(n3293), .A2(\registers[29][17] ), .B1(n3290), .B2(
        \registers[28][17] ), .ZN(n1872) );
  AOI22_X1 U2376 ( .A1(n3293), .A2(\registers[29][18] ), .B1(n3290), .B2(
        \registers[28][18] ), .ZN(n1855) );
  AOI22_X1 U2377 ( .A1(n3293), .A2(\registers[29][19] ), .B1(n3290), .B2(
        \registers[28][19] ), .ZN(n1838) );
  AOI22_X1 U2378 ( .A1(n3293), .A2(\registers[29][20] ), .B1(n3290), .B2(
        \registers[28][20] ), .ZN(n1821) );
  AOI22_X1 U2379 ( .A1(n3293), .A2(\registers[29][21] ), .B1(n3290), .B2(
        \registers[28][21] ), .ZN(n1804) );
  AOI22_X1 U2380 ( .A1(n1018), .A2(\registers[29][0] ), .B1(n1015), .B2(
        \registers[28][0] ), .ZN(n2761) );
  AOI22_X1 U2381 ( .A1(n1018), .A2(\registers[29][1] ), .B1(n1015), .B2(
        \registers[28][1] ), .ZN(n2735) );
  AOI22_X1 U2382 ( .A1(n1018), .A2(\registers[29][2] ), .B1(n1015), .B2(
        \registers[28][2] ), .ZN(n2718) );
  AOI22_X1 U2383 ( .A1(n1018), .A2(\registers[29][3] ), .B1(n1015), .B2(
        \registers[28][3] ), .ZN(n2701) );
  AOI22_X1 U2384 ( .A1(n1018), .A2(\registers[29][4] ), .B1(n1015), .B2(
        \registers[28][4] ), .ZN(n2684) );
  AOI22_X1 U2385 ( .A1(n1018), .A2(\registers[29][5] ), .B1(n1015), .B2(
        \registers[28][5] ), .ZN(n2667) );
  AOI22_X1 U2386 ( .A1(n1018), .A2(\registers[29][6] ), .B1(n1015), .B2(
        \registers[28][6] ), .ZN(n2650) );
  AOI22_X1 U2387 ( .A1(n1018), .A2(\registers[29][7] ), .B1(n1015), .B2(
        \registers[28][7] ), .ZN(n2633) );
  AOI22_X1 U2388 ( .A1(n1018), .A2(\registers[29][8] ), .B1(n1015), .B2(
        \registers[28][8] ), .ZN(n2616) );
  AOI22_X1 U2389 ( .A1(n1018), .A2(\registers[29][9] ), .B1(n1015), .B2(
        \registers[28][9] ), .ZN(n2599) );
  AOI22_X1 U2390 ( .A1(n1018), .A2(\registers[29][10] ), .B1(n1015), .B2(
        \registers[28][10] ), .ZN(n2582) );
  AOI22_X1 U2391 ( .A1(n1019), .A2(\registers[29][11] ), .B1(n1016), .B2(
        \registers[28][11] ), .ZN(n2565) );
  AOI22_X1 U2392 ( .A1(n1019), .A2(\registers[29][12] ), .B1(n1016), .B2(
        \registers[28][12] ), .ZN(n2548) );
  AOI22_X1 U2393 ( .A1(n1019), .A2(\registers[29][13] ), .B1(n1016), .B2(
        \registers[28][13] ), .ZN(n2531) );
  AOI22_X1 U2394 ( .A1(n1019), .A2(\registers[29][14] ), .B1(n1016), .B2(
        \registers[28][14] ), .ZN(n2514) );
  AOI22_X1 U2395 ( .A1(n1019), .A2(\registers[29][15] ), .B1(n1016), .B2(
        \registers[28][15] ), .ZN(n2497) );
  AOI22_X1 U2396 ( .A1(n1019), .A2(\registers[29][16] ), .B1(n1016), .B2(
        \registers[28][16] ), .ZN(n2480) );
  AOI22_X1 U2397 ( .A1(n1019), .A2(\registers[29][17] ), .B1(n1016), .B2(
        \registers[28][17] ), .ZN(n2463) );
  AOI22_X1 U2398 ( .A1(n1019), .A2(\registers[29][18] ), .B1(n1016), .B2(
        \registers[28][18] ), .ZN(n2446) );
  AOI22_X1 U2399 ( .A1(n1019), .A2(\registers[29][19] ), .B1(n1016), .B2(
        \registers[28][19] ), .ZN(n2429) );
  AOI22_X1 U2400 ( .A1(n1019), .A2(\registers[29][20] ), .B1(n1016), .B2(
        \registers[28][20] ), .ZN(n2412) );
  AOI22_X1 U2401 ( .A1(n1019), .A2(\registers[29][21] ), .B1(n1016), .B2(
        \registers[28][21] ), .ZN(n2395) );
  OAI22_X1 U2402 ( .A1(n3584), .A2(n4201), .B1(n3581), .B2(n982), .ZN(n2784)
         );
  OAI22_X1 U2403 ( .A1(n3582), .A2(n790), .B1(n3580), .B2(n981), .ZN(n2785) );
  OAI22_X1 U2404 ( .A1(n3583), .A2(n4199), .B1(n3579), .B2(n980), .ZN(n2786)
         );
  OAI22_X1 U2405 ( .A1(n3582), .A2(n4198), .B1(n3579), .B2(n979), .ZN(n2787)
         );
  OAI22_X1 U2406 ( .A1(n3582), .A2(n4197), .B1(n3580), .B2(n978), .ZN(n2788)
         );
  OAI22_X1 U2407 ( .A1(n3582), .A2(n4196), .B1(n3581), .B2(n977), .ZN(n2789)
         );
  OAI22_X1 U2408 ( .A1(n3582), .A2(n4195), .B1(n3579), .B2(n976), .ZN(n2790)
         );
  OAI22_X1 U2409 ( .A1(n3584), .A2(n4194), .B1(n3580), .B2(n975), .ZN(n2791)
         );
  OAI22_X1 U2410 ( .A1(n3583), .A2(n4193), .B1(n3581), .B2(n974), .ZN(n2792)
         );
  OAI22_X1 U2411 ( .A1(n3584), .A2(n677), .B1(n3579), .B2(n973), .ZN(n2793) );
  OAI22_X1 U2412 ( .A1(n3582), .A2(n687), .B1(n3579), .B2(n972), .ZN(n2794) );
  OAI22_X1 U2413 ( .A1(n3583), .A2(n257), .B1(n3580), .B2(n971), .ZN(n2795) );
  OAI22_X1 U2414 ( .A1(n3584), .A2(n4189), .B1(n3581), .B2(n970), .ZN(n2796)
         );
  OAI22_X1 U2415 ( .A1(n3584), .A2(n285), .B1(n3581), .B2(n969), .ZN(n2797) );
  OAI22_X1 U2416 ( .A1(n3582), .A2(n4187), .B1(n3579), .B2(n968), .ZN(n2798)
         );
  OAI22_X1 U2417 ( .A1(n3582), .A2(n282), .B1(n3579), .B2(n967), .ZN(n2799) );
  OAI22_X1 U2418 ( .A1(n3583), .A2(n684), .B1(n3580), .B2(n966), .ZN(n2800) );
  OAI22_X1 U2419 ( .A1(n3582), .A2(n271), .B1(n3581), .B2(n965), .ZN(n2801) );
  OAI22_X1 U2420 ( .A1(n3582), .A2(n683), .B1(n3580), .B2(n964), .ZN(n2802) );
  OAI22_X1 U2421 ( .A1(n3584), .A2(n376), .B1(n3579), .B2(n963), .ZN(n2803) );
  OAI22_X1 U2422 ( .A1(n3582), .A2(n681), .B1(n3580), .B2(n962), .ZN(n2804) );
  OAI22_X1 U2423 ( .A1(n3584), .A2(n713), .B1(n3581), .B2(n961), .ZN(n2805) );
  OAI22_X1 U2424 ( .A1(n3582), .A2(n4211), .B1(n3581), .B2(n992), .ZN(n2774)
         );
  OAI22_X1 U2425 ( .A1(n3582), .A2(n4210), .B1(n3580), .B2(n991), .ZN(n2775)
         );
  OAI22_X1 U2426 ( .A1(n3583), .A2(n4209), .B1(n3581), .B2(n990), .ZN(n2776)
         );
  OAI22_X1 U2427 ( .A1(n3583), .A2(n691), .B1(n3581), .B2(n989), .ZN(n2777) );
  OAI22_X1 U2428 ( .A1(n3582), .A2(n356), .B1(n3579), .B2(n988), .ZN(n2778) );
  OAI22_X1 U2429 ( .A1(n3584), .A2(n4206), .B1(n3580), .B2(n987), .ZN(n2779)
         );
  OAI22_X1 U2430 ( .A1(n3582), .A2(n714), .B1(n3580), .B2(n986), .ZN(n2780) );
  OAI22_X1 U2431 ( .A1(n3584), .A2(n4204), .B1(n3579), .B2(n985), .ZN(n2781)
         );
  OAI22_X1 U2432 ( .A1(n3582), .A2(n689), .B1(n3579), .B2(n984), .ZN(n2782) );
  OAI22_X1 U2433 ( .A1(n3583), .A2(n370), .B1(n3580), .B2(n983), .ZN(n2783) );
  AND2_X1 U2434 ( .A1(ADD_RD2[0]), .A2(n2171), .ZN(n2169) );
  AND2_X1 U2435 ( .A1(ADD_RD1[0]), .A2(n2762), .ZN(n2760) );
  NAND4_X1 U2436 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(N343)
         );
  AOI221_X1 U2437 ( .B1(n1252), .B2(\registers[9][22] ), .C1(n1143), .C2(
        \registers[8][22] ), .A(n1792), .ZN(n1776) );
  AOI221_X1 U2438 ( .B1(n1353), .B2(\registers[13][22] ), .C1(n1349), .C2(
        \registers[12][22] ), .A(n1791), .ZN(n1777) );
  AOI211_X1 U2439 ( .C1(n3288), .C2(\registers[1][22] ), .A(n1788), .B(n1789), 
        .ZN(n1778) );
  NAND4_X1 U2440 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(N344)
         );
  AOI221_X1 U2441 ( .B1(n1252), .B2(\registers[9][23] ), .C1(n1143), .C2(
        \registers[8][23] ), .A(n1775), .ZN(n1759) );
  AOI221_X1 U2442 ( .B1(n1353), .B2(\registers[13][23] ), .C1(n1349), .C2(
        \registers[12][23] ), .A(n1774), .ZN(n1760) );
  AOI211_X1 U2443 ( .C1(n3288), .C2(\registers[1][23] ), .A(n1771), .B(n1772), 
        .ZN(n1761) );
  NAND4_X1 U2444 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(N345)
         );
  AOI221_X1 U2445 ( .B1(n1252), .B2(\registers[9][24] ), .C1(n1143), .C2(
        \registers[8][24] ), .A(n1758), .ZN(n1742) );
  AOI221_X1 U2446 ( .B1(n1353), .B2(\registers[13][24] ), .C1(n1349), .C2(
        \registers[12][24] ), .A(n1757), .ZN(n1743) );
  AOI211_X1 U2447 ( .C1(n3288), .C2(\registers[1][24] ), .A(n1754), .B(n1755), 
        .ZN(n1744) );
  NAND4_X1 U2448 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(N346)
         );
  AOI221_X1 U2449 ( .B1(n1252), .B2(\registers[9][25] ), .C1(n1143), .C2(
        \registers[8][25] ), .A(n1741), .ZN(n1725) );
  AOI221_X1 U2450 ( .B1(n1353), .B2(\registers[13][25] ), .C1(n1349), .C2(
        \registers[12][25] ), .A(n1740), .ZN(n1726) );
  AOI211_X1 U2451 ( .C1(n3288), .C2(\registers[1][25] ), .A(n1737), .B(n1738), 
        .ZN(n1727) );
  NAND4_X1 U2452 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(N347)
         );
  AOI221_X1 U2453 ( .B1(n1252), .B2(\registers[9][26] ), .C1(n1143), .C2(
        \registers[8][26] ), .A(n1724), .ZN(n1708) );
  AOI221_X1 U2454 ( .B1(n1353), .B2(\registers[13][26] ), .C1(n1349), .C2(
        \registers[12][26] ), .A(n1723), .ZN(n1709) );
  AOI211_X1 U2455 ( .C1(n3288), .C2(\registers[1][26] ), .A(n1720), .B(n1721), 
        .ZN(n1710) );
  NAND4_X1 U2456 ( .A1(n1691), .A2(n1692), .A3(n1693), .A4(n1694), .ZN(N348)
         );
  AOI221_X1 U2457 ( .B1(n1252), .B2(\registers[9][27] ), .C1(n1143), .C2(
        \registers[8][27] ), .A(n1707), .ZN(n1691) );
  AOI221_X1 U2458 ( .B1(n1353), .B2(\registers[13][27] ), .C1(n1349), .C2(
        \registers[12][27] ), .A(n1706), .ZN(n1692) );
  AOI211_X1 U2459 ( .C1(n3288), .C2(\registers[1][27] ), .A(n1703), .B(n1704), 
        .ZN(n1693) );
  NAND4_X1 U2460 ( .A1(n1674), .A2(n1675), .A3(n1676), .A4(n1677), .ZN(N349)
         );
  AOI221_X1 U2461 ( .B1(n1252), .B2(\registers[9][28] ), .C1(n1143), .C2(
        \registers[8][28] ), .A(n1690), .ZN(n1674) );
  AOI221_X1 U2462 ( .B1(n1353), .B2(\registers[13][28] ), .C1(n1349), .C2(
        \registers[12][28] ), .A(n1689), .ZN(n1675) );
  AOI211_X1 U2463 ( .C1(n3288), .C2(\registers[1][28] ), .A(n1686), .B(n1687), 
        .ZN(n1676) );
  NAND4_X1 U2464 ( .A1(n1657), .A2(n1658), .A3(n1659), .A4(n1660), .ZN(N350)
         );
  AOI221_X1 U2465 ( .B1(n1252), .B2(\registers[9][29] ), .C1(n1143), .C2(
        \registers[8][29] ), .A(n1673), .ZN(n1657) );
  AOI221_X1 U2466 ( .B1(n1353), .B2(\registers[13][29] ), .C1(n1349), .C2(
        \registers[12][29] ), .A(n1672), .ZN(n1658) );
  AOI211_X1 U2467 ( .C1(n3288), .C2(\registers[1][29] ), .A(n1669), .B(n1670), 
        .ZN(n1659) );
  NAND4_X1 U2468 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .ZN(N351)
         );
  AOI221_X1 U2469 ( .B1(n1252), .B2(\registers[9][30] ), .C1(n1143), .C2(
        \registers[8][30] ), .A(n1656), .ZN(n1640) );
  AOI221_X1 U2470 ( .B1(n1353), .B2(\registers[13][30] ), .C1(n1349), .C2(
        \registers[12][30] ), .A(n1655), .ZN(n1641) );
  AOI211_X1 U2471 ( .C1(n3288), .C2(\registers[1][30] ), .A(n1652), .B(n1653), 
        .ZN(n1642) );
  NAND4_X1 U2472 ( .A1(n1592), .A2(n1593), .A3(n1594), .A4(n1595), .ZN(N352)
         );
  AOI221_X1 U2473 ( .B1(n1252), .B2(\registers[9][31] ), .C1(n1143), .C2(
        \registers[8][31] ), .A(n1637), .ZN(n1592) );
  AOI221_X1 U2474 ( .B1(n1353), .B2(\registers[13][31] ), .C1(n1349), .C2(
        \registers[12][31] ), .A(n1632), .ZN(n1593) );
  AOI211_X1 U2475 ( .C1(n3288), .C2(\registers[1][31] ), .A(n1621), .B(n1622), 
        .ZN(n1594) );
  NAND4_X1 U2476 ( .A1(n2367), .A2(n2368), .A3(n2369), .A4(n2370), .ZN(N208)
         );
  AOI221_X1 U2477 ( .B1(n917), .B2(\registers[9][22] ), .C1(n914), .C2(
        \registers[8][22] ), .A(n2383), .ZN(n2367) );
  AOI221_X1 U2478 ( .B1(n993), .B2(\registers[13][22] ), .C1(n926), .C2(
        \registers[12][22] ), .A(n2382), .ZN(n2368) );
  AOI211_X1 U2479 ( .C1(n1014), .C2(\registers[1][22] ), .A(n2379), .B(n2380), 
        .ZN(n2369) );
  NAND4_X1 U2480 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(N209)
         );
  AOI221_X1 U2481 ( .B1(n917), .B2(\registers[9][23] ), .C1(n914), .C2(
        \registers[8][23] ), .A(n2366), .ZN(n2350) );
  AOI221_X1 U2482 ( .B1(n993), .B2(\registers[13][23] ), .C1(n926), .C2(
        \registers[12][23] ), .A(n2365), .ZN(n2351) );
  AOI211_X1 U2483 ( .C1(n1014), .C2(\registers[1][23] ), .A(n2362), .B(n2363), 
        .ZN(n2352) );
  NAND4_X1 U2484 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(N210)
         );
  AOI221_X1 U2485 ( .B1(n917), .B2(\registers[9][24] ), .C1(n914), .C2(
        \registers[8][24] ), .A(n2349), .ZN(n2333) );
  AOI221_X1 U2486 ( .B1(n993), .B2(\registers[13][24] ), .C1(n926), .C2(
        \registers[12][24] ), .A(n2348), .ZN(n2334) );
  AOI211_X1 U2487 ( .C1(n1014), .C2(\registers[1][24] ), .A(n2345), .B(n2346), 
        .ZN(n2335) );
  NAND4_X1 U2488 ( .A1(n2316), .A2(n2317), .A3(n2318), .A4(n2319), .ZN(N211)
         );
  AOI221_X1 U2489 ( .B1(n917), .B2(\registers[9][25] ), .C1(n914), .C2(
        \registers[8][25] ), .A(n2332), .ZN(n2316) );
  AOI221_X1 U2490 ( .B1(n993), .B2(\registers[13][25] ), .C1(n926), .C2(
        \registers[12][25] ), .A(n2331), .ZN(n2317) );
  AOI211_X1 U2491 ( .C1(n1014), .C2(\registers[1][25] ), .A(n2328), .B(n2329), 
        .ZN(n2318) );
  NAND4_X1 U2492 ( .A1(n2299), .A2(n2300), .A3(n2301), .A4(n2302), .ZN(N212)
         );
  AOI221_X1 U2493 ( .B1(n917), .B2(\registers[9][26] ), .C1(n914), .C2(
        \registers[8][26] ), .A(n2315), .ZN(n2299) );
  AOI221_X1 U2494 ( .B1(n993), .B2(\registers[13][26] ), .C1(n926), .C2(
        \registers[12][26] ), .A(n2314), .ZN(n2300) );
  AOI211_X1 U2495 ( .C1(n1014), .C2(\registers[1][26] ), .A(n2311), .B(n2312), 
        .ZN(n2301) );
  NAND4_X1 U2496 ( .A1(n2282), .A2(n2283), .A3(n2284), .A4(n2285), .ZN(N213)
         );
  AOI221_X1 U2497 ( .B1(n917), .B2(\registers[9][27] ), .C1(n914), .C2(
        \registers[8][27] ), .A(n2298), .ZN(n2282) );
  AOI221_X1 U2498 ( .B1(n993), .B2(\registers[13][27] ), .C1(n926), .C2(
        \registers[12][27] ), .A(n2297), .ZN(n2283) );
  AOI211_X1 U2499 ( .C1(n1014), .C2(\registers[1][27] ), .A(n2294), .B(n2295), 
        .ZN(n2284) );
  NAND4_X1 U2500 ( .A1(n2265), .A2(n2266), .A3(n2267), .A4(n2268), .ZN(N214)
         );
  AOI221_X1 U2501 ( .B1(n917), .B2(\registers[9][28] ), .C1(n914), .C2(
        \registers[8][28] ), .A(n2281), .ZN(n2265) );
  AOI221_X1 U2502 ( .B1(n993), .B2(\registers[13][28] ), .C1(n926), .C2(
        \registers[12][28] ), .A(n2280), .ZN(n2266) );
  AOI211_X1 U2503 ( .C1(n1014), .C2(\registers[1][28] ), .A(n2277), .B(n2278), 
        .ZN(n2267) );
  NAND4_X1 U2504 ( .A1(n2248), .A2(n2249), .A3(n2250), .A4(n2251), .ZN(N215)
         );
  AOI221_X1 U2505 ( .B1(n917), .B2(\registers[9][29] ), .C1(n914), .C2(
        \registers[8][29] ), .A(n2264), .ZN(n2248) );
  AOI221_X1 U2506 ( .B1(n993), .B2(\registers[13][29] ), .C1(n926), .C2(
        \registers[12][29] ), .A(n2263), .ZN(n2249) );
  AOI211_X1 U2507 ( .C1(n1014), .C2(\registers[1][29] ), .A(n2260), .B(n2261), 
        .ZN(n2250) );
  NAND4_X1 U2508 ( .A1(n2231), .A2(n2232), .A3(n2233), .A4(n2234), .ZN(N216)
         );
  AOI221_X1 U2509 ( .B1(n917), .B2(\registers[9][30] ), .C1(n914), .C2(
        \registers[8][30] ), .A(n2247), .ZN(n2231) );
  AOI221_X1 U2510 ( .B1(n993), .B2(\registers[13][30] ), .C1(n926), .C2(
        \registers[12][30] ), .A(n2246), .ZN(n2232) );
  AOI211_X1 U2511 ( .C1(n1014), .C2(\registers[1][30] ), .A(n2243), .B(n2244), 
        .ZN(n2233) );
  NAND4_X1 U2512 ( .A1(n2183), .A2(n2184), .A3(n2185), .A4(n2186), .ZN(N217)
         );
  AOI221_X1 U2513 ( .B1(n917), .B2(\registers[9][31] ), .C1(n914), .C2(
        \registers[8][31] ), .A(n2228), .ZN(n2183) );
  AOI221_X1 U2514 ( .B1(n993), .B2(\registers[13][31] ), .C1(n926), .C2(
        \registers[12][31] ), .A(n2223), .ZN(n2184) );
  AOI211_X1 U2515 ( .C1(n1014), .C2(\registers[1][31] ), .A(n2212), .B(n2213), 
        .ZN(n2185) );
  NAND4_X1 U2516 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .ZN(N321)
         );
  AOI221_X1 U2517 ( .B1(n1248), .B2(\registers[9][0] ), .C1(n1113), .C2(
        \registers[8][0] ), .A(n2181), .ZN(n2150) );
  AOI221_X1 U2518 ( .B1(n1350), .B2(\registers[13][0] ), .C1(n1285), .C2(
        \registers[12][0] ), .A(n2178), .ZN(n2151) );
  AOI211_X1 U2519 ( .C1(n3286), .C2(\registers[1][0] ), .A(n2172), .B(n2173), 
        .ZN(n2152) );
  NAND4_X1 U2520 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(N322)
         );
  AOI221_X1 U2521 ( .B1(n1248), .B2(\registers[9][1] ), .C1(n1113), .C2(
        \registers[8][1] ), .A(n2149), .ZN(n2133) );
  AOI221_X1 U2522 ( .B1(n1350), .B2(\registers[13][1] ), .C1(n1285), .C2(
        \registers[12][1] ), .A(n2148), .ZN(n2134) );
  AOI211_X1 U2523 ( .C1(n3286), .C2(\registers[1][1] ), .A(n2145), .B(n2146), 
        .ZN(n2135) );
  NAND4_X1 U2524 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(N323)
         );
  AOI221_X1 U2525 ( .B1(n1248), .B2(\registers[9][2] ), .C1(n1113), .C2(
        \registers[8][2] ), .A(n2132), .ZN(n2116) );
  AOI221_X1 U2526 ( .B1(n1350), .B2(\registers[13][2] ), .C1(n1285), .C2(
        \registers[12][2] ), .A(n2131), .ZN(n2117) );
  AOI211_X1 U2527 ( .C1(n3286), .C2(\registers[1][2] ), .A(n2128), .B(n2129), 
        .ZN(n2118) );
  NAND4_X1 U2528 ( .A1(n2099), .A2(n2100), .A3(n2101), .A4(n2102), .ZN(N324)
         );
  AOI221_X1 U2529 ( .B1(n1248), .B2(\registers[9][3] ), .C1(n1113), .C2(
        \registers[8][3] ), .A(n2115), .ZN(n2099) );
  AOI221_X1 U2530 ( .B1(n1350), .B2(\registers[13][3] ), .C1(n1285), .C2(
        \registers[12][3] ), .A(n2114), .ZN(n2100) );
  AOI211_X1 U2531 ( .C1(n3286), .C2(\registers[1][3] ), .A(n2111), .B(n2112), 
        .ZN(n2101) );
  NAND4_X1 U2532 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(N325)
         );
  AOI221_X1 U2533 ( .B1(n1248), .B2(\registers[9][4] ), .C1(n1113), .C2(
        \registers[8][4] ), .A(n2098), .ZN(n2082) );
  AOI221_X1 U2534 ( .B1(n1350), .B2(\registers[13][4] ), .C1(n1285), .C2(
        \registers[12][4] ), .A(n2097), .ZN(n2083) );
  AOI211_X1 U2535 ( .C1(n3286), .C2(\registers[1][4] ), .A(n2094), .B(n2095), 
        .ZN(n2084) );
  NAND4_X1 U2536 ( .A1(n2065), .A2(n2066), .A3(n2067), .A4(n2068), .ZN(N326)
         );
  AOI221_X1 U2537 ( .B1(n1248), .B2(\registers[9][5] ), .C1(n1113), .C2(
        \registers[8][5] ), .A(n2081), .ZN(n2065) );
  AOI221_X1 U2538 ( .B1(n1350), .B2(\registers[13][5] ), .C1(n1285), .C2(
        \registers[12][5] ), .A(n2080), .ZN(n2066) );
  AOI211_X1 U2539 ( .C1(n3286), .C2(\registers[1][5] ), .A(n2077), .B(n2078), 
        .ZN(n2067) );
  NAND4_X1 U2540 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(N327)
         );
  AOI221_X1 U2541 ( .B1(n1248), .B2(\registers[9][6] ), .C1(n1113), .C2(
        \registers[8][6] ), .A(n2064), .ZN(n2048) );
  AOI221_X1 U2542 ( .B1(n1350), .B2(\registers[13][6] ), .C1(n1285), .C2(
        \registers[12][6] ), .A(n2063), .ZN(n2049) );
  AOI211_X1 U2543 ( .C1(n3286), .C2(\registers[1][6] ), .A(n2060), .B(n2061), 
        .ZN(n2050) );
  NAND4_X1 U2544 ( .A1(n2031), .A2(n2032), .A3(n2033), .A4(n2034), .ZN(N328)
         );
  AOI221_X1 U2545 ( .B1(n1248), .B2(\registers[9][7] ), .C1(n1113), .C2(
        \registers[8][7] ), .A(n2047), .ZN(n2031) );
  AOI221_X1 U2546 ( .B1(n1350), .B2(\registers[13][7] ), .C1(n1285), .C2(
        \registers[12][7] ), .A(n2046), .ZN(n2032) );
  AOI211_X1 U2547 ( .C1(n3286), .C2(\registers[1][7] ), .A(n2043), .B(n2044), 
        .ZN(n2033) );
  NAND4_X1 U2548 ( .A1(n2014), .A2(n2015), .A3(n2016), .A4(n2017), .ZN(N329)
         );
  AOI221_X1 U2549 ( .B1(n1248), .B2(\registers[9][8] ), .C1(n1113), .C2(
        \registers[8][8] ), .A(n2030), .ZN(n2014) );
  AOI221_X1 U2550 ( .B1(n1350), .B2(\registers[13][8] ), .C1(n1285), .C2(
        \registers[12][8] ), .A(n2029), .ZN(n2015) );
  AOI211_X1 U2551 ( .C1(n3286), .C2(\registers[1][8] ), .A(n2026), .B(n2027), 
        .ZN(n2016) );
  NAND4_X1 U2552 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(N330)
         );
  AOI221_X1 U2553 ( .B1(n1248), .B2(\registers[9][9] ), .C1(n1113), .C2(
        \registers[8][9] ), .A(n2013), .ZN(n1997) );
  AOI221_X1 U2554 ( .B1(n1350), .B2(\registers[13][9] ), .C1(n1285), .C2(
        \registers[12][9] ), .A(n2012), .ZN(n1998) );
  AOI211_X1 U2555 ( .C1(n3286), .C2(\registers[1][9] ), .A(n2009), .B(n2010), 
        .ZN(n1999) );
  NAND4_X1 U2556 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .ZN(N331)
         );
  AOI221_X1 U2557 ( .B1(n1248), .B2(\registers[9][10] ), .C1(n1113), .C2(
        \registers[8][10] ), .A(n1996), .ZN(n1980) );
  AOI221_X1 U2558 ( .B1(n1350), .B2(\registers[13][10] ), .C1(n1285), .C2(
        \registers[12][10] ), .A(n1995), .ZN(n1981) );
  AOI211_X1 U2559 ( .C1(n3286), .C2(\registers[1][10] ), .A(n1992), .B(n1993), 
        .ZN(n1982) );
  NAND4_X1 U2560 ( .A1(n1963), .A2(n1964), .A3(n1965), .A4(n1966), .ZN(N332)
         );
  AOI221_X1 U2561 ( .B1(n1250), .B2(\registers[9][11] ), .C1(n1141), .C2(
        \registers[8][11] ), .A(n1979), .ZN(n1963) );
  AOI221_X1 U2562 ( .B1(n1351), .B2(\registers[13][11] ), .C1(n1320), .C2(
        \registers[12][11] ), .A(n1978), .ZN(n1964) );
  AOI211_X1 U2563 ( .C1(n3287), .C2(\registers[1][11] ), .A(n1975), .B(n1976), 
        .ZN(n1965) );
  NAND4_X1 U2564 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(N333)
         );
  AOI221_X1 U2565 ( .B1(n1250), .B2(\registers[9][12] ), .C1(n1141), .C2(
        \registers[8][12] ), .A(n1962), .ZN(n1946) );
  AOI221_X1 U2566 ( .B1(n1351), .B2(\registers[13][12] ), .C1(n1320), .C2(
        \registers[12][12] ), .A(n1961), .ZN(n1947) );
  AOI211_X1 U2567 ( .C1(n3287), .C2(\registers[1][12] ), .A(n1958), .B(n1959), 
        .ZN(n1948) );
  NAND4_X1 U2568 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(N334)
         );
  AOI221_X1 U2569 ( .B1(n1250), .B2(\registers[9][13] ), .C1(n1141), .C2(
        \registers[8][13] ), .A(n1945), .ZN(n1929) );
  AOI221_X1 U2570 ( .B1(n1351), .B2(\registers[13][13] ), .C1(n1320), .C2(
        \registers[12][13] ), .A(n1944), .ZN(n1930) );
  AOI211_X1 U2571 ( .C1(n3287), .C2(\registers[1][13] ), .A(n1941), .B(n1942), 
        .ZN(n1931) );
  NAND4_X1 U2572 ( .A1(n1912), .A2(n1913), .A3(n1914), .A4(n1915), .ZN(N335)
         );
  AOI221_X1 U2573 ( .B1(n1250), .B2(\registers[9][14] ), .C1(n1141), .C2(
        \registers[8][14] ), .A(n1928), .ZN(n1912) );
  AOI221_X1 U2574 ( .B1(n1351), .B2(\registers[13][14] ), .C1(n1320), .C2(
        \registers[12][14] ), .A(n1927), .ZN(n1913) );
  AOI211_X1 U2575 ( .C1(n3287), .C2(\registers[1][14] ), .A(n1924), .B(n1925), 
        .ZN(n1914) );
  NAND4_X1 U2576 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(N336)
         );
  AOI221_X1 U2577 ( .B1(n1250), .B2(\registers[9][15] ), .C1(n1141), .C2(
        \registers[8][15] ), .A(n1911), .ZN(n1895) );
  AOI221_X1 U2578 ( .B1(n1351), .B2(\registers[13][15] ), .C1(n1320), .C2(
        \registers[12][15] ), .A(n1910), .ZN(n1896) );
  AOI211_X1 U2579 ( .C1(n3287), .C2(\registers[1][15] ), .A(n1907), .B(n1908), 
        .ZN(n1897) );
  NAND4_X1 U2580 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .ZN(N337)
         );
  AOI221_X1 U2581 ( .B1(n1250), .B2(\registers[9][16] ), .C1(n1141), .C2(
        \registers[8][16] ), .A(n1894), .ZN(n1878) );
  AOI221_X1 U2582 ( .B1(n1351), .B2(\registers[13][16] ), .C1(n1320), .C2(
        \registers[12][16] ), .A(n1893), .ZN(n1879) );
  AOI211_X1 U2583 ( .C1(n3287), .C2(\registers[1][16] ), .A(n1890), .B(n1891), 
        .ZN(n1880) );
  NAND4_X1 U2584 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .ZN(N338)
         );
  AOI221_X1 U2585 ( .B1(n1250), .B2(\registers[9][17] ), .C1(n1141), .C2(
        \registers[8][17] ), .A(n1877), .ZN(n1861) );
  AOI221_X1 U2586 ( .B1(n1351), .B2(\registers[13][17] ), .C1(n1320), .C2(
        \registers[12][17] ), .A(n1876), .ZN(n1862) );
  AOI211_X1 U2587 ( .C1(n3287), .C2(\registers[1][17] ), .A(n1873), .B(n1874), 
        .ZN(n1863) );
  NAND4_X1 U2588 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .ZN(N339)
         );
  AOI221_X1 U2589 ( .B1(n1250), .B2(\registers[9][18] ), .C1(n1141), .C2(
        \registers[8][18] ), .A(n1860), .ZN(n1844) );
  AOI221_X1 U2590 ( .B1(n1351), .B2(\registers[13][18] ), .C1(n1320), .C2(
        \registers[12][18] ), .A(n1859), .ZN(n1845) );
  AOI211_X1 U2591 ( .C1(n3287), .C2(\registers[1][18] ), .A(n1856), .B(n1857), 
        .ZN(n1846) );
  NAND4_X1 U2592 ( .A1(n1827), .A2(n1828), .A3(n1829), .A4(n1830), .ZN(N340)
         );
  AOI221_X1 U2593 ( .B1(n1250), .B2(\registers[9][19] ), .C1(n1141), .C2(
        \registers[8][19] ), .A(n1843), .ZN(n1827) );
  AOI221_X1 U2594 ( .B1(n1351), .B2(\registers[13][19] ), .C1(n1320), .C2(
        \registers[12][19] ), .A(n1842), .ZN(n1828) );
  AOI211_X1 U2595 ( .C1(n3287), .C2(\registers[1][19] ), .A(n1839), .B(n1840), 
        .ZN(n1829) );
  NAND4_X1 U2596 ( .A1(n1810), .A2(n1811), .A3(n1812), .A4(n1813), .ZN(N341)
         );
  AOI221_X1 U2597 ( .B1(n1250), .B2(\registers[9][20] ), .C1(n1141), .C2(
        \registers[8][20] ), .A(n1826), .ZN(n1810) );
  AOI221_X1 U2598 ( .B1(n1351), .B2(\registers[13][20] ), .C1(n1320), .C2(
        \registers[12][20] ), .A(n1825), .ZN(n1811) );
  AOI211_X1 U2599 ( .C1(n3287), .C2(\registers[1][20] ), .A(n1822), .B(n1823), 
        .ZN(n1812) );
  NAND4_X1 U2600 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .ZN(N342)
         );
  AOI221_X1 U2601 ( .B1(n1250), .B2(\registers[9][21] ), .C1(n1141), .C2(
        \registers[8][21] ), .A(n1809), .ZN(n1793) );
  AOI221_X1 U2602 ( .B1(n1351), .B2(\registers[13][21] ), .C1(n1320), .C2(
        \registers[12][21] ), .A(n1808), .ZN(n1794) );
  AOI211_X1 U2603 ( .C1(n3287), .C2(\registers[1][21] ), .A(n1805), .B(n1806), 
        .ZN(n1795) );
  NAND4_X1 U2604 ( .A1(n2741), .A2(n2742), .A3(n2743), .A4(n2744), .ZN(N186)
         );
  AOI221_X1 U2605 ( .B1(n915), .B2(\registers[9][0] ), .C1(n912), .C2(
        \registers[8][0] ), .A(n2772), .ZN(n2741) );
  AOI221_X1 U2606 ( .B1(n927), .B2(\registers[13][0] ), .C1(n924), .C2(
        \registers[12][0] ), .A(n2769), .ZN(n2742) );
  AOI211_X1 U2607 ( .C1(n1012), .C2(\registers[1][0] ), .A(n2763), .B(n2764), 
        .ZN(n2743) );
  NAND4_X1 U2608 ( .A1(n2724), .A2(n2725), .A3(n2726), .A4(n2727), .ZN(N187)
         );
  AOI221_X1 U2609 ( .B1(n915), .B2(\registers[9][1] ), .C1(n912), .C2(
        \registers[8][1] ), .A(n2740), .ZN(n2724) );
  AOI221_X1 U2610 ( .B1(n927), .B2(\registers[13][1] ), .C1(n924), .C2(
        \registers[12][1] ), .A(n2739), .ZN(n2725) );
  AOI211_X1 U2611 ( .C1(n1012), .C2(\registers[1][1] ), .A(n2736), .B(n2737), 
        .ZN(n2726) );
  NAND4_X1 U2612 ( .A1(n2707), .A2(n2708), .A3(n2709), .A4(n2710), .ZN(N188)
         );
  AOI221_X1 U2613 ( .B1(n915), .B2(\registers[9][2] ), .C1(n912), .C2(
        \registers[8][2] ), .A(n2723), .ZN(n2707) );
  AOI221_X1 U2614 ( .B1(n927), .B2(\registers[13][2] ), .C1(n924), .C2(
        \registers[12][2] ), .A(n2722), .ZN(n2708) );
  AOI211_X1 U2615 ( .C1(n1012), .C2(\registers[1][2] ), .A(n2719), .B(n2720), 
        .ZN(n2709) );
  NAND4_X1 U2616 ( .A1(n2690), .A2(n2691), .A3(n2692), .A4(n2693), .ZN(N189)
         );
  AOI221_X1 U2617 ( .B1(n915), .B2(\registers[9][3] ), .C1(n912), .C2(
        \registers[8][3] ), .A(n2706), .ZN(n2690) );
  AOI221_X1 U2618 ( .B1(n927), .B2(\registers[13][3] ), .C1(n924), .C2(
        \registers[12][3] ), .A(n2705), .ZN(n2691) );
  AOI211_X1 U2619 ( .C1(n1012), .C2(\registers[1][3] ), .A(n2702), .B(n2703), 
        .ZN(n2692) );
  NAND4_X1 U2620 ( .A1(n2673), .A2(n2674), .A3(n2675), .A4(n2676), .ZN(N190)
         );
  AOI221_X1 U2621 ( .B1(n915), .B2(\registers[9][4] ), .C1(n912), .C2(
        \registers[8][4] ), .A(n2689), .ZN(n2673) );
  AOI221_X1 U2622 ( .B1(n927), .B2(\registers[13][4] ), .C1(n924), .C2(
        \registers[12][4] ), .A(n2688), .ZN(n2674) );
  AOI211_X1 U2623 ( .C1(n1012), .C2(\registers[1][4] ), .A(n2685), .B(n2686), 
        .ZN(n2675) );
  NAND4_X1 U2624 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(N191)
         );
  AOI221_X1 U2625 ( .B1(n915), .B2(\registers[9][5] ), .C1(n912), .C2(
        \registers[8][5] ), .A(n2672), .ZN(n2656) );
  AOI221_X1 U2626 ( .B1(n927), .B2(\registers[13][5] ), .C1(n924), .C2(
        \registers[12][5] ), .A(n2671), .ZN(n2657) );
  AOI211_X1 U2627 ( .C1(n1012), .C2(\registers[1][5] ), .A(n2668), .B(n2669), 
        .ZN(n2658) );
  NAND4_X1 U2628 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2642), .ZN(N192)
         );
  AOI221_X1 U2629 ( .B1(n915), .B2(\registers[9][6] ), .C1(n912), .C2(
        \registers[8][6] ), .A(n2655), .ZN(n2639) );
  AOI221_X1 U2630 ( .B1(n927), .B2(\registers[13][6] ), .C1(n924), .C2(
        \registers[12][6] ), .A(n2654), .ZN(n2640) );
  AOI211_X1 U2631 ( .C1(n1012), .C2(\registers[1][6] ), .A(n2651), .B(n2652), 
        .ZN(n2641) );
  NAND4_X1 U2632 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(N193)
         );
  AOI221_X1 U2633 ( .B1(n915), .B2(\registers[9][7] ), .C1(n912), .C2(
        \registers[8][7] ), .A(n2638), .ZN(n2622) );
  AOI221_X1 U2634 ( .B1(n927), .B2(\registers[13][7] ), .C1(n924), .C2(
        \registers[12][7] ), .A(n2637), .ZN(n2623) );
  AOI211_X1 U2635 ( .C1(n1012), .C2(\registers[1][7] ), .A(n2634), .B(n2635), 
        .ZN(n2624) );
  NAND4_X1 U2636 ( .A1(n2605), .A2(n2606), .A3(n2607), .A4(n2608), .ZN(N194)
         );
  AOI221_X1 U2637 ( .B1(n915), .B2(\registers[9][8] ), .C1(n912), .C2(
        \registers[8][8] ), .A(n2621), .ZN(n2605) );
  AOI221_X1 U2638 ( .B1(n927), .B2(\registers[13][8] ), .C1(n924), .C2(
        \registers[12][8] ), .A(n2620), .ZN(n2606) );
  AOI211_X1 U2639 ( .C1(n1012), .C2(\registers[1][8] ), .A(n2617), .B(n2618), 
        .ZN(n2607) );
  NAND4_X1 U2640 ( .A1(n2588), .A2(n2589), .A3(n2590), .A4(n2591), .ZN(N195)
         );
  AOI221_X1 U2641 ( .B1(n915), .B2(\registers[9][9] ), .C1(n912), .C2(
        \registers[8][9] ), .A(n2604), .ZN(n2588) );
  AOI221_X1 U2642 ( .B1(n927), .B2(\registers[13][9] ), .C1(n924), .C2(
        \registers[12][9] ), .A(n2603), .ZN(n2589) );
  AOI211_X1 U2643 ( .C1(n1012), .C2(\registers[1][9] ), .A(n2600), .B(n2601), 
        .ZN(n2590) );
  NAND4_X1 U2644 ( .A1(n2571), .A2(n2572), .A3(n2573), .A4(n2574), .ZN(N196)
         );
  AOI221_X1 U2645 ( .B1(n915), .B2(\registers[9][10] ), .C1(n912), .C2(
        \registers[8][10] ), .A(n2587), .ZN(n2571) );
  AOI221_X1 U2646 ( .B1(n927), .B2(\registers[13][10] ), .C1(n924), .C2(
        \registers[12][10] ), .A(n2586), .ZN(n2572) );
  AOI211_X1 U2647 ( .C1(n1012), .C2(\registers[1][10] ), .A(n2583), .B(n2584), 
        .ZN(n2573) );
  NAND4_X1 U2648 ( .A1(n2554), .A2(n2555), .A3(n2556), .A4(n2557), .ZN(N197)
         );
  AOI221_X1 U2649 ( .B1(n916), .B2(\registers[9][11] ), .C1(n913), .C2(
        \registers[8][11] ), .A(n2570), .ZN(n2554) );
  AOI221_X1 U2650 ( .B1(n928), .B2(\registers[13][11] ), .C1(n925), .C2(
        \registers[12][11] ), .A(n2569), .ZN(n2555) );
  AOI211_X1 U2651 ( .C1(n1013), .C2(\registers[1][11] ), .A(n2566), .B(n2567), 
        .ZN(n2556) );
  NAND4_X1 U2652 ( .A1(n2537), .A2(n2538), .A3(n2539), .A4(n2540), .ZN(N198)
         );
  AOI221_X1 U2653 ( .B1(n916), .B2(\registers[9][12] ), .C1(n913), .C2(
        \registers[8][12] ), .A(n2553), .ZN(n2537) );
  AOI221_X1 U2654 ( .B1(n928), .B2(\registers[13][12] ), .C1(n925), .C2(
        \registers[12][12] ), .A(n2552), .ZN(n2538) );
  AOI211_X1 U2655 ( .C1(n1013), .C2(\registers[1][12] ), .A(n2549), .B(n2550), 
        .ZN(n2539) );
  NAND4_X1 U2656 ( .A1(n2520), .A2(n2521), .A3(n2522), .A4(n2523), .ZN(N199)
         );
  AOI221_X1 U2657 ( .B1(n916), .B2(\registers[9][13] ), .C1(n913), .C2(
        \registers[8][13] ), .A(n2536), .ZN(n2520) );
  AOI221_X1 U2658 ( .B1(n928), .B2(\registers[13][13] ), .C1(n925), .C2(
        \registers[12][13] ), .A(n2535), .ZN(n2521) );
  AOI211_X1 U2659 ( .C1(n1013), .C2(\registers[1][13] ), .A(n2532), .B(n2533), 
        .ZN(n2522) );
  NAND4_X1 U2660 ( .A1(n2503), .A2(n2504), .A3(n2505), .A4(n2506), .ZN(N200)
         );
  AOI221_X1 U2661 ( .B1(n916), .B2(\registers[9][14] ), .C1(n913), .C2(
        \registers[8][14] ), .A(n2519), .ZN(n2503) );
  AOI221_X1 U2662 ( .B1(n928), .B2(\registers[13][14] ), .C1(n925), .C2(
        \registers[12][14] ), .A(n2518), .ZN(n2504) );
  AOI211_X1 U2663 ( .C1(n1013), .C2(\registers[1][14] ), .A(n2515), .B(n2516), 
        .ZN(n2505) );
  NAND4_X1 U2664 ( .A1(n2486), .A2(n2487), .A3(n2488), .A4(n2489), .ZN(N201)
         );
  AOI221_X1 U2665 ( .B1(n916), .B2(\registers[9][15] ), .C1(n913), .C2(
        \registers[8][15] ), .A(n2502), .ZN(n2486) );
  AOI221_X1 U2666 ( .B1(n928), .B2(\registers[13][15] ), .C1(n925), .C2(
        \registers[12][15] ), .A(n2501), .ZN(n2487) );
  AOI211_X1 U2667 ( .C1(n1013), .C2(\registers[1][15] ), .A(n2498), .B(n2499), 
        .ZN(n2488) );
  NAND4_X1 U2668 ( .A1(n2469), .A2(n2470), .A3(n2471), .A4(n2472), .ZN(N202)
         );
  AOI221_X1 U2669 ( .B1(n916), .B2(\registers[9][16] ), .C1(n913), .C2(
        \registers[8][16] ), .A(n2485), .ZN(n2469) );
  AOI221_X1 U2670 ( .B1(n928), .B2(\registers[13][16] ), .C1(n925), .C2(
        \registers[12][16] ), .A(n2484), .ZN(n2470) );
  AOI211_X1 U2671 ( .C1(n1013), .C2(\registers[1][16] ), .A(n2481), .B(n2482), 
        .ZN(n2471) );
  NAND4_X1 U2672 ( .A1(n2452), .A2(n2453), .A3(n2454), .A4(n2455), .ZN(N203)
         );
  AOI221_X1 U2673 ( .B1(n916), .B2(\registers[9][17] ), .C1(n913), .C2(
        \registers[8][17] ), .A(n2468), .ZN(n2452) );
  AOI221_X1 U2674 ( .B1(n928), .B2(\registers[13][17] ), .C1(n925), .C2(
        \registers[12][17] ), .A(n2467), .ZN(n2453) );
  AOI211_X1 U2675 ( .C1(n1013), .C2(\registers[1][17] ), .A(n2464), .B(n2465), 
        .ZN(n2454) );
  NAND4_X1 U2676 ( .A1(n2435), .A2(n2436), .A3(n2437), .A4(n2438), .ZN(N204)
         );
  AOI221_X1 U2677 ( .B1(n916), .B2(\registers[9][18] ), .C1(n913), .C2(
        \registers[8][18] ), .A(n2451), .ZN(n2435) );
  AOI221_X1 U2678 ( .B1(n928), .B2(\registers[13][18] ), .C1(n925), .C2(
        \registers[12][18] ), .A(n2450), .ZN(n2436) );
  AOI211_X1 U2679 ( .C1(n1013), .C2(\registers[1][18] ), .A(n2447), .B(n2448), 
        .ZN(n2437) );
  NAND4_X1 U2680 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(N205)
         );
  AOI221_X1 U2681 ( .B1(n916), .B2(\registers[9][19] ), .C1(n913), .C2(
        \registers[8][19] ), .A(n2434), .ZN(n2418) );
  AOI221_X1 U2682 ( .B1(n928), .B2(\registers[13][19] ), .C1(n925), .C2(
        \registers[12][19] ), .A(n2433), .ZN(n2419) );
  AOI211_X1 U2683 ( .C1(n1013), .C2(\registers[1][19] ), .A(n2430), .B(n2431), 
        .ZN(n2420) );
  NAND4_X1 U2684 ( .A1(n2401), .A2(n2402), .A3(n2403), .A4(n2404), .ZN(N206)
         );
  AOI221_X1 U2685 ( .B1(n916), .B2(\registers[9][20] ), .C1(n913), .C2(
        \registers[8][20] ), .A(n2417), .ZN(n2401) );
  AOI221_X1 U2686 ( .B1(n928), .B2(\registers[13][20] ), .C1(n925), .C2(
        \registers[12][20] ), .A(n2416), .ZN(n2402) );
  AOI211_X1 U2687 ( .C1(n1013), .C2(\registers[1][20] ), .A(n2413), .B(n2414), 
        .ZN(n2403) );
  NAND4_X1 U2688 ( .A1(n2384), .A2(n2385), .A3(n2386), .A4(n2387), .ZN(N207)
         );
  AOI221_X1 U2689 ( .B1(n916), .B2(\registers[9][21] ), .C1(n913), .C2(
        \registers[8][21] ), .A(n2400), .ZN(n2384) );
  AOI221_X1 U2690 ( .B1(n928), .B2(\registers[13][21] ), .C1(n925), .C2(
        \registers[12][21] ), .A(n2399), .ZN(n2385) );
  AOI211_X1 U2691 ( .C1(n1013), .C2(\registers[1][21] ), .A(n2396), .B(n2397), 
        .ZN(n2386) );
  NOR2_X1 U2692 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n2177) );
  NOR2_X1 U2693 ( .A1(n4177), .A2(ADD_RD2[4]), .ZN(n2182) );
  NOR2_X1 U2694 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n2768) );
  NOR2_X1 U2695 ( .A1(n4174), .A2(ADD_RD1[4]), .ZN(n2773) );
  AND2_X1 U2696 ( .A1(n2166), .A2(ADD_RD2[0]), .ZN(n2161) );
  AND2_X1 U2697 ( .A1(n2177), .A2(ADD_RD2[0]), .ZN(n2174) );
  AND2_X1 U2698 ( .A1(n2182), .A2(ADD_RD2[0]), .ZN(n2179) );
  AND2_X1 U2699 ( .A1(n2757), .A2(ADD_RD1[0]), .ZN(n2752) );
  AND2_X1 U2700 ( .A1(n2768), .A2(ADD_RD1[0]), .ZN(n2765) );
  AND2_X1 U2701 ( .A1(n2773), .A2(ADD_RD1[0]), .ZN(n2770) );
  INV_X1 U2702 ( .A(ADD_RD2[0]), .ZN(n4179) );
  INV_X1 U2703 ( .A(ADD_RD1[0]), .ZN(n4176) );
  INV_X1 U2704 ( .A(ADD_RD2[3]), .ZN(n4177) );
  INV_X1 U2705 ( .A(ADD_RD2[1]), .ZN(n4178) );
  INV_X1 U2706 ( .A(ADD_RD1[3]), .ZN(n4174) );
  INV_X1 U2707 ( .A(ADD_RD1[1]), .ZN(n4175) );
  AND2_X1 U2708 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n2171) );
  AND2_X1 U2709 ( .A1(ADD_RD2[4]), .A2(n4177), .ZN(n2166) );
  AND2_X1 U2710 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2762) );
  AND2_X1 U2711 ( .A1(ADD_RD1[4]), .A2(n4174), .ZN(n2757) );
  INV_X1 U2712 ( .A(n1073), .ZN(n4138) );
  AOI22_X1 U2713 ( .A1(n754), .A2(DATAIN[0]), .B1(n3572), .B2(
        \registers[29][0] ), .ZN(n1073) );
  INV_X1 U2714 ( .A(n1075), .ZN(n4139) );
  AOI22_X1 U2715 ( .A1(n892), .A2(n3566), .B1(n3570), .B2(\registers[29][1] ), 
        .ZN(n1075) );
  INV_X1 U2716 ( .A(n1076), .ZN(n4140) );
  AOI22_X1 U2717 ( .A1(n375), .A2(n3565), .B1(n3567), .B2(\registers[29][2] ), 
        .ZN(n1076) );
  INV_X1 U2718 ( .A(n1077), .ZN(n4141) );
  AOI22_X1 U2719 ( .A1(n800), .A2(n3565), .B1(n554), .B2(\registers[29][3] ), 
        .ZN(n1077) );
  INV_X1 U2720 ( .A(n1078), .ZN(n4142) );
  AOI22_X1 U2721 ( .A1(n590), .A2(n745), .B1(n554), .B2(\registers[29][4] ), 
        .ZN(n1078) );
  INV_X1 U2722 ( .A(n1079), .ZN(n4143) );
  AOI22_X1 U2723 ( .A1(n798), .A2(n3565), .B1(n3567), .B2(\registers[29][5] ), 
        .ZN(n1079) );
  INV_X1 U2724 ( .A(n1080), .ZN(n4144) );
  AOI22_X1 U2725 ( .A1(n228), .A2(n3564), .B1(n554), .B2(\registers[29][6] ), 
        .ZN(n1080) );
  INV_X1 U2726 ( .A(n1081), .ZN(n4145) );
  AOI22_X1 U2727 ( .A1(n199), .A2(n3566), .B1(n3569), .B2(\registers[29][7] ), 
        .ZN(n1081) );
  INV_X1 U2728 ( .A(n1107), .ZN(n4107) );
  AOI22_X1 U2729 ( .A1(DATAIN[0]), .A2(n545), .B1(n229), .B2(
        \registers[28][0] ), .ZN(n1107) );
  INV_X1 U2730 ( .A(n1109), .ZN(n4108) );
  AOI22_X1 U2731 ( .A1(n892), .A2(n395), .B1(n3561), .B2(\registers[28][1] ), 
        .ZN(n1109) );
  INV_X1 U2732 ( .A(n1110), .ZN(n4109) );
  AOI22_X1 U2733 ( .A1(n890), .A2(n545), .B1(n229), .B2(\registers[28][2] ), 
        .ZN(n1110) );
  INV_X1 U2734 ( .A(n1111), .ZN(n4110) );
  AOI22_X1 U2735 ( .A1(n800), .A2(n3559), .B1(n229), .B2(\registers[28][3] ), 
        .ZN(n1111) );
  INV_X1 U2736 ( .A(n1112), .ZN(n4111) );
  AOI22_X1 U2737 ( .A1(n545), .A2(n882), .B1(n229), .B2(\registers[28][4] ), 
        .ZN(n1112) );
  INV_X1 U2738 ( .A(n1114), .ZN(n4112) );
  AOI22_X1 U2739 ( .A1(n881), .A2(n3559), .B1(n182), .B2(\registers[28][6] ), 
        .ZN(n1114) );
  INV_X1 U2740 ( .A(n1115), .ZN(n4113) );
  AOI22_X1 U2741 ( .A1(n3558), .A2(n796), .B1(n3562), .B2(\registers[28][7] ), 
        .ZN(n1115) );
  INV_X1 U2742 ( .A(n1145), .ZN(n4075) );
  AOI22_X1 U2743 ( .A1(DATAIN[0]), .A2(n3534), .B1(n386), .B2(
        \registers[25][0] ), .ZN(n1145) );
  INV_X1 U2744 ( .A(n1147), .ZN(n4076) );
  AOI22_X1 U2745 ( .A1(n892), .A2(n719), .B1(n3536), .B2(\registers[25][1] ), 
        .ZN(n1147) );
  INV_X1 U2746 ( .A(n1148), .ZN(n4077) );
  AOI22_X1 U2747 ( .A1(n375), .A2(n3534), .B1(n386), .B2(\registers[25][2] ), 
        .ZN(n1148) );
  INV_X1 U2748 ( .A(n1149), .ZN(n4078) );
  AOI22_X1 U2749 ( .A1(n800), .A2(n3533), .B1(n386), .B2(\registers[25][3] ), 
        .ZN(n1149) );
  INV_X1 U2750 ( .A(n1150), .ZN(n4079) );
  AOI22_X1 U2751 ( .A1(n882), .A2(n762), .B1(n386), .B2(\registers[25][4] ), 
        .ZN(n1150) );
  INV_X1 U2752 ( .A(n1151), .ZN(n4080) );
  AOI22_X1 U2753 ( .A1(n798), .A2(n719), .B1(n386), .B2(\registers[25][5] ), 
        .ZN(n1151) );
  INV_X1 U2754 ( .A(n1152), .ZN(n4081) );
  AOI22_X1 U2755 ( .A1(n881), .A2(n762), .B1(n386), .B2(\registers[25][6] ), 
        .ZN(n1152) );
  INV_X1 U2756 ( .A(n1153), .ZN(n4082) );
  AOI22_X1 U2757 ( .A1(n31), .A2(n198), .B1(n3535), .B2(\registers[25][7] ), 
        .ZN(n1153) );
  INV_X1 U2758 ( .A(n1214), .ZN(n4011) );
  AOI22_X1 U2759 ( .A1(DATAIN[0]), .A2(n3517), .B1(n3521), .B2(
        \registers[23][0] ), .ZN(n1214) );
  INV_X1 U2760 ( .A(n1216), .ZN(n4012) );
  AOI22_X1 U2761 ( .A1(n892), .A2(n750), .B1(n3521), .B2(\registers[23][1] ), 
        .ZN(n1216) );
  INV_X1 U2762 ( .A(n1217), .ZN(n4013) );
  AOI22_X1 U2763 ( .A1(n375), .A2(n3518), .B1(n3520), .B2(\registers[23][2] ), 
        .ZN(n1217) );
  INV_X1 U2764 ( .A(n1218), .ZN(n4014) );
  AOI22_X1 U2765 ( .A1(n800), .A2(n173), .B1(n3520), .B2(\registers[23][3] ), 
        .ZN(n1218) );
  INV_X1 U2766 ( .A(n1219), .ZN(n4015) );
  AOI22_X1 U2767 ( .A1(n882), .A2(n750), .B1(n3522), .B2(\registers[23][4] ), 
        .ZN(n1219) );
  INV_X1 U2768 ( .A(n1220), .ZN(n4016) );
  AOI22_X1 U2769 ( .A1(n798), .A2(n3518), .B1(n3520), .B2(\registers[23][5] ), 
        .ZN(n1220) );
  INV_X1 U2770 ( .A(n1221), .ZN(n4017) );
  AOI22_X1 U2771 ( .A1(n228), .A2(n173), .B1(n3521), .B2(\registers[23][6] ), 
        .ZN(n1221) );
  INV_X1 U2772 ( .A(n1222), .ZN(n4018) );
  AOI22_X1 U2773 ( .A1(n199), .A2(n3519), .B1(n3520), .B2(\registers[23][7] ), 
        .ZN(n1222) );
  INV_X1 U2774 ( .A(n1251), .ZN(n3986) );
  AOI22_X1 U2775 ( .A1(n890), .A2(n362), .B1(n3516), .B2(\registers[22][2] ), 
        .ZN(n1251) );
  INV_X1 U2776 ( .A(n1253), .ZN(n3987) );
  AOI22_X1 U2777 ( .A1(n362), .A2(n590), .B1(n361), .B2(\registers[22][4] ), 
        .ZN(n1253) );
  INV_X1 U2778 ( .A(n1255), .ZN(n3988) );
  AOI22_X1 U2779 ( .A1(n227), .A2(n364), .B1(n361), .B2(\registers[22][6] ), 
        .ZN(n1255) );
  INV_X1 U2780 ( .A(n1256), .ZN(n3989) );
  AOI22_X1 U2781 ( .A1(n199), .A2(n185), .B1(n3514), .B2(\registers[22][7] ), 
        .ZN(n1256) );
  INV_X1 U2782 ( .A(n1354), .ZN(n3797) );
  AOI22_X1 U2783 ( .A1(DATAIN[0]), .A2(n3441), .B1(n3444), .B2(
        \registers[13][0] ), .ZN(n1354) );
  INV_X1 U2784 ( .A(n1356), .ZN(n3798) );
  AOI22_X1 U2785 ( .A1(n892), .A2(n3439), .B1(n3444), .B2(\registers[13][1] ), 
        .ZN(n1356) );
  INV_X1 U2786 ( .A(n1358), .ZN(n3799) );
  AOI22_X1 U2787 ( .A1(n800), .A2(n391), .B1(n11), .B2(\registers[13][3] ), 
        .ZN(n1358) );
  INV_X1 U2788 ( .A(n1359), .ZN(n3800) );
  AOI22_X1 U2789 ( .A1(n718), .A2(n590), .B1(n12), .B2(\registers[13][4] ), 
        .ZN(n1359) );
  INV_X1 U2790 ( .A(n1360), .ZN(n3801) );
  AOI22_X1 U2791 ( .A1(n718), .A2(n798), .B1(n12), .B2(\registers[13][5] ), 
        .ZN(n1360) );
  INV_X1 U2792 ( .A(n1361), .ZN(n3802) );
  AOI22_X1 U2793 ( .A1(n881), .A2(n3441), .B1(n3444), .B2(\registers[13][6] ), 
        .ZN(n1361) );
  INV_X1 U2794 ( .A(n1362), .ZN(n3803) );
  AOI22_X1 U2795 ( .A1(n198), .A2(n3440), .B1(n3444), .B2(\registers[13][7] ), 
        .ZN(n1362) );
  INV_X1 U2796 ( .A(n1389), .ZN(n3769) );
  AOI22_X1 U2797 ( .A1(n892), .A2(n695), .B1(n3434), .B2(\registers[12][1] ), 
        .ZN(n1389) );
  INV_X1 U2798 ( .A(n1390), .ZN(n3770) );
  AOI22_X1 U2799 ( .A1(n375), .A2(n751), .B1(n3434), .B2(\registers[12][2] ), 
        .ZN(n1390) );
  INV_X1 U2800 ( .A(n1391), .ZN(n3771) );
  AOI22_X1 U2801 ( .A1(n800), .A2(n751), .B1(n3434), .B2(\registers[12][3] ), 
        .ZN(n1391) );
  INV_X1 U2802 ( .A(n1392), .ZN(n3772) );
  AOI22_X1 U2803 ( .A1(n882), .A2(n747), .B1(n3434), .B2(\registers[12][4] ), 
        .ZN(n1392) );
  INV_X1 U2804 ( .A(n1393), .ZN(n3773) );
  AOI22_X1 U2805 ( .A1(n798), .A2(n3433), .B1(n274), .B2(\registers[12][5] ), 
        .ZN(n1393) );
  INV_X1 U2806 ( .A(n1394), .ZN(n3774) );
  AOI22_X1 U2807 ( .A1(n696), .A2(n881), .B1(n276), .B2(\registers[12][6] ), 
        .ZN(n1394) );
  INV_X1 U2808 ( .A(n1395), .ZN(n3775) );
  AOI22_X1 U2809 ( .A1(n796), .A2(n747), .B1(n276), .B2(\registers[12][7] ), 
        .ZN(n1395) );
  INV_X1 U2810 ( .A(n1488), .ZN(n3891) );
  AOI22_X1 U2811 ( .A1(DATAIN[0]), .A2(n3390), .B1(n3391), .B2(
        \registers[7][0] ), .ZN(n1488) );
  INV_X1 U2812 ( .A(n1490), .ZN(n3892) );
  AOI22_X1 U2813 ( .A1(n892), .A2(n3390), .B1(n3391), .B2(\registers[7][1] ), 
        .ZN(n1490) );
  INV_X1 U2814 ( .A(n1491), .ZN(n3893) );
  AOI22_X1 U2815 ( .A1(n890), .A2(n358), .B1(n3391), .B2(\registers[7][2] ), 
        .ZN(n1491) );
  INV_X1 U2816 ( .A(n1492), .ZN(n3894) );
  AOI22_X1 U2817 ( .A1(n800), .A2(n3390), .B1(n3391), .B2(\registers[7][3] ), 
        .ZN(n1492) );
  INV_X1 U2818 ( .A(n1493), .ZN(n3895) );
  AOI22_X1 U2819 ( .A1(n882), .A2(n3390), .B1(n3391), .B2(\registers[7][4] ), 
        .ZN(n1493) );
  INV_X1 U2820 ( .A(n1494), .ZN(n3896) );
  AOI22_X1 U2821 ( .A1(n798), .A2(n358), .B1(n3392), .B2(\registers[7][5] ), 
        .ZN(n1494) );
  INV_X1 U2822 ( .A(n1495), .ZN(n3897) );
  AOI22_X1 U2823 ( .A1(n881), .A2(n3390), .B1(n3392), .B2(\registers[7][6] ), 
        .ZN(n1495) );
  INV_X1 U2824 ( .A(n1496), .ZN(n3898) );
  AOI22_X1 U2825 ( .A1(n199), .A2(n358), .B1(n3392), .B2(\registers[7][7] ), 
        .ZN(n1496) );
  INV_X1 U2826 ( .A(n1522), .ZN(n3859) );
  AOI22_X1 U2827 ( .A1(n3384), .A2(DATAIN[0]), .B1(n3386), .B2(
        \registers[6][0] ), .ZN(n1522) );
  INV_X1 U2828 ( .A(n1524), .ZN(n3860) );
  AOI22_X1 U2829 ( .A1(n892), .A2(n547), .B1(n3385), .B2(\registers[6][1] ), 
        .ZN(n1524) );
  INV_X1 U2830 ( .A(n1525), .ZN(n3861) );
  AOI22_X1 U2831 ( .A1(n3384), .A2(n375), .B1(n3386), .B2(\registers[6][2] ), 
        .ZN(n1525) );
  INV_X1 U2832 ( .A(n1526), .ZN(n3862) );
  AOI22_X1 U2833 ( .A1(n800), .A2(n547), .B1(n3388), .B2(\registers[6][3] ), 
        .ZN(n1526) );
  INV_X1 U2834 ( .A(n1527), .ZN(n3863) );
  AOI22_X1 U2835 ( .A1(n398), .A2(n590), .B1(n3386), .B2(\registers[6][4] ), 
        .ZN(n1527) );
  INV_X1 U2836 ( .A(n1528), .ZN(n3864) );
  AOI22_X1 U2837 ( .A1(n798), .A2(n398), .B1(n3385), .B2(\registers[6][5] ), 
        .ZN(n1528) );
  INV_X1 U2838 ( .A(n1529), .ZN(n3865) );
  AOI22_X1 U2839 ( .A1(n227), .A2(n196), .B1(n3388), .B2(\registers[6][6] ), 
        .ZN(n1529) );
  INV_X1 U2840 ( .A(n1530), .ZN(n3866) );
  AOI22_X1 U2841 ( .A1(n196), .A2(n198), .B1(n3385), .B2(\registers[6][7] ), 
        .ZN(n1530) );
  INV_X1 U2842 ( .A(n1425), .ZN(n3743) );
  AOI22_X1 U2843 ( .A1(n890), .A2(n3409), .B1(n3412), .B2(\registers[9][2] ), 
        .ZN(n1425) );
  INV_X1 U2844 ( .A(n1426), .ZN(n3744) );
  AOI22_X1 U2845 ( .A1(n800), .A2(n3408), .B1(n381), .B2(\registers[9][3] ), 
        .ZN(n1426) );
  INV_X1 U2846 ( .A(n1428), .ZN(n3745) );
  AOI22_X1 U2847 ( .A1(n798), .A2(n561), .B1(n3412), .B2(\registers[9][5] ), 
        .ZN(n1428) );
  INV_X1 U2848 ( .A(n1430), .ZN(n3746) );
  AOI22_X1 U2849 ( .A1(n796), .A2(n3408), .B1(n354), .B2(\registers[9][7] ), 
        .ZN(n1430) );
  INV_X1 U2850 ( .A(n1559), .ZN(n3827) );
  AOI22_X1 U2851 ( .A1(n165), .A2(n3338), .B1(n3340), .B2(\registers[1][0] ), 
        .ZN(n1559) );
  INV_X1 U2852 ( .A(n1561), .ZN(n3828) );
  AOI22_X1 U2853 ( .A1(n366), .A2(n892), .B1(n3340), .B2(\registers[1][1] ), 
        .ZN(n1561) );
  INV_X1 U2854 ( .A(n1562), .ZN(n3829) );
  AOI22_X1 U2855 ( .A1(n375), .A2(n366), .B1(n262), .B2(\registers[1][2] ), 
        .ZN(n1562) );
  INV_X1 U2856 ( .A(n1563), .ZN(n3830) );
  AOI22_X1 U2857 ( .A1(n800), .A2(n3338), .B1(n3340), .B2(\registers[1][3] ), 
        .ZN(n1563) );
  INV_X1 U2858 ( .A(n1564), .ZN(n3831) );
  AOI22_X1 U2859 ( .A1(n590), .A2(n3338), .B1(n3340), .B2(\registers[1][4] ), 
        .ZN(n1564) );
  INV_X1 U2860 ( .A(n1565), .ZN(n3832) );
  AOI22_X1 U2861 ( .A1(n366), .A2(n798), .B1(n262), .B2(\registers[1][5] ), 
        .ZN(n1565) );
  INV_X1 U2862 ( .A(n1566), .ZN(n3833) );
  AOI22_X1 U2863 ( .A1(n365), .A2(n228), .B1(n3340), .B2(\registers[1][6] ), 
        .ZN(n1566) );
  INV_X1 U2864 ( .A(n1567), .ZN(n3834) );
  AOI22_X1 U2865 ( .A1(n366), .A2(n199), .B1(n3340), .B2(\registers[1][7] ), 
        .ZN(n1567) );
  INV_X1 U2866 ( .A(n1283), .ZN(n3955) );
  AOI22_X1 U2867 ( .A1(n165), .A2(n725), .B1(n4), .B2(\registers[19][0] ), 
        .ZN(n1283) );
  INV_X1 U2868 ( .A(n1286), .ZN(n3956) );
  AOI22_X1 U2869 ( .A1(n890), .A2(n3486), .B1(n4), .B2(\registers[19][2] ), 
        .ZN(n1286) );
  INV_X1 U2870 ( .A(n1287), .ZN(n3957) );
  AOI22_X1 U2871 ( .A1(n800), .A2(n3487), .B1(n3), .B2(\registers[19][3] ), 
        .ZN(n1287) );
  INV_X1 U2872 ( .A(n1288), .ZN(n3958) );
  AOI22_X1 U2873 ( .A1(n882), .A2(n765), .B1(n4), .B2(\registers[19][4] ), 
        .ZN(n1288) );
  INV_X1 U2874 ( .A(n1289), .ZN(n3959) );
  AOI22_X1 U2875 ( .A1(n798), .A2(n396), .B1(n19), .B2(\registers[19][5] ), 
        .ZN(n1289) );
  INV_X1 U2876 ( .A(n1290), .ZN(n3960) );
  AOI22_X1 U2877 ( .A1(n227), .A2(n546), .B1(n19), .B2(\registers[19][6] ), 
        .ZN(n1290) );
  INV_X1 U2878 ( .A(n1291), .ZN(n3961) );
  AOI22_X1 U2879 ( .A1(n198), .A2(n3485), .B1(n19), .B2(\registers[19][7] ), 
        .ZN(n1291) );
  INV_X1 U2880 ( .A(n1316), .ZN(n3924) );
  AOI22_X1 U2881 ( .A1(DATAIN[0]), .A2(n3477), .B1(n3480), .B2(
        \registers[18][0] ), .ZN(n1316) );
  INV_X1 U2882 ( .A(n1318), .ZN(n3925) );
  AOI22_X1 U2883 ( .A1(n892), .A2(n763), .B1(n3480), .B2(\registers[18][1] ), 
        .ZN(n1318) );
  INV_X1 U2884 ( .A(n1319), .ZN(n3926) );
  AOI22_X1 U2885 ( .A1(n890), .A2(n3479), .B1(n3480), .B2(\registers[18][2] ), 
        .ZN(n1319) );
  INV_X1 U2886 ( .A(n1321), .ZN(n3927) );
  AOI22_X1 U2887 ( .A1(n590), .A2(n763), .B1(n3480), .B2(\registers[18][4] ), 
        .ZN(n1321) );
  INV_X1 U2888 ( .A(n1322), .ZN(n3928) );
  AOI22_X1 U2889 ( .A1(n798), .A2(n596), .B1(n3481), .B2(\registers[18][5] ), 
        .ZN(n1322) );
  INV_X1 U2890 ( .A(n1323), .ZN(n3929) );
  AOI22_X1 U2891 ( .A1(n730), .A2(n881), .B1(n3481), .B2(\registers[18][6] ), 
        .ZN(n1323) );
  INV_X1 U2892 ( .A(n1324), .ZN(n3930) );
  AOI22_X1 U2893 ( .A1(n729), .A2(n796), .B1(n3481), .B2(\registers[18][7] ), 
        .ZN(n1324) );
  INV_X1 U2894 ( .A(n1082), .ZN(n4146) );
  AOI22_X1 U2895 ( .A1(n204), .A2(n755), .B1(n3568), .B2(\registers[29][8] ), 
        .ZN(n1082) );
  INV_X1 U2896 ( .A(n1083), .ZN(n4147) );
  AOI22_X1 U2897 ( .A1(n589), .A2(n745), .B1(n3571), .B2(\registers[29][9] ), 
        .ZN(n1083) );
  INV_X1 U2898 ( .A(n1084), .ZN(n4148) );
  AOI22_X1 U2899 ( .A1(DATAIN[10]), .A2(n755), .B1(n3571), .B2(
        \registers[29][10] ), .ZN(n1084) );
  INV_X1 U2900 ( .A(n1085), .ZN(n4149) );
  AOI22_X1 U2901 ( .A1(DATAIN[11]), .A2(n3564), .B1(n3569), .B2(
        \registers[29][11] ), .ZN(n1085) );
  INV_X1 U2902 ( .A(n1086), .ZN(n4150) );
  AOI22_X1 U2903 ( .A1(n708), .A2(n3564), .B1(n3569), .B2(\registers[29][12] ), 
        .ZN(n1086) );
  INV_X1 U2904 ( .A(n1087), .ZN(n4151) );
  AOI22_X1 U2905 ( .A1(n706), .A2(n197), .B1(n3569), .B2(\registers[29][13] ), 
        .ZN(n1087) );
  INV_X1 U2906 ( .A(n1088), .ZN(n4152) );
  AOI22_X1 U2907 ( .A1(n704), .A2(n197), .B1(n3570), .B2(\registers[29][14] ), 
        .ZN(n1088) );
  INV_X1 U2908 ( .A(n1089), .ZN(n4153) );
  AOI22_X1 U2909 ( .A1(n702), .A2(n746), .B1(n3567), .B2(\registers[29][15] ), 
        .ZN(n1089) );
  INV_X1 U2910 ( .A(n1090), .ZN(n4154) );
  AOI22_X1 U2911 ( .A1(n712), .A2(n197), .B1(n3571), .B2(\registers[29][16] ), 
        .ZN(n1090) );
  INV_X1 U2912 ( .A(n1091), .ZN(n4155) );
  AOI22_X1 U2913 ( .A1(n710), .A2(n755), .B1(n3568), .B2(\registers[29][17] ), 
        .ZN(n1091) );
  INV_X1 U2914 ( .A(n1092), .ZN(n4156) );
  AOI22_X1 U2915 ( .A1(n700), .A2(n3566), .B1(n3567), .B2(\registers[29][18] ), 
        .ZN(n1092) );
  INV_X1 U2916 ( .A(n1093), .ZN(n4157) );
  AOI22_X1 U2917 ( .A1(n792), .A2(n746), .B1(n3571), .B2(\registers[29][19] ), 
        .ZN(n1093) );
  INV_X1 U2918 ( .A(n1094), .ZN(n4158) );
  AOI22_X1 U2919 ( .A1(n876), .A2(n745), .B1(n3568), .B2(\registers[29][20] ), 
        .ZN(n1094) );
  INV_X1 U2920 ( .A(n1095), .ZN(n4159) );
  AOI22_X1 U2921 ( .A1(n888), .A2(n746), .B1(n3568), .B2(\registers[29][21] ), 
        .ZN(n1095) );
  INV_X1 U2922 ( .A(n1096), .ZN(n4160) );
  AOI22_X1 U2923 ( .A1(n588), .A2(n754), .B1(n3570), .B2(\registers[29][22] ), 
        .ZN(n1096) );
  INV_X1 U2924 ( .A(n1097), .ZN(n4161) );
  AOI22_X1 U2925 ( .A1(n887), .A2(n3565), .B1(n3569), .B2(\registers[29][23] ), 
        .ZN(n1097) );
  INV_X1 U2926 ( .A(n1098), .ZN(n4162) );
  AOI22_X1 U2927 ( .A1(n746), .A2(n872), .B1(n3570), .B2(\registers[29][24] ), 
        .ZN(n1098) );
  INV_X1 U2928 ( .A(n1099), .ZN(n4163) );
  AOI22_X1 U2929 ( .A1(n755), .A2(n886), .B1(n3571), .B2(\registers[29][25] ), 
        .ZN(n1099) );
  INV_X1 U2930 ( .A(n1100), .ZN(n4164) );
  AOI22_X1 U2931 ( .A1(n870), .A2(n754), .B1(n554), .B2(\registers[29][26] ), 
        .ZN(n1100) );
  INV_X1 U2932 ( .A(n1101), .ZN(n4165) );
  AOI22_X1 U2933 ( .A1(n885), .A2(n3566), .B1(n554), .B2(\registers[29][27] ), 
        .ZN(n1101) );
  INV_X1 U2934 ( .A(n1102), .ZN(n4166) );
  AOI22_X1 U2935 ( .A1(n868), .A2(n754), .B1(n3567), .B2(\registers[29][28] ), 
        .ZN(n1102) );
  INV_X1 U2936 ( .A(n1103), .ZN(n4167) );
  AOI22_X1 U2937 ( .A1(n397), .A2(n197), .B1(n3568), .B2(\registers[29][29] ), 
        .ZN(n1103) );
  INV_X1 U2938 ( .A(n1104), .ZN(n4168) );
  AOI22_X1 U2939 ( .A1(n745), .A2(n288), .B1(n3572), .B2(\registers[29][30] ), 
        .ZN(n1104) );
  INV_X1 U2940 ( .A(n1105), .ZN(n4169) );
  AOI22_X1 U2941 ( .A1(n878), .A2(n3564), .B1(n3570), .B2(\registers[29][31] ), 
        .ZN(n1105) );
  INV_X1 U2942 ( .A(n1116), .ZN(n4114) );
  AOI22_X1 U2943 ( .A1(n794), .A2(n3559), .B1(n182), .B2(\registers[28][8] ), 
        .ZN(n1116) );
  INV_X1 U2944 ( .A(n1117), .ZN(n4115) );
  AOI22_X1 U2945 ( .A1(n3559), .A2(n589), .B1(n3561), .B2(\registers[28][9] ), 
        .ZN(n1117) );
  INV_X1 U2946 ( .A(n1118), .ZN(n4116) );
  AOI22_X1 U2947 ( .A1(DATAIN[10]), .A2(n3558), .B1(n231), .B2(
        \registers[28][10] ), .ZN(n1118) );
  INV_X1 U2948 ( .A(n1119), .ZN(n4117) );
  AOI22_X1 U2949 ( .A1(DATAIN[11]), .A2(n753), .B1(n3561), .B2(
        \registers[28][11] ), .ZN(n1119) );
  INV_X1 U2950 ( .A(n1120), .ZN(n4118) );
  AOI22_X1 U2951 ( .A1(n708), .A2(n395), .B1(n3562), .B2(\registers[28][12] ), 
        .ZN(n1120) );
  INV_X1 U2952 ( .A(n1121), .ZN(n4119) );
  AOI22_X1 U2953 ( .A1(n545), .A2(n706), .B1(n230), .B2(\registers[28][13] ), 
        .ZN(n1121) );
  INV_X1 U2954 ( .A(n1122), .ZN(n4120) );
  AOI22_X1 U2955 ( .A1(n3558), .A2(n704), .B1(n3561), .B2(\registers[28][14] ), 
        .ZN(n1122) );
  INV_X1 U2956 ( .A(n1123), .ZN(n4121) );
  AOI22_X1 U2957 ( .A1(n748), .A2(n702), .B1(n230), .B2(\registers[28][15] ), 
        .ZN(n1123) );
  INV_X1 U2958 ( .A(n1124), .ZN(n4122) );
  AOI22_X1 U2959 ( .A1(n712), .A2(n752), .B1(n231), .B2(\registers[28][16] ), 
        .ZN(n1124) );
  INV_X1 U2960 ( .A(n1125), .ZN(n4123) );
  AOI22_X1 U2961 ( .A1(n710), .A2(n395), .B1(n3561), .B2(\registers[28][17] ), 
        .ZN(n1125) );
  INV_X1 U2962 ( .A(n1126), .ZN(n4124) );
  AOI22_X1 U2963 ( .A1(n748), .A2(n700), .B1(n3561), .B2(\registers[28][18] ), 
        .ZN(n1126) );
  INV_X1 U2964 ( .A(n1127), .ZN(n4125) );
  AOI22_X1 U2965 ( .A1(n792), .A2(n748), .B1(n3562), .B2(\registers[28][19] ), 
        .ZN(n1127) );
  INV_X1 U2966 ( .A(n1128), .ZN(n4126) );
  AOI22_X1 U2967 ( .A1(n876), .A2(n748), .B1(n182), .B2(\registers[28][20] ), 
        .ZN(n1128) );
  INV_X1 U2968 ( .A(n1129), .ZN(n4127) );
  AOI22_X1 U2969 ( .A1(n888), .A2(n753), .B1(n3561), .B2(\registers[28][21] ), 
        .ZN(n1129) );
  INV_X1 U2970 ( .A(n1130), .ZN(n4128) );
  AOI22_X1 U2971 ( .A1(n587), .A2(n748), .B1(n182), .B2(\registers[28][22] ), 
        .ZN(n1130) );
  INV_X1 U2972 ( .A(n1131), .ZN(n4129) );
  AOI22_X1 U2973 ( .A1(n752), .A2(n371), .B1(n3561), .B2(\registers[28][23] ), 
        .ZN(n1131) );
  INV_X1 U2974 ( .A(n1132), .ZN(n4130) );
  AOI22_X1 U2975 ( .A1(n236), .A2(n752), .B1(n231), .B2(\registers[28][24] ), 
        .ZN(n1132) );
  INV_X1 U2976 ( .A(n1133), .ZN(n4131) );
  AOI22_X1 U2977 ( .A1(n545), .A2(n886), .B1(n3562), .B2(\registers[28][25] ), 
        .ZN(n1133) );
  INV_X1 U2978 ( .A(n1134), .ZN(n4132) );
  AOI22_X1 U2979 ( .A1(n870), .A2(n3558), .B1(n3562), .B2(\registers[28][26] ), 
        .ZN(n1134) );
  INV_X1 U2980 ( .A(n1135), .ZN(n4133) );
  AOI22_X1 U2981 ( .A1(n251), .A2(n395), .B1(n230), .B2(\registers[28][27] ), 
        .ZN(n1135) );
  INV_X1 U2982 ( .A(n1136), .ZN(n4134) );
  AOI22_X1 U2983 ( .A1(n3558), .A2(n250), .B1(n3561), .B2(\registers[28][28] ), 
        .ZN(n1136) );
  INV_X1 U2984 ( .A(n1137), .ZN(n4135) );
  AOI22_X1 U2985 ( .A1(n397), .A2(n753), .B1(n3561), .B2(\registers[28][29] ), 
        .ZN(n1137) );
  INV_X1 U2986 ( .A(n1138), .ZN(n4136) );
  AOI22_X1 U2987 ( .A1(n866), .A2(n3559), .B1(n231), .B2(\registers[28][30] ), 
        .ZN(n1138) );
  INV_X1 U2988 ( .A(n1139), .ZN(n4137) );
  AOI22_X1 U2989 ( .A1(n252), .A2(n752), .B1(n3562), .B2(\registers[28][31] ), 
        .ZN(n1139) );
  INV_X1 U2990 ( .A(n1154), .ZN(n4083) );
  AOI22_X1 U2991 ( .A1(n203), .A2(n3534), .B1(n3536), .B2(\registers[25][8] ), 
        .ZN(n1154) );
  INV_X1 U2992 ( .A(n1155), .ZN(n4084) );
  AOI22_X1 U2993 ( .A1(n589), .A2(n31), .B1(n386), .B2(\registers[25][9] ), 
        .ZN(n1155) );
  INV_X1 U2994 ( .A(n1156), .ZN(n4085) );
  AOI22_X1 U2995 ( .A1(DATAIN[10]), .A2(n762), .B1(n3536), .B2(
        \registers[25][10] ), .ZN(n1156) );
  INV_X1 U2996 ( .A(n1157), .ZN(n4086) );
  AOI22_X1 U2997 ( .A1(DATAIN[11]), .A2(n762), .B1(n386), .B2(
        \registers[25][11] ), .ZN(n1157) );
  INV_X1 U2998 ( .A(n1158), .ZN(n4087) );
  AOI22_X1 U2999 ( .A1(n788), .A2(n591), .B1(n3536), .B2(\registers[25][12] ), 
        .ZN(n1158) );
  INV_X1 U3000 ( .A(n1159), .ZN(n4088) );
  AOI22_X1 U3001 ( .A1(n705), .A2(n3534), .B1(n3536), .B2(\registers[25][13] ), 
        .ZN(n1159) );
  INV_X1 U3002 ( .A(n1160), .ZN(n4089) );
  AOI22_X1 U3003 ( .A1(n783), .A2(n591), .B1(n3536), .B2(\registers[25][14] ), 
        .ZN(n1160) );
  INV_X1 U3004 ( .A(n1161), .ZN(n4090) );
  AOI22_X1 U3005 ( .A1(n720), .A2(n780), .B1(n3535), .B2(\registers[25][15] ), 
        .ZN(n1161) );
  INV_X1 U3006 ( .A(n1162), .ZN(n4091) );
  AOI22_X1 U3007 ( .A1(n777), .A2(n761), .B1(n386), .B2(\registers[25][16] ), 
        .ZN(n1162) );
  INV_X1 U3008 ( .A(n1163), .ZN(n4092) );
  AOI22_X1 U3009 ( .A1(n774), .A2(n761), .B1(n3536), .B2(\registers[25][17] ), 
        .ZN(n1163) );
  INV_X1 U3010 ( .A(n1164), .ZN(n4093) );
  AOI22_X1 U3011 ( .A1(n771), .A2(n3533), .B1(n3536), .B2(\registers[25][18] ), 
        .ZN(n1164) );
  INV_X1 U3012 ( .A(n1165), .ZN(n4094) );
  AOI22_X1 U3013 ( .A1(n792), .A2(n720), .B1(n3535), .B2(\registers[25][19] ), 
        .ZN(n1165) );
  INV_X1 U3014 ( .A(n1166), .ZN(n4095) );
  AOI22_X1 U3015 ( .A1(n876), .A2(n719), .B1(n386), .B2(\registers[25][20] ), 
        .ZN(n1166) );
  INV_X1 U3016 ( .A(n1167), .ZN(n4096) );
  AOI22_X1 U3017 ( .A1(n889), .A2(n31), .B1(n3536), .B2(\registers[25][21] ), 
        .ZN(n1167) );
  INV_X1 U3018 ( .A(n1168), .ZN(n4097) );
  AOI22_X1 U3019 ( .A1(n587), .A2(n3533), .B1(n3536), .B2(\registers[25][22] ), 
        .ZN(n1168) );
  INV_X1 U3020 ( .A(n1169), .ZN(n4098) );
  AOI22_X1 U3021 ( .A1(n887), .A2(n720), .B1(n386), .B2(\registers[25][23] ), 
        .ZN(n1169) );
  INV_X1 U3022 ( .A(n1170), .ZN(n4099) );
  AOI22_X1 U3023 ( .A1(n872), .A2(n719), .B1(n386), .B2(\registers[25][24] ), 
        .ZN(n1170) );
  INV_X1 U3024 ( .A(n1171), .ZN(n4100) );
  AOI22_X1 U3025 ( .A1(n367), .A2(n31), .B1(n386), .B2(\registers[25][25] ), 
        .ZN(n1171) );
  INV_X1 U3026 ( .A(n1172), .ZN(n4101) );
  AOI22_X1 U3027 ( .A1(n870), .A2(n720), .B1(n3535), .B2(\registers[25][26] ), 
        .ZN(n1172) );
  INV_X1 U3028 ( .A(n1173), .ZN(n4102) );
  AOI22_X1 U3029 ( .A1(n885), .A2(n591), .B1(n3536), .B2(\registers[25][27] ), 
        .ZN(n1173) );
  INV_X1 U3030 ( .A(n1174), .ZN(n4103) );
  AOI22_X1 U3031 ( .A1(n868), .A2(n3533), .B1(n3536), .B2(\registers[25][28] ), 
        .ZN(n1174) );
  INV_X1 U3032 ( .A(n1175), .ZN(n4104) );
  AOI22_X1 U3033 ( .A1(n397), .A2(n761), .B1(n3536), .B2(\registers[25][29] ), 
        .ZN(n1175) );
  INV_X1 U3034 ( .A(n1176), .ZN(n4105) );
  AOI22_X1 U3035 ( .A1(n288), .A2(n591), .B1(n386), .B2(\registers[25][30] ), 
        .ZN(n1176) );
  INV_X1 U3036 ( .A(n1177), .ZN(n4106) );
  AOI22_X1 U3037 ( .A1(n878), .A2(n761), .B1(n3536), .B2(\registers[25][31] ), 
        .ZN(n1177) );
  INV_X1 U3038 ( .A(n1223), .ZN(n4019) );
  AOI22_X1 U3039 ( .A1(n204), .A2(n750), .B1(n3522), .B2(\registers[23][8] ), 
        .ZN(n1223) );
  INV_X1 U3040 ( .A(n1224), .ZN(n4020) );
  AOI22_X1 U3041 ( .A1(n879), .A2(n173), .B1(n3520), .B2(\registers[23][9] ), 
        .ZN(n1224) );
  INV_X1 U3042 ( .A(n1225), .ZN(n4021) );
  AOI22_X1 U3043 ( .A1(DATAIN[10]), .A2(n3518), .B1(n3521), .B2(
        \registers[23][10] ), .ZN(n1225) );
  INV_X1 U3044 ( .A(n1226), .ZN(n4022) );
  AOI22_X1 U3045 ( .A1(DATAIN[11]), .A2(n749), .B1(n3522), .B2(
        \registers[23][11] ), .ZN(n1226) );
  INV_X1 U3046 ( .A(n1227), .ZN(n4023) );
  AOI22_X1 U3047 ( .A1(n708), .A2(n3517), .B1(n3522), .B2(\registers[23][12] ), 
        .ZN(n1227) );
  INV_X1 U3048 ( .A(n1228), .ZN(n4024) );
  AOI22_X1 U3049 ( .A1(n706), .A2(n749), .B1(n3520), .B2(\registers[23][13] ), 
        .ZN(n1228) );
  INV_X1 U3050 ( .A(n1229), .ZN(n4025) );
  AOI22_X1 U3051 ( .A1(n704), .A2(n173), .B1(n3522), .B2(\registers[23][14] ), 
        .ZN(n1229) );
  INV_X1 U3052 ( .A(n1230), .ZN(n4026) );
  AOI22_X1 U3053 ( .A1(n702), .A2(n173), .B1(n3520), .B2(\registers[23][15] ), 
        .ZN(n1230) );
  INV_X1 U3054 ( .A(n1231), .ZN(n4027) );
  AOI22_X1 U3055 ( .A1(n712), .A2(n749), .B1(n3520), .B2(\registers[23][16] ), 
        .ZN(n1231) );
  INV_X1 U3056 ( .A(n1232), .ZN(n4028) );
  AOI22_X1 U3057 ( .A1(n710), .A2(n749), .B1(n3521), .B2(\registers[23][17] ), 
        .ZN(n1232) );
  INV_X1 U3058 ( .A(n1233), .ZN(n4029) );
  AOI22_X1 U3059 ( .A1(n700), .A2(n3519), .B1(n3522), .B2(\registers[23][18] ), 
        .ZN(n1233) );
  INV_X1 U3060 ( .A(n1234), .ZN(n4030) );
  AOI22_X1 U3061 ( .A1(n792), .A2(n750), .B1(n3522), .B2(\registers[23][19] ), 
        .ZN(n1234) );
  INV_X1 U3062 ( .A(n1235), .ZN(n4031) );
  AOI22_X1 U3063 ( .A1(n875), .A2(n3519), .B1(n3522), .B2(\registers[23][20] ), 
        .ZN(n1235) );
  INV_X1 U3064 ( .A(n1236), .ZN(n4032) );
  AOI22_X1 U3065 ( .A1(n888), .A2(n3519), .B1(n3521), .B2(\registers[23][21] ), 
        .ZN(n1236) );
  INV_X1 U3066 ( .A(n1237), .ZN(n4033) );
  AOI22_X1 U3067 ( .A1(n586), .A2(n749), .B1(n3520), .B2(\registers[23][22] ), 
        .ZN(n1237) );
  INV_X1 U3068 ( .A(n1238), .ZN(n4034) );
  AOI22_X1 U3069 ( .A1(n371), .A2(n3517), .B1(n3521), .B2(\registers[23][23] ), 
        .ZN(n1238) );
  INV_X1 U3070 ( .A(n1239), .ZN(n4035) );
  AOI22_X1 U3071 ( .A1(n236), .A2(n3517), .B1(n3520), .B2(\registers[23][24] ), 
        .ZN(n1239) );
  INV_X1 U3072 ( .A(n1240), .ZN(n4036) );
  AOI22_X1 U3073 ( .A1(n886), .A2(n173), .B1(n3522), .B2(\registers[23][25] ), 
        .ZN(n1240) );
  INV_X1 U3074 ( .A(n1241), .ZN(n4037) );
  AOI22_X1 U3075 ( .A1(n870), .A2(n3519), .B1(n3522), .B2(\registers[23][26] ), 
        .ZN(n1241) );
  INV_X1 U3076 ( .A(n1242), .ZN(n4038) );
  AOI22_X1 U3077 ( .A1(n251), .A2(n3518), .B1(n3521), .B2(\registers[23][27] ), 
        .ZN(n1242) );
  INV_X1 U3078 ( .A(n1243), .ZN(n4039) );
  AOI22_X1 U3079 ( .A1(n250), .A2(n3518), .B1(n3522), .B2(\registers[23][28] ), 
        .ZN(n1243) );
  INV_X1 U3080 ( .A(n1244), .ZN(n4040) );
  AOI22_X1 U3081 ( .A1(n397), .A2(n3518), .B1(n3521), .B2(\registers[23][29] ), 
        .ZN(n1244) );
  INV_X1 U3082 ( .A(n1245), .ZN(n4041) );
  AOI22_X1 U3083 ( .A1(n288), .A2(n3517), .B1(n3521), .B2(\registers[23][30] ), 
        .ZN(n1245) );
  INV_X1 U3084 ( .A(n1246), .ZN(n4042) );
  AOI22_X1 U3085 ( .A1(n252), .A2(n750), .B1(n3520), .B2(\registers[23][31] ), 
        .ZN(n1246) );
  INV_X1 U3086 ( .A(n1257), .ZN(n3990) );
  AOI22_X1 U3087 ( .A1(n194), .A2(n794), .B1(n3515), .B2(\registers[22][8] ), 
        .ZN(n1257) );
  INV_X1 U3088 ( .A(n1259), .ZN(n3991) );
  AOI22_X1 U3089 ( .A1(n363), .A2(DATAIN[10]), .B1(n211), .B2(
        \registers[22][10] ), .ZN(n1259) );
  INV_X1 U3090 ( .A(n1260), .ZN(n3992) );
  AOI22_X1 U3091 ( .A1(n184), .A2(DATAIN[11]), .B1(n211), .B2(
        \registers[22][11] ), .ZN(n1260) );
  INV_X1 U3092 ( .A(n1261), .ZN(n3993) );
  AOI22_X1 U3093 ( .A1(n708), .A2(n184), .B1(n3514), .B2(\registers[22][12] ), 
        .ZN(n1261) );
  INV_X1 U3094 ( .A(n1262), .ZN(n3994) );
  AOI22_X1 U3095 ( .A1(n194), .A2(n706), .B1(n387), .B2(\registers[22][13] ), 
        .ZN(n1262) );
  INV_X1 U3096 ( .A(n1263), .ZN(n3995) );
  AOI22_X1 U3097 ( .A1(n704), .A2(n185), .B1(n3514), .B2(\registers[22][14] ), 
        .ZN(n1263) );
  INV_X1 U3098 ( .A(n1264), .ZN(n3996) );
  AOI22_X1 U3099 ( .A1(n702), .A2(n185), .B1(n3516), .B2(\registers[22][15] ), 
        .ZN(n1264) );
  INV_X1 U3100 ( .A(n1265), .ZN(n3997) );
  AOI22_X1 U3101 ( .A1(n712), .A2(n364), .B1(n361), .B2(\registers[22][16] ), 
        .ZN(n1265) );
  INV_X1 U3102 ( .A(n1267), .ZN(n3998) );
  AOI22_X1 U3103 ( .A1(n700), .A2(n388), .B1(n3516), .B2(\registers[22][18] ), 
        .ZN(n1267) );
  INV_X1 U3104 ( .A(n1268), .ZN(n3999) );
  AOI22_X1 U3105 ( .A1(n792), .A2(n184), .B1(n3514), .B2(\registers[22][19] ), 
        .ZN(n1268) );
  INV_X1 U3106 ( .A(n1269), .ZN(n4000) );
  AOI22_X1 U3107 ( .A1(n876), .A2(n3513), .B1(n361), .B2(\registers[22][20] ), 
        .ZN(n1269) );
  INV_X1 U3108 ( .A(n1270), .ZN(n4001) );
  AOI22_X1 U3109 ( .A1(n888), .A2(n3513), .B1(n3515), .B2(\registers[22][21] ), 
        .ZN(n1270) );
  INV_X1 U3110 ( .A(n1271), .ZN(n4002) );
  AOI22_X1 U3111 ( .A1(n374), .A2(n3513), .B1(n3515), .B2(\registers[22][22] ), 
        .ZN(n1271) );
  INV_X1 U3112 ( .A(n1272), .ZN(n4003) );
  AOI22_X1 U3113 ( .A1(n887), .A2(n3513), .B1(n211), .B2(\registers[22][23] ), 
        .ZN(n1272) );
  INV_X1 U3114 ( .A(n1273), .ZN(n4004) );
  AOI22_X1 U3115 ( .A1(n872), .A2(n388), .B1(n3516), .B2(\registers[22][24] ), 
        .ZN(n1273) );
  INV_X1 U3116 ( .A(n1274), .ZN(n4005) );
  AOI22_X1 U3117 ( .A1(n367), .A2(n388), .B1(n3516), .B2(\registers[22][25] ), 
        .ZN(n1274) );
  INV_X1 U3118 ( .A(n1275), .ZN(n4006) );
  AOI22_X1 U3119 ( .A1(n870), .A2(n388), .B1(n3515), .B2(\registers[22][26] ), 
        .ZN(n1275) );
  INV_X1 U3120 ( .A(n1276), .ZN(n4007) );
  AOI22_X1 U3121 ( .A1(n885), .A2(n388), .B1(n387), .B2(\registers[22][27] ), 
        .ZN(n1276) );
  INV_X1 U3122 ( .A(n1277), .ZN(n4008) );
  AOI22_X1 U3123 ( .A1(n868), .A2(n388), .B1(n361), .B2(\registers[22][28] ), 
        .ZN(n1277) );
  INV_X1 U3124 ( .A(n1278), .ZN(n4009) );
  AOI22_X1 U3125 ( .A1(n397), .A2(n3513), .B1(n211), .B2(\registers[22][29] ), 
        .ZN(n1278) );
  INV_X1 U3126 ( .A(n1279), .ZN(n4010) );
  AOI22_X1 U3127 ( .A1(n190), .A2(n3513), .B1(n387), .B2(\registers[22][30] ), 
        .ZN(n1279) );
  INV_X1 U3128 ( .A(n1363), .ZN(n3804) );
  AOI22_X1 U3129 ( .A1(n204), .A2(n3441), .B1(n3443), .B2(\registers[13][8] ), 
        .ZN(n1363) );
  INV_X1 U3130 ( .A(n1364), .ZN(n3805) );
  AOI22_X1 U3131 ( .A1(n589), .A2(n391), .B1(n3444), .B2(\registers[13][9] ), 
        .ZN(n1364) );
  INV_X1 U3132 ( .A(n1365), .ZN(n3806) );
  AOI22_X1 U3133 ( .A1(n717), .A2(DATAIN[10]), .B1(n12), .B2(
        \registers[13][10] ), .ZN(n1365) );
  INV_X1 U3134 ( .A(n1366), .ZN(n3807) );
  AOI22_X1 U3135 ( .A1(n717), .A2(DATAIN[11]), .B1(n12), .B2(
        \registers[13][11] ), .ZN(n1366) );
  INV_X1 U3136 ( .A(n1368), .ZN(n3808) );
  AOI22_X1 U3137 ( .A1(n706), .A2(n3440), .B1(n3443), .B2(\registers[13][13] ), 
        .ZN(n1368) );
  INV_X1 U3138 ( .A(n1369), .ZN(n3809) );
  AOI22_X1 U3139 ( .A1(n718), .A2(n704), .B1(n13), .B2(\registers[13][14] ), 
        .ZN(n1369) );
  INV_X1 U3140 ( .A(n1370), .ZN(n3810) );
  AOI22_X1 U3141 ( .A1(n702), .A2(n3439), .B1(n13), .B2(\registers[13][15] ), 
        .ZN(n1370) );
  INV_X1 U3142 ( .A(n1371), .ZN(n3811) );
  AOI22_X1 U3143 ( .A1(n712), .A2(n3440), .B1(n3444), .B2(\registers[13][16] ), 
        .ZN(n1371) );
  INV_X1 U3144 ( .A(n1372), .ZN(n3812) );
  AOI22_X1 U3145 ( .A1(n710), .A2(n3440), .B1(n3444), .B2(\registers[13][17] ), 
        .ZN(n1372) );
  INV_X1 U3146 ( .A(n1373), .ZN(n3813) );
  AOI22_X1 U3147 ( .A1(n718), .A2(n700), .B1(n11), .B2(\registers[13][18] ), 
        .ZN(n1373) );
  INV_X1 U3148 ( .A(n1374), .ZN(n3814) );
  AOI22_X1 U3149 ( .A1(n792), .A2(n391), .B1(n3443), .B2(\registers[13][19] ), 
        .ZN(n1374) );
  INV_X1 U3150 ( .A(n1375), .ZN(n3815) );
  AOI22_X1 U3151 ( .A1(n876), .A2(n3441), .B1(n3443), .B2(\registers[13][20] ), 
        .ZN(n1375) );
  INV_X1 U3152 ( .A(n1376), .ZN(n3816) );
  AOI22_X1 U3153 ( .A1(n717), .A2(n889), .B1(n3443), .B2(\registers[13][21] ), 
        .ZN(n1376) );
  INV_X1 U3154 ( .A(n1377), .ZN(n3817) );
  AOI22_X1 U3155 ( .A1(n717), .A2(n588), .B1(n11), .B2(\registers[13][22] ), 
        .ZN(n1377) );
  INV_X1 U3156 ( .A(n1378), .ZN(n3818) );
  AOI22_X1 U3157 ( .A1(n887), .A2(n391), .B1(n3444), .B2(\registers[13][23] ), 
        .ZN(n1378) );
  INV_X1 U3158 ( .A(n1379), .ZN(n3819) );
  AOI22_X1 U3159 ( .A1(n872), .A2(n3439), .B1(n13), .B2(\registers[13][24] ), 
        .ZN(n1379) );
  INV_X1 U3160 ( .A(n1380), .ZN(n3820) );
  AOI22_X1 U3161 ( .A1(n886), .A2(n3439), .B1(n3444), .B2(\registers[13][25] ), 
        .ZN(n1380) );
  INV_X1 U3162 ( .A(n1381), .ZN(n3821) );
  AOI22_X1 U3163 ( .A1(n870), .A2(n391), .B1(n3444), .B2(\registers[13][26] ), 
        .ZN(n1381) );
  INV_X1 U3164 ( .A(n1382), .ZN(n3822) );
  AOI22_X1 U3165 ( .A1(n251), .A2(n3440), .B1(n13), .B2(\registers[13][27] ), 
        .ZN(n1382) );
  INV_X1 U3166 ( .A(n1383), .ZN(n3823) );
  AOI22_X1 U3167 ( .A1(n718), .A2(n868), .B1(n11), .B2(\registers[13][28] ), 
        .ZN(n1383) );
  INV_X1 U3168 ( .A(n1384), .ZN(n3824) );
  AOI22_X1 U3169 ( .A1(n883), .A2(n3441), .B1(n3443), .B2(\registers[13][29] ), 
        .ZN(n1384) );
  INV_X1 U3170 ( .A(n1385), .ZN(n3825) );
  AOI22_X1 U3171 ( .A1(n190), .A2(n3439), .B1(n3443), .B2(\registers[13][30] ), 
        .ZN(n1385) );
  INV_X1 U3172 ( .A(n1386), .ZN(n3826) );
  AOI22_X1 U3173 ( .A1(n717), .A2(n252), .B1(n12), .B2(\registers[13][31] ), 
        .ZN(n1386) );
  INV_X1 U3174 ( .A(n1396), .ZN(n3776) );
  AOI22_X1 U3175 ( .A1(n204), .A2(n751), .B1(n275), .B2(\registers[12][8] ), 
        .ZN(n1396) );
  INV_X1 U3176 ( .A(n1397), .ZN(n3777) );
  AOI22_X1 U3177 ( .A1(n589), .A2(n751), .B1(n181), .B2(\registers[12][9] ), 
        .ZN(n1397) );
  INV_X1 U3178 ( .A(n1398), .ZN(n3778) );
  AOI22_X1 U3179 ( .A1(DATAIN[10]), .A2(n584), .B1(n3436), .B2(
        \registers[12][10] ), .ZN(n1398) );
  INV_X1 U3180 ( .A(n1400), .ZN(n3779) );
  AOI22_X1 U3181 ( .A1(n708), .A2(n216), .B1(n3436), .B2(\registers[12][12] ), 
        .ZN(n1400) );
  INV_X1 U3182 ( .A(n1401), .ZN(n3780) );
  AOI22_X1 U3183 ( .A1(n584), .A2(n706), .B1(n3436), .B2(\registers[12][13] ), 
        .ZN(n1401) );
  INV_X1 U3184 ( .A(n1402), .ZN(n3781) );
  AOI22_X1 U3185 ( .A1(n704), .A2(n217), .B1(n3436), .B2(\registers[12][14] ), 
        .ZN(n1402) );
  INV_X1 U3186 ( .A(n1405), .ZN(n3782) );
  AOI22_X1 U3187 ( .A1(n710), .A2(n216), .B1(n220), .B2(\registers[12][17] ), 
        .ZN(n1405) );
  INV_X1 U3188 ( .A(n1406), .ZN(n3783) );
  AOI22_X1 U3189 ( .A1(n700), .A2(n695), .B1(n278), .B2(\registers[12][18] ), 
        .ZN(n1406) );
  INV_X1 U3190 ( .A(n1407), .ZN(n3784) );
  AOI22_X1 U3191 ( .A1(n792), .A2(n695), .B1(n278), .B2(\registers[12][19] ), 
        .ZN(n1407) );
  INV_X1 U3192 ( .A(n1408), .ZN(n3785) );
  AOI22_X1 U3193 ( .A1(n876), .A2(n696), .B1(n181), .B2(\registers[12][20] ), 
        .ZN(n1408) );
  INV_X1 U3194 ( .A(n1409), .ZN(n3786) );
  AOI22_X1 U3195 ( .A1(n696), .A2(n888), .B1(n3434), .B2(\registers[12][21] ), 
        .ZN(n1409) );
  INV_X1 U3196 ( .A(n1410), .ZN(n3787) );
  AOI22_X1 U3197 ( .A1(n374), .A2(n751), .B1(n274), .B2(\registers[12][22] ), 
        .ZN(n1410) );
  INV_X1 U3198 ( .A(n1411), .ZN(n3788) );
  AOI22_X1 U3199 ( .A1(n371), .A2(n3433), .B1(n277), .B2(\registers[12][23] ), 
        .ZN(n1411) );
  INV_X1 U3200 ( .A(n1412), .ZN(n3789) );
  AOI22_X1 U3201 ( .A1(n236), .A2(n695), .B1(n3436), .B2(\registers[12][24] ), 
        .ZN(n1412) );
  INV_X1 U3202 ( .A(n1413), .ZN(n3790) );
  AOI22_X1 U3203 ( .A1(n367), .A2(n3433), .B1(n3436), .B2(\registers[12][25] ), 
        .ZN(n1413) );
  INV_X1 U3204 ( .A(n1414), .ZN(n3791) );
  AOI22_X1 U3205 ( .A1(n870), .A2(n696), .B1(n220), .B2(\registers[12][26] ), 
        .ZN(n1414) );
  INV_X1 U3206 ( .A(n1415), .ZN(n3792) );
  AOI22_X1 U3207 ( .A1(n696), .A2(n885), .B1(n276), .B2(\registers[12][27] ), 
        .ZN(n1415) );
  INV_X1 U3208 ( .A(n1416), .ZN(n3793) );
  AOI22_X1 U3209 ( .A1(n696), .A2(n250), .B1(n274), .B2(\registers[12][28] ), 
        .ZN(n1416) );
  INV_X1 U3210 ( .A(n1417), .ZN(n3794) );
  AOI22_X1 U3211 ( .A1(n883), .A2(n217), .B1(n3436), .B2(\registers[12][29] ), 
        .ZN(n1417) );
  INV_X1 U3212 ( .A(n1418), .ZN(n3795) );
  AOI22_X1 U3213 ( .A1(n866), .A2(n3433), .B1(n275), .B2(\registers[12][30] ), 
        .ZN(n1418) );
  INV_X1 U3214 ( .A(n1419), .ZN(n3796) );
  AOI22_X1 U3215 ( .A1(n878), .A2(n3433), .B1(n275), .B2(\registers[12][31] ), 
        .ZN(n1419) );
  INV_X1 U3216 ( .A(n1497), .ZN(n3899) );
  AOI22_X1 U3217 ( .A1(n203), .A2(n3389), .B1(n3392), .B2(\registers[7][8] ), 
        .ZN(n1497) );
  INV_X1 U3218 ( .A(n1498), .ZN(n3900) );
  AOI22_X1 U3219 ( .A1(n879), .A2(n3389), .B1(n3392), .B2(\registers[7][9] ), 
        .ZN(n1498) );
  INV_X1 U3220 ( .A(n1499), .ZN(n3901) );
  AOI22_X1 U3221 ( .A1(DATAIN[10]), .A2(n3389), .B1(n3393), .B2(
        \registers[7][10] ), .ZN(n1499) );
  INV_X1 U3222 ( .A(n1500), .ZN(n3902) );
  AOI22_X1 U3223 ( .A1(DATAIN[11]), .A2(n3389), .B1(n3393), .B2(
        \registers[7][11] ), .ZN(n1500) );
  INV_X1 U3224 ( .A(n1501), .ZN(n3903) );
  AOI22_X1 U3225 ( .A1(n708), .A2(n3389), .B1(n3393), .B2(\registers[7][12] ), 
        .ZN(n1501) );
  INV_X1 U3226 ( .A(n1502), .ZN(n3904) );
  AOI22_X1 U3227 ( .A1(n706), .A2(n3389), .B1(n3393), .B2(\registers[7][13] ), 
        .ZN(n1502) );
  INV_X1 U3228 ( .A(n1503), .ZN(n3905) );
  AOI22_X1 U3229 ( .A1(n704), .A2(n3389), .B1(n3393), .B2(\registers[7][14] ), 
        .ZN(n1503) );
  INV_X1 U3230 ( .A(n1504), .ZN(n3906) );
  AOI22_X1 U3231 ( .A1(n702), .A2(n3389), .B1(n3394), .B2(\registers[7][15] ), 
        .ZN(n1504) );
  INV_X1 U3232 ( .A(n1505), .ZN(n3907) );
  AOI22_X1 U3233 ( .A1(n712), .A2(n358), .B1(n3394), .B2(\registers[7][16] ), 
        .ZN(n1505) );
  INV_X1 U3234 ( .A(n1506), .ZN(n3908) );
  AOI22_X1 U3235 ( .A1(n710), .A2(n3390), .B1(n3394), .B2(\registers[7][17] ), 
        .ZN(n1506) );
  INV_X1 U3236 ( .A(n1507), .ZN(n3909) );
  AOI22_X1 U3237 ( .A1(n700), .A2(n3390), .B1(n3394), .B2(\registers[7][18] ), 
        .ZN(n1507) );
  INV_X1 U3238 ( .A(n1508), .ZN(n3910) );
  AOI22_X1 U3239 ( .A1(n792), .A2(n3390), .B1(n3394), .B2(\registers[7][19] ), 
        .ZN(n1508) );
  INV_X1 U3240 ( .A(n1509), .ZN(n3911) );
  AOI22_X1 U3241 ( .A1(n876), .A2(n3390), .B1(n3395), .B2(\registers[7][20] ), 
        .ZN(n1509) );
  INV_X1 U3242 ( .A(n1510), .ZN(n3912) );
  AOI22_X1 U3243 ( .A1(n888), .A2(n358), .B1(n3395), .B2(\registers[7][21] ), 
        .ZN(n1510) );
  INV_X1 U3244 ( .A(n1511), .ZN(n3913) );
  AOI22_X1 U3245 ( .A1(n586), .A2(n3390), .B1(n3395), .B2(\registers[7][22] ), 
        .ZN(n1511) );
  INV_X1 U3246 ( .A(n1512), .ZN(n3914) );
  AOI22_X1 U3247 ( .A1(n887), .A2(n3390), .B1(n3395), .B2(\registers[7][23] ), 
        .ZN(n1512) );
  INV_X1 U3248 ( .A(n1513), .ZN(n3915) );
  AOI22_X1 U3249 ( .A1(n872), .A2(n3390), .B1(n3395), .B2(\registers[7][24] ), 
        .ZN(n1513) );
  INV_X1 U3250 ( .A(n1514), .ZN(n3916) );
  AOI22_X1 U3251 ( .A1(n886), .A2(n3390), .B1(n3396), .B2(\registers[7][25] ), 
        .ZN(n1514) );
  INV_X1 U3252 ( .A(n1515), .ZN(n3917) );
  AOI22_X1 U3253 ( .A1(n869), .A2(n358), .B1(n3396), .B2(\registers[7][26] ), 
        .ZN(n1515) );
  INV_X1 U3254 ( .A(n1516), .ZN(n3918) );
  AOI22_X1 U3255 ( .A1(n885), .A2(n358), .B1(n3396), .B2(\registers[7][27] ), 
        .ZN(n1516) );
  INV_X1 U3256 ( .A(n1517), .ZN(n3919) );
  AOI22_X1 U3257 ( .A1(n868), .A2(n3389), .B1(n3396), .B2(\registers[7][28] ), 
        .ZN(n1517) );
  INV_X1 U3258 ( .A(n1518), .ZN(n3920) );
  AOI22_X1 U3259 ( .A1(n883), .A2(n358), .B1(n3396), .B2(\registers[7][29] ), 
        .ZN(n1518) );
  INV_X1 U3260 ( .A(n1519), .ZN(n3921) );
  AOI22_X1 U3261 ( .A1(n190), .A2(n3390), .B1(n3397), .B2(\registers[7][30] ), 
        .ZN(n1519) );
  INV_X1 U3262 ( .A(n1520), .ZN(n3922) );
  AOI22_X1 U3263 ( .A1(n252), .A2(n358), .B1(n3397), .B2(\registers[7][31] ), 
        .ZN(n1520) );
  INV_X1 U3264 ( .A(n1531), .ZN(n3867) );
  AOI22_X1 U3265 ( .A1(n3382), .A2(n203), .B1(n3386), .B2(\registers[6][8] ), 
        .ZN(n1531) );
  INV_X1 U3266 ( .A(n1532), .ZN(n3868) );
  AOI22_X1 U3267 ( .A1(n3384), .A2(n879), .B1(n3386), .B2(\registers[6][9] ), 
        .ZN(n1532) );
  INV_X1 U3268 ( .A(n1533), .ZN(n3869) );
  AOI22_X1 U3269 ( .A1(n599), .A2(DATAIN[10]), .B1(n3385), .B2(
        \registers[6][10] ), .ZN(n1533) );
  INV_X1 U3270 ( .A(n1534), .ZN(n3870) );
  AOI22_X1 U3271 ( .A1(n598), .A2(DATAIN[11]), .B1(n3385), .B2(
        \registers[6][11] ), .ZN(n1534) );
  INV_X1 U3272 ( .A(n1535), .ZN(n3871) );
  AOI22_X1 U3273 ( .A1(n398), .A2(n708), .B1(n3385), .B2(\registers[6][12] ), 
        .ZN(n1535) );
  INV_X1 U3274 ( .A(n1536), .ZN(n3872) );
  AOI22_X1 U3275 ( .A1(n598), .A2(n706), .B1(n3386), .B2(\registers[6][13] ), 
        .ZN(n1536) );
  INV_X1 U3276 ( .A(n1537), .ZN(n3873) );
  AOI22_X1 U3277 ( .A1(n398), .A2(n704), .B1(n3386), .B2(\registers[6][14] ), 
        .ZN(n1537) );
  INV_X1 U3278 ( .A(n1538), .ZN(n3874) );
  AOI22_X1 U3279 ( .A1(n576), .A2(n702), .B1(n3388), .B2(\registers[6][15] ), 
        .ZN(n1538) );
  INV_X1 U3280 ( .A(n1539), .ZN(n3875) );
  AOI22_X1 U3281 ( .A1(n599), .A2(n712), .B1(n3388), .B2(\registers[6][16] ), 
        .ZN(n1539) );
  INV_X1 U3282 ( .A(n1540), .ZN(n3876) );
  AOI22_X1 U3283 ( .A1(n598), .A2(n710), .B1(n3385), .B2(\registers[6][17] ), 
        .ZN(n1540) );
  INV_X1 U3284 ( .A(n1541), .ZN(n3877) );
  AOI22_X1 U3285 ( .A1(n3384), .A2(n700), .B1(n3386), .B2(\registers[6][18] ), 
        .ZN(n1541) );
  INV_X1 U3286 ( .A(n1542), .ZN(n3878) );
  AOI22_X1 U3287 ( .A1(n792), .A2(n547), .B1(n3388), .B2(\registers[6][19] ), 
        .ZN(n1542) );
  INV_X1 U3288 ( .A(n1543), .ZN(n3879) );
  AOI22_X1 U3289 ( .A1(n876), .A2(n195), .B1(n3388), .B2(\registers[6][20] ), 
        .ZN(n1543) );
  INV_X1 U3290 ( .A(n1544), .ZN(n3880) );
  AOI22_X1 U3291 ( .A1(n576), .A2(n889), .B1(n3388), .B2(\registers[6][21] ), 
        .ZN(n1544) );
  INV_X1 U3292 ( .A(n1545), .ZN(n3881) );
  AOI22_X1 U3293 ( .A1(n195), .A2(n373), .B1(n3385), .B2(\registers[6][22] ), 
        .ZN(n1545) );
  INV_X1 U3294 ( .A(n1546), .ZN(n3882) );
  AOI22_X1 U3295 ( .A1(n3383), .A2(n371), .B1(n3386), .B2(\registers[6][23] ), 
        .ZN(n1546) );
  INV_X1 U3296 ( .A(n1547), .ZN(n3883) );
  AOI22_X1 U3297 ( .A1(n576), .A2(n236), .B1(n3386), .B2(\registers[6][24] ), 
        .ZN(n1547) );
  INV_X1 U3298 ( .A(n1548), .ZN(n3884) );
  AOI22_X1 U3299 ( .A1(n598), .A2(n367), .B1(n3388), .B2(\registers[6][25] ), 
        .ZN(n1548) );
  INV_X1 U3300 ( .A(n1549), .ZN(n3885) );
  AOI22_X1 U3301 ( .A1(n870), .A2(n3383), .B1(n3385), .B2(\registers[6][26] ), 
        .ZN(n1549) );
  INV_X1 U3302 ( .A(n1550), .ZN(n3886) );
  AOI22_X1 U3303 ( .A1(n547), .A2(n251), .B1(n3388), .B2(\registers[6][27] ), 
        .ZN(n1550) );
  INV_X1 U3304 ( .A(n1551), .ZN(n3887) );
  AOI22_X1 U3305 ( .A1(n576), .A2(n250), .B1(n3388), .B2(\registers[6][28] ), 
        .ZN(n1551) );
  INV_X1 U3306 ( .A(n1552), .ZN(n3888) );
  AOI22_X1 U3307 ( .A1(n3382), .A2(n883), .B1(n3388), .B2(\registers[6][29] ), 
        .ZN(n1552) );
  INV_X1 U3308 ( .A(n1553), .ZN(n3889) );
  AOI22_X1 U3309 ( .A1(n599), .A2(n866), .B1(n3385), .B2(\registers[6][30] ), 
        .ZN(n1553) );
  INV_X1 U3310 ( .A(n1554), .ZN(n3890) );
  AOI22_X1 U3311 ( .A1(n599), .A2(n252), .B1(n3386), .B2(\registers[6][31] ), 
        .ZN(n1554) );
  INV_X1 U3312 ( .A(n1431), .ZN(n3747) );
  AOI22_X1 U3313 ( .A1(n794), .A2(n382), .B1(n354), .B2(\registers[9][8] ), 
        .ZN(n1431) );
  INV_X1 U3314 ( .A(n1433), .ZN(n3748) );
  AOI22_X1 U3315 ( .A1(DATAIN[10]), .A2(n3408), .B1(n354), .B2(
        \registers[9][10] ), .ZN(n1433) );
  INV_X1 U3316 ( .A(n1434), .ZN(n3749) );
  AOI22_X1 U3317 ( .A1(DATAIN[11]), .A2(n3408), .B1(n3412), .B2(
        \registers[9][11] ), .ZN(n1434) );
  INV_X1 U3318 ( .A(n1435), .ZN(n3750) );
  AOI22_X1 U3319 ( .A1(n708), .A2(n384), .B1(n381), .B2(\registers[9][12] ), 
        .ZN(n1435) );
  INV_X1 U3320 ( .A(n1436), .ZN(n3751) );
  AOI22_X1 U3321 ( .A1(n706), .A2(n3408), .B1(n3410), .B2(\registers[9][13] ), 
        .ZN(n1436) );
  INV_X1 U3322 ( .A(n1437), .ZN(n3752) );
  AOI22_X1 U3323 ( .A1(n704), .A2(n561), .B1(n3411), .B2(\registers[9][14] ), 
        .ZN(n1437) );
  INV_X1 U3324 ( .A(n1438), .ZN(n3753) );
  AOI22_X1 U3325 ( .A1(n702), .A2(n3409), .B1(n3411), .B2(\registers[9][15] ), 
        .ZN(n1438) );
  INV_X1 U3326 ( .A(n1439), .ZN(n3754) );
  AOI22_X1 U3327 ( .A1(n712), .A2(n384), .B1(n3411), .B2(\registers[9][16] ), 
        .ZN(n1439) );
  INV_X1 U3328 ( .A(n1440), .ZN(n3755) );
  AOI22_X1 U3329 ( .A1(n710), .A2(n3408), .B1(n385), .B2(\registers[9][17] ), 
        .ZN(n1440) );
  INV_X1 U3330 ( .A(n1441), .ZN(n3756) );
  AOI22_X1 U3331 ( .A1(n382), .A2(n700), .B1(n385), .B2(\registers[9][18] ), 
        .ZN(n1441) );
  INV_X1 U3332 ( .A(n1442), .ZN(n3757) );
  AOI22_X1 U3333 ( .A1(n792), .A2(n382), .B1(n385), .B2(\registers[9][19] ), 
        .ZN(n1442) );
  INV_X1 U3334 ( .A(n1443), .ZN(n3758) );
  AOI22_X1 U3335 ( .A1(n876), .A2(n3409), .B1(n3412), .B2(\registers[9][20] ), 
        .ZN(n1443) );
  INV_X1 U3336 ( .A(n1444), .ZN(n3759) );
  AOI22_X1 U3337 ( .A1(n889), .A2(n3409), .B1(n381), .B2(\registers[9][21] ), 
        .ZN(n1444) );
  INV_X1 U3338 ( .A(n1446), .ZN(n3760) );
  AOI22_X1 U3339 ( .A1(n561), .A2(n887), .B1(n385), .B2(\registers[9][23] ), 
        .ZN(n1446) );
  INV_X1 U3340 ( .A(n1447), .ZN(n3761) );
  AOI22_X1 U3341 ( .A1(n3409), .A2(n872), .B1(n385), .B2(\registers[9][24] ), 
        .ZN(n1447) );
  INV_X1 U3342 ( .A(n1448), .ZN(n3762) );
  AOI22_X1 U3343 ( .A1(n561), .A2(n886), .B1(n385), .B2(\registers[9][25] ), 
        .ZN(n1448) );
  INV_X1 U3344 ( .A(n1449), .ZN(n3763) );
  AOI22_X1 U3345 ( .A1(n870), .A2(n384), .B1(n385), .B2(\registers[9][26] ), 
        .ZN(n1449) );
  INV_X1 U3346 ( .A(n1450), .ZN(n3764) );
  AOI22_X1 U3347 ( .A1(n885), .A2(n384), .B1(n3410), .B2(\registers[9][27] ), 
        .ZN(n1450) );
  INV_X1 U3348 ( .A(n1451), .ZN(n3765) );
  AOI22_X1 U3349 ( .A1(n382), .A2(n868), .B1(n385), .B2(\registers[9][28] ), 
        .ZN(n1451) );
  INV_X1 U3350 ( .A(n1452), .ZN(n3766) );
  AOI22_X1 U3351 ( .A1(n3409), .A2(n883), .B1(n385), .B2(\registers[9][29] ), 
        .ZN(n1452) );
  INV_X1 U3352 ( .A(n1453), .ZN(n3767) );
  AOI22_X1 U3353 ( .A1(n866), .A2(n561), .B1(n3410), .B2(\registers[9][30] ), 
        .ZN(n1453) );
  INV_X1 U3354 ( .A(n1454), .ZN(n3768) );
  AOI22_X1 U3355 ( .A1(n878), .A2(n382), .B1(n3411), .B2(\registers[9][31] ), 
        .ZN(n1454) );
  INV_X1 U3356 ( .A(n1568), .ZN(n3835) );
  AOI22_X1 U3357 ( .A1(n794), .A2(n365), .B1(n264), .B2(\registers[1][8] ), 
        .ZN(n1568) );
  INV_X1 U3358 ( .A(n1569), .ZN(n3836) );
  AOI22_X1 U3359 ( .A1(n589), .A2(n3337), .B1(n262), .B2(\registers[1][9] ), 
        .ZN(n1569) );
  INV_X1 U3360 ( .A(n1570), .ZN(n3837) );
  AOI22_X1 U3361 ( .A1(DATAIN[10]), .A2(n3337), .B1(n3340), .B2(
        \registers[1][10] ), .ZN(n1570) );
  INV_X1 U3362 ( .A(n1571), .ZN(n3838) );
  AOI22_X1 U3363 ( .A1(n365), .A2(DATAIN[11]), .B1(n3340), .B2(
        \registers[1][11] ), .ZN(n1571) );
  INV_X1 U3364 ( .A(n1572), .ZN(n3839) );
  AOI22_X1 U3365 ( .A1(n708), .A2(n380), .B1(n3340), .B2(\registers[1][12] ), 
        .ZN(n1572) );
  INV_X1 U3366 ( .A(n1573), .ZN(n3840) );
  AOI22_X1 U3367 ( .A1(n706), .A2(n380), .B1(n3340), .B2(\registers[1][13] ), 
        .ZN(n1573) );
  INV_X1 U3368 ( .A(n1574), .ZN(n3841) );
  AOI22_X1 U3369 ( .A1(n704), .A2(n3339), .B1(n3340), .B2(\registers[1][14] ), 
        .ZN(n1574) );
  INV_X1 U3370 ( .A(n1575), .ZN(n3842) );
  AOI22_X1 U3371 ( .A1(n702), .A2(n3337), .B1(n3340), .B2(\registers[1][15] ), 
        .ZN(n1575) );
  INV_X1 U3372 ( .A(n1576), .ZN(n3843) );
  AOI22_X1 U3373 ( .A1(n712), .A2(n3339), .B1(n3340), .B2(\registers[1][16] ), 
        .ZN(n1576) );
  INV_X1 U3374 ( .A(n1577), .ZN(n3844) );
  AOI22_X1 U3375 ( .A1(n710), .A2(n3339), .B1(n3340), .B2(\registers[1][17] ), 
        .ZN(n1577) );
  INV_X1 U3376 ( .A(n1578), .ZN(n3845) );
  AOI22_X1 U3377 ( .A1(n700), .A2(n365), .B1(n263), .B2(\registers[1][18] ), 
        .ZN(n1578) );
  INV_X1 U3378 ( .A(n1579), .ZN(n3846) );
  AOI22_X1 U3379 ( .A1(n792), .A2(n3337), .B1(n3340), .B2(\registers[1][19] ), 
        .ZN(n1579) );
  INV_X1 U3380 ( .A(n1580), .ZN(n3847) );
  AOI22_X1 U3381 ( .A1(n876), .A2(n366), .B1(n1), .B2(\registers[1][20] ), 
        .ZN(n1580) );
  INV_X1 U3382 ( .A(n1581), .ZN(n3848) );
  AOI22_X1 U3383 ( .A1(n889), .A2(n3339), .B1(n3340), .B2(\registers[1][21] ), 
        .ZN(n1581) );
  INV_X1 U3384 ( .A(n1582), .ZN(n3849) );
  AOI22_X1 U3385 ( .A1(n365), .A2(n373), .B1(n3340), .B2(\registers[1][22] ), 
        .ZN(n1582) );
  INV_X1 U3386 ( .A(n1583), .ZN(n3850) );
  AOI22_X1 U3387 ( .A1(n371), .A2(n366), .B1(n1), .B2(\registers[1][23] ), 
        .ZN(n1583) );
  INV_X1 U3388 ( .A(n1584), .ZN(n3851) );
  AOI22_X1 U3389 ( .A1(n236), .A2(n380), .B1(n3340), .B2(\registers[1][24] ), 
        .ZN(n1584) );
  INV_X1 U3390 ( .A(n1585), .ZN(n3852) );
  AOI22_X1 U3391 ( .A1(n367), .A2(n380), .B1(n264), .B2(\registers[1][25] ), 
        .ZN(n1585) );
  INV_X1 U3392 ( .A(n1586), .ZN(n3853) );
  AOI22_X1 U3393 ( .A1(n870), .A2(n3339), .B1(n3340), .B2(\registers[1][26] ), 
        .ZN(n1586) );
  INV_X1 U3394 ( .A(n1587), .ZN(n3854) );
  AOI22_X1 U3395 ( .A1(n251), .A2(n3338), .B1(n1), .B2(\registers[1][27] ), 
        .ZN(n1587) );
  INV_X1 U3396 ( .A(n1588), .ZN(n3855) );
  AOI22_X1 U3397 ( .A1(n250), .A2(n380), .B1(n3340), .B2(\registers[1][28] ), 
        .ZN(n1588) );
  INV_X1 U3398 ( .A(n1589), .ZN(n3856) );
  AOI22_X1 U3399 ( .A1(n883), .A2(n3338), .B1(n263), .B2(\registers[1][29] ), 
        .ZN(n1589) );
  INV_X1 U3400 ( .A(n1590), .ZN(n3857) );
  AOI22_X1 U3401 ( .A1(n288), .A2(n3337), .B1(n264), .B2(\registers[1][30] ), 
        .ZN(n1590) );
  INV_X1 U3402 ( .A(n1591), .ZN(n3858) );
  AOI22_X1 U3403 ( .A1(n878), .A2(n365), .B1(n263), .B2(\registers[1][31] ), 
        .ZN(n1591) );
  INV_X1 U3404 ( .A(n1292), .ZN(n3962) );
  AOI22_X1 U3405 ( .A1(n204), .A2(n546), .B1(n19), .B2(\registers[19][8] ), 
        .ZN(n1292) );
  INV_X1 U3406 ( .A(n1293), .ZN(n3963) );
  AOI22_X1 U3407 ( .A1(n879), .A2(n597), .B1(n19), .B2(\registers[19][9] ), 
        .ZN(n1293) );
  INV_X1 U3408 ( .A(n1294), .ZN(n3964) );
  AOI22_X1 U3409 ( .A1(DATAIN[10]), .A2(n396), .B1(n3), .B2(
        \registers[19][10] ), .ZN(n1294) );
  INV_X1 U3410 ( .A(n1295), .ZN(n3965) );
  AOI22_X1 U3411 ( .A1(n202), .A2(DATAIN[11]), .B1(n19), .B2(
        \registers[19][11] ), .ZN(n1295) );
  INV_X1 U3412 ( .A(n1296), .ZN(n3966) );
  AOI22_X1 U3413 ( .A1(n708), .A2(n546), .B1(n2), .B2(\registers[19][12] ), 
        .ZN(n1296) );
  INV_X1 U3414 ( .A(n1297), .ZN(n3967) );
  AOI22_X1 U3415 ( .A1(n706), .A2(n724), .B1(n163), .B2(\registers[19][13] ), 
        .ZN(n1297) );
  INV_X1 U3416 ( .A(n1298), .ZN(n3968) );
  AOI22_X1 U3417 ( .A1(n704), .A2(n724), .B1(n2), .B2(\registers[19][14] ), 
        .ZN(n1298) );
  INV_X1 U3418 ( .A(n1299), .ZN(n3969) );
  AOI22_X1 U3419 ( .A1(n702), .A2(n3487), .B1(n163), .B2(\registers[19][15] ), 
        .ZN(n1299) );
  INV_X1 U3420 ( .A(n1300), .ZN(n3970) );
  AOI22_X1 U3421 ( .A1(n712), .A2(n725), .B1(n161), .B2(\registers[19][16] ), 
        .ZN(n1300) );
  INV_X1 U3422 ( .A(n1301), .ZN(n3971) );
  AOI22_X1 U3423 ( .A1(n710), .A2(n725), .B1(n4), .B2(\registers[19][17] ), 
        .ZN(n1301) );
  INV_X1 U3424 ( .A(n1302), .ZN(n3972) );
  AOI22_X1 U3425 ( .A1(n700), .A2(n724), .B1(n162), .B2(\registers[19][18] ), 
        .ZN(n1302) );
  INV_X1 U3426 ( .A(n1303), .ZN(n3973) );
  AOI22_X1 U3427 ( .A1(n792), .A2(n3486), .B1(n3), .B2(\registers[19][19] ), 
        .ZN(n1303) );
  INV_X1 U3428 ( .A(n1304), .ZN(n3974) );
  AOI22_X1 U3429 ( .A1(n876), .A2(n765), .B1(n162), .B2(\registers[19][20] ), 
        .ZN(n1304) );
  INV_X1 U3430 ( .A(n1305), .ZN(n3975) );
  AOI22_X1 U3431 ( .A1(n889), .A2(n765), .B1(n163), .B2(\registers[19][21] ), 
        .ZN(n1305) );
  INV_X1 U3432 ( .A(n1306), .ZN(n3976) );
  AOI22_X1 U3433 ( .A1(n373), .A2(n3485), .B1(n162), .B2(\registers[19][22] ), 
        .ZN(n1306) );
  INV_X1 U3434 ( .A(n1307), .ZN(n3977) );
  AOI22_X1 U3435 ( .A1(n887), .A2(n597), .B1(n163), .B2(\registers[19][23] ), 
        .ZN(n1307) );
  INV_X1 U3436 ( .A(n1308), .ZN(n3978) );
  AOI22_X1 U3437 ( .A1(n872), .A2(n396), .B1(n162), .B2(\registers[19][24] ), 
        .ZN(n1308) );
  INV_X1 U3438 ( .A(n1309), .ZN(n3979) );
  AOI22_X1 U3439 ( .A1(n367), .A2(n202), .B1(n161), .B2(\registers[19][25] ), 
        .ZN(n1309) );
  INV_X1 U3440 ( .A(n1310), .ZN(n3980) );
  AOI22_X1 U3441 ( .A1(n870), .A2(n546), .B1(n2), .B2(\registers[19][26] ), 
        .ZN(n1310) );
  INV_X1 U3442 ( .A(n1311), .ZN(n3981) );
  AOI22_X1 U3443 ( .A1(n885), .A2(n3486), .B1(n161), .B2(\registers[19][27] ), 
        .ZN(n1311) );
  INV_X1 U3444 ( .A(n1312), .ZN(n3982) );
  AOI22_X1 U3445 ( .A1(n868), .A2(n3487), .B1(n2), .B2(\registers[19][28] ), 
        .ZN(n1312) );
  INV_X1 U3446 ( .A(n1313), .ZN(n3983) );
  AOI22_X1 U3447 ( .A1(n397), .A2(n597), .B1(n161), .B2(\registers[19][29] ), 
        .ZN(n1313) );
  INV_X1 U3448 ( .A(n1314), .ZN(n3984) );
  AOI22_X1 U3449 ( .A1(n190), .A2(n3485), .B1(n3491), .B2(\registers[19][30] ), 
        .ZN(n1314) );
  INV_X1 U3450 ( .A(n1315), .ZN(n3985) );
  AOI22_X1 U3451 ( .A1(n252), .A2(n724), .B1(n3491), .B2(\registers[19][31] ), 
        .ZN(n1315) );
  INV_X1 U3452 ( .A(n1325), .ZN(n3931) );
  AOI22_X1 U3453 ( .A1(n729), .A2(n203), .B1(n3481), .B2(\registers[18][8] ), 
        .ZN(n1325) );
  INV_X1 U3454 ( .A(n1326), .ZN(n3932) );
  AOI22_X1 U3455 ( .A1(n3478), .A2(n879), .B1(n3481), .B2(\registers[18][9] ), 
        .ZN(n1326) );
  INV_X1 U3456 ( .A(n1327), .ZN(n3933) );
  AOI22_X1 U3457 ( .A1(DATAIN[10]), .A2(n596), .B1(n3480), .B2(
        \registers[18][10] ), .ZN(n1327) );
  INV_X1 U3458 ( .A(n1328), .ZN(n3934) );
  AOI22_X1 U3459 ( .A1(n3479), .A2(DATAIN[11]), .B1(n3481), .B2(
        \registers[18][11] ), .ZN(n1328) );
  INV_X1 U3460 ( .A(n1329), .ZN(n3935) );
  AOI22_X1 U3461 ( .A1(n708), .A2(n596), .B1(n3480), .B2(\registers[18][12] ), 
        .ZN(n1329) );
  INV_X1 U3462 ( .A(n1330), .ZN(n3936) );
  AOI22_X1 U3463 ( .A1(n706), .A2(n596), .B1(n3482), .B2(\registers[18][13] ), 
        .ZN(n1330) );
  INV_X1 U3464 ( .A(n1331), .ZN(n3937) );
  AOI22_X1 U3465 ( .A1(n704), .A2(n3478), .B1(n3483), .B2(\registers[18][14] ), 
        .ZN(n1331) );
  INV_X1 U3466 ( .A(n1332), .ZN(n3938) );
  AOI22_X1 U3467 ( .A1(n702), .A2(n764), .B1(n3482), .B2(\registers[18][15] ), 
        .ZN(n1332) );
  INV_X1 U3468 ( .A(n1333), .ZN(n3939) );
  AOI22_X1 U3469 ( .A1(n712), .A2(n763), .B1(n3483), .B2(\registers[18][16] ), 
        .ZN(n1333) );
  INV_X1 U3470 ( .A(n1334), .ZN(n3940) );
  AOI22_X1 U3471 ( .A1(n710), .A2(n3478), .B1(n3480), .B2(\registers[18][17] ), 
        .ZN(n1334) );
  INV_X1 U3472 ( .A(n1335), .ZN(n3941) );
  AOI22_X1 U3473 ( .A1(n700), .A2(n764), .B1(n3482), .B2(\registers[18][18] ), 
        .ZN(n1335) );
  INV_X1 U3474 ( .A(n1336), .ZN(n3942) );
  AOI22_X1 U3475 ( .A1(n792), .A2(n763), .B1(n3480), .B2(\registers[18][19] ), 
        .ZN(n1336) );
  INV_X1 U3476 ( .A(n1337), .ZN(n3943) );
  AOI22_X1 U3477 ( .A1(n876), .A2(n730), .B1(n3482), .B2(\registers[18][20] ), 
        .ZN(n1337) );
  INV_X1 U3478 ( .A(n1338), .ZN(n3944) );
  AOI22_X1 U3479 ( .A1(n888), .A2(n764), .B1(n3482), .B2(\registers[18][21] ), 
        .ZN(n1338) );
  INV_X1 U3480 ( .A(n1339), .ZN(n3945) );
  AOI22_X1 U3481 ( .A1(n586), .A2(n3477), .B1(n3482), .B2(\registers[18][22] ), 
        .ZN(n1339) );
  INV_X1 U3482 ( .A(n1340), .ZN(n3946) );
  AOI22_X1 U3483 ( .A1(n371), .A2(n3477), .B1(n3482), .B2(\registers[18][23] ), 
        .ZN(n1340) );
  INV_X1 U3484 ( .A(n1341), .ZN(n3947) );
  AOI22_X1 U3485 ( .A1(n236), .A2(n3477), .B1(n3482), .B2(\registers[18][24] ), 
        .ZN(n1341) );
  INV_X1 U3486 ( .A(n1342), .ZN(n3948) );
  AOI22_X1 U3487 ( .A1(n886), .A2(n3478), .B1(n3483), .B2(\registers[18][25] ), 
        .ZN(n1342) );
  INV_X1 U3488 ( .A(n1343), .ZN(n3949) );
  AOI22_X1 U3489 ( .A1(n870), .A2(n730), .B1(n3483), .B2(\registers[18][26] ), 
        .ZN(n1343) );
  INV_X1 U3490 ( .A(n1344), .ZN(n3950) );
  AOI22_X1 U3491 ( .A1(n764), .A2(n251), .B1(n3483), .B2(\registers[18][27] ), 
        .ZN(n1344) );
  INV_X1 U3492 ( .A(n1345), .ZN(n3951) );
  AOI22_X1 U3493 ( .A1(n729), .A2(n250), .B1(n3483), .B2(\registers[18][28] ), 
        .ZN(n1345) );
  INV_X1 U3494 ( .A(n1346), .ZN(n3952) );
  AOI22_X1 U3495 ( .A1(n730), .A2(n397), .B1(n3483), .B2(\registers[18][29] ), 
        .ZN(n1346) );
  INV_X1 U3496 ( .A(n1347), .ZN(n3953) );
  AOI22_X1 U3497 ( .A1(n3479), .A2(n866), .B1(n3484), .B2(\registers[18][30] ), 
        .ZN(n1347) );
  INV_X1 U3498 ( .A(n1348), .ZN(n3954) );
  AOI22_X1 U3499 ( .A1(n729), .A2(n878), .B1(n3484), .B2(\registers[18][31] ), 
        .ZN(n1348) );
  INV_X1 U3500 ( .A(n1179), .ZN(n4043) );
  AOI22_X1 U3501 ( .A1(DATAIN[0]), .A2(n17), .B1(n3530), .B2(
        \registers[24][0] ), .ZN(n1179) );
  INV_X1 U3502 ( .A(n1181), .ZN(n4044) );
  AOI22_X1 U3503 ( .A1(n892), .A2(n604), .B1(n3531), .B2(\registers[24][1] ), 
        .ZN(n1181) );
  INV_X1 U3504 ( .A(n1182), .ZN(n4045) );
  AOI22_X1 U3505 ( .A1(n890), .A2(n604), .B1(n3529), .B2(\registers[24][2] ), 
        .ZN(n1182) );
  INV_X1 U3506 ( .A(n1455), .ZN(n3711) );
  AOI22_X1 U3507 ( .A1(n180), .A2(n675), .B1(n23), .B2(\registers[8][0] ), 
        .ZN(n1455) );
  INV_X1 U3508 ( .A(n1457), .ZN(n3712) );
  AOI22_X1 U3509 ( .A1(n892), .A2(n675), .B1(n3404), .B2(\registers[8][1] ), 
        .ZN(n1457) );
  INV_X1 U3510 ( .A(n1458), .ZN(n3713) );
  AOI22_X1 U3511 ( .A1(n375), .A2(n3398), .B1(n3406), .B2(\registers[8][2] ), 
        .ZN(n1458) );
  INV_X1 U3512 ( .A(n1190), .ZN(n4053) );
  AOI22_X1 U3513 ( .A1(DATAIN[10]), .A2(n3524), .B1(n3527), .B2(
        \registers[24][10] ), .ZN(n1190) );
  INV_X1 U3514 ( .A(n1191), .ZN(n4054) );
  AOI22_X1 U3515 ( .A1(DATAIN[11]), .A2(n3525), .B1(n557), .B2(
        \registers[24][11] ), .ZN(n1191) );
  INV_X1 U3516 ( .A(n1192), .ZN(n4055) );
  AOI22_X1 U3517 ( .A1(n788), .A2(n3525), .B1(n3527), .B2(\registers[24][12] ), 
        .ZN(n1192) );
  INV_X1 U3518 ( .A(n1193), .ZN(n4056) );
  AOI22_X1 U3519 ( .A1(n705), .A2(n17), .B1(n557), .B2(\registers[24][13] ), 
        .ZN(n1193) );
  INV_X1 U3520 ( .A(n1194), .ZN(n4057) );
  AOI22_X1 U3521 ( .A1(n783), .A2(n604), .B1(n3530), .B2(\registers[24][14] ), 
        .ZN(n1194) );
  INV_X1 U3522 ( .A(n1195), .ZN(n4058) );
  AOI22_X1 U3523 ( .A1(n780), .A2(n17), .B1(n3531), .B2(\registers[24][15] ), 
        .ZN(n1195) );
  INV_X1 U3524 ( .A(n1196), .ZN(n4059) );
  AOI22_X1 U3525 ( .A1(n712), .A2(n3526), .B1(n3529), .B2(\registers[24][16] ), 
        .ZN(n1196) );
  INV_X1 U3526 ( .A(n1197), .ZN(n4060) );
  AOI22_X1 U3527 ( .A1(n774), .A2(n3525), .B1(n3531), .B2(\registers[24][17] ), 
        .ZN(n1197) );
  INV_X1 U3528 ( .A(n1198), .ZN(n4061) );
  AOI22_X1 U3529 ( .A1(n771), .A2(n17), .B1(n3529), .B2(\registers[24][18] ), 
        .ZN(n1198) );
  INV_X1 U3530 ( .A(n1199), .ZN(n4062) );
  AOI22_X1 U3531 ( .A1(n792), .A2(n3526), .B1(n3528), .B2(\registers[24][19] ), 
        .ZN(n1199) );
  INV_X1 U3532 ( .A(n1200), .ZN(n4063) );
  AOI22_X1 U3533 ( .A1(n876), .A2(n604), .B1(n3528), .B2(\registers[24][20] ), 
        .ZN(n1200) );
  INV_X1 U3534 ( .A(n1201), .ZN(n4064) );
  AOI22_X1 U3535 ( .A1(n889), .A2(n603), .B1(n3527), .B2(\registers[24][21] ), 
        .ZN(n1201) );
  INV_X1 U3536 ( .A(n1202), .ZN(n4065) );
  AOI22_X1 U3537 ( .A1(n588), .A2(n603), .B1(n3529), .B2(\registers[24][22] ), 
        .ZN(n1202) );
  INV_X1 U3538 ( .A(n1203), .ZN(n4066) );
  AOI22_X1 U3539 ( .A1(n371), .A2(n3524), .B1(n3528), .B2(\registers[24][23] ), 
        .ZN(n1203) );
  INV_X1 U3540 ( .A(n1204), .ZN(n4067) );
  AOI22_X1 U3541 ( .A1(n236), .A2(n604), .B1(n557), .B2(\registers[24][24] ), 
        .ZN(n1204) );
  INV_X1 U3542 ( .A(n1205), .ZN(n4068) );
  AOI22_X1 U3543 ( .A1(n886), .A2(n603), .B1(n3527), .B2(\registers[24][25] ), 
        .ZN(n1205) );
  INV_X1 U3544 ( .A(n1206), .ZN(n4069) );
  AOI22_X1 U3545 ( .A1(n870), .A2(n3524), .B1(n3531), .B2(\registers[24][26] ), 
        .ZN(n1206) );
  INV_X1 U3546 ( .A(n1207), .ZN(n4070) );
  AOI22_X1 U3547 ( .A1(n251), .A2(n604), .B1(n3531), .B2(\registers[24][27] ), 
        .ZN(n1207) );
  INV_X1 U3548 ( .A(n1208), .ZN(n4071) );
  AOI22_X1 U3549 ( .A1(n250), .A2(n17), .B1(n3530), .B2(\registers[24][28] ), 
        .ZN(n1208) );
  INV_X1 U3550 ( .A(n1209), .ZN(n4072) );
  AOI22_X1 U3551 ( .A1(n883), .A2(n3525), .B1(n557), .B2(\registers[24][29] ), 
        .ZN(n1209) );
  INV_X1 U3552 ( .A(n1210), .ZN(n4073) );
  AOI22_X1 U3553 ( .A1(n288), .A2(n3524), .B1(n3528), .B2(\registers[24][30] ), 
        .ZN(n1210) );
  INV_X1 U3554 ( .A(n1466), .ZN(n3721) );
  AOI22_X1 U3555 ( .A1(DATAIN[10]), .A2(n3399), .B1(n3404), .B2(
        \registers[8][10] ), .ZN(n1466) );
  INV_X1 U3556 ( .A(n1467), .ZN(n3722) );
  AOI22_X1 U3557 ( .A1(DATAIN[11]), .A2(n676), .B1(n3406), .B2(
        \registers[8][11] ), .ZN(n1467) );
  INV_X1 U3558 ( .A(n1468), .ZN(n3723) );
  AOI22_X1 U3559 ( .A1(n788), .A2(n675), .B1(n3401), .B2(\registers[8][12] ), 
        .ZN(n1468) );
  INV_X1 U3560 ( .A(n1469), .ZN(n3724) );
  AOI22_X1 U3561 ( .A1(n705), .A2(n3398), .B1(n3403), .B2(\registers[8][13] ), 
        .ZN(n1469) );
  INV_X1 U3562 ( .A(n1470), .ZN(n3725) );
  AOI22_X1 U3563 ( .A1(n783), .A2(n3399), .B1(n23), .B2(\registers[8][14] ), 
        .ZN(n1470) );
  INV_X1 U3564 ( .A(n1471), .ZN(n3726) );
  AOI22_X1 U3565 ( .A1(n780), .A2(n3400), .B1(n3404), .B2(\registers[8][15] ), 
        .ZN(n1471) );
  INV_X1 U3566 ( .A(n1472), .ZN(n3727) );
  AOI22_X1 U3567 ( .A1(n777), .A2(n675), .B1(n3406), .B2(\registers[8][16] ), 
        .ZN(n1472) );
  INV_X1 U3568 ( .A(n1473), .ZN(n3728) );
  AOI22_X1 U3569 ( .A1(n206), .A2(n675), .B1(n3401), .B2(\registers[8][17] ), 
        .ZN(n1473) );
  INV_X1 U3570 ( .A(n1474), .ZN(n3729) );
  AOI22_X1 U3571 ( .A1(n771), .A2(n3400), .B1(n3403), .B2(\registers[8][18] ), 
        .ZN(n1474) );
  INV_X1 U3572 ( .A(n1475), .ZN(n3730) );
  AOI22_X1 U3573 ( .A1(n792), .A2(n760), .B1(n23), .B2(\registers[8][19] ), 
        .ZN(n1475) );
  INV_X1 U3574 ( .A(n1476), .ZN(n3731) );
  AOI22_X1 U3575 ( .A1(n876), .A2(n676), .B1(n189), .B2(\registers[8][20] ), 
        .ZN(n1476) );
  INV_X1 U3576 ( .A(n1477), .ZN(n3732) );
  AOI22_X1 U3577 ( .A1(n889), .A2(n676), .B1(n3405), .B2(\registers[8][21] ), 
        .ZN(n1477) );
  INV_X1 U3578 ( .A(n1478), .ZN(n3733) );
  AOI22_X1 U3579 ( .A1(n587), .A2(n760), .B1(n3405), .B2(\registers[8][22] ), 
        .ZN(n1478) );
  INV_X1 U3580 ( .A(n1479), .ZN(n3734) );
  AOI22_X1 U3581 ( .A1(n887), .A2(n676), .B1(n3405), .B2(\registers[8][23] ), 
        .ZN(n1479) );
  INV_X1 U3582 ( .A(n1480), .ZN(n3735) );
  AOI22_X1 U3583 ( .A1(n872), .A2(n3399), .B1(n3405), .B2(\registers[8][24] ), 
        .ZN(n1480) );
  INV_X1 U3584 ( .A(n1481), .ZN(n3736) );
  AOI22_X1 U3585 ( .A1(n367), .A2(n676), .B1(n3404), .B2(\registers[8][25] ), 
        .ZN(n1481) );
  INV_X1 U3586 ( .A(n1482), .ZN(n3737) );
  AOI22_X1 U3587 ( .A1(n870), .A2(n3398), .B1(n3406), .B2(\registers[8][26] ), 
        .ZN(n1482) );
  INV_X1 U3588 ( .A(n1483), .ZN(n3738) );
  AOI22_X1 U3589 ( .A1(n885), .A2(n760), .B1(n3401), .B2(\registers[8][27] ), 
        .ZN(n1483) );
  INV_X1 U3590 ( .A(n1484), .ZN(n3739) );
  AOI22_X1 U3591 ( .A1(n868), .A2(n760), .B1(n3403), .B2(\registers[8][28] ), 
        .ZN(n1484) );
  INV_X1 U3592 ( .A(n1485), .ZN(n3740) );
  AOI22_X1 U3593 ( .A1(n397), .A2(n3400), .B1(n23), .B2(\registers[8][29] ), 
        .ZN(n1485) );
  INV_X1 U3594 ( .A(n1486), .ZN(n3741) );
  AOI22_X1 U3595 ( .A1(n190), .A2(n3399), .B1(n189), .B2(\registers[8][30] ), 
        .ZN(n1486) );
  INV_X1 U3596 ( .A(n1459), .ZN(n3714) );
  AOI22_X1 U3597 ( .A1(n800), .A2(n3400), .B1(n3401), .B2(\registers[8][3] ), 
        .ZN(n1459) );
  INV_X1 U3598 ( .A(n1460), .ZN(n3715) );
  AOI22_X1 U3599 ( .A1(n882), .A2(n3399), .B1(n3403), .B2(\registers[8][4] ), 
        .ZN(n1460) );
  INV_X1 U3600 ( .A(n1461), .ZN(n3716) );
  AOI22_X1 U3601 ( .A1(n798), .A2(n676), .B1(n189), .B2(\registers[8][5] ), 
        .ZN(n1461) );
  INV_X1 U3602 ( .A(n1462), .ZN(n3717) );
  AOI22_X1 U3603 ( .A1(n227), .A2(n3398), .B1(n3402), .B2(\registers[8][6] ), 
        .ZN(n1462) );
  INV_X1 U3604 ( .A(n1463), .ZN(n3718) );
  AOI22_X1 U3605 ( .A1(n198), .A2(n3400), .B1(n3402), .B2(\registers[8][7] ), 
        .ZN(n1463) );
  INV_X1 U3606 ( .A(n1464), .ZN(n3719) );
  AOI22_X1 U3607 ( .A1(n203), .A2(n3398), .B1(n3402), .B2(\registers[8][8] ), 
        .ZN(n1464) );
  INV_X1 U3608 ( .A(n1465), .ZN(n3720) );
  AOI22_X1 U3609 ( .A1(n879), .A2(n675), .B1(n3402), .B2(\registers[8][9] ), 
        .ZN(n1465) );
  INV_X1 U3610 ( .A(n1487), .ZN(n3742) );
  AOI22_X1 U3611 ( .A1(n252), .A2(n760), .B1(n189), .B2(\registers[8][31] ), 
        .ZN(n1487) );
  INV_X1 U3612 ( .A(n1183), .ZN(n4046) );
  AOI22_X1 U3613 ( .A1(n800), .A2(n3526), .B1(n3529), .B2(\registers[24][3] ), 
        .ZN(n1183) );
  INV_X1 U3614 ( .A(n1184), .ZN(n4047) );
  AOI22_X1 U3615 ( .A1(n590), .A2(n3526), .B1(n3527), .B2(\registers[24][4] ), 
        .ZN(n1184) );
  INV_X1 U3616 ( .A(n1185), .ZN(n4048) );
  AOI22_X1 U3617 ( .A1(n798), .A2(n603), .B1(n3530), .B2(\registers[24][5] ), 
        .ZN(n1185) );
  INV_X1 U3618 ( .A(n1186), .ZN(n4049) );
  AOI22_X1 U3619 ( .A1(n228), .A2(n3524), .B1(n3527), .B2(\registers[24][6] ), 
        .ZN(n1186) );
  INV_X1 U3620 ( .A(n1187), .ZN(n4050) );
  AOI22_X1 U3621 ( .A1(n796), .A2(n3525), .B1(n3528), .B2(\registers[24][7] ), 
        .ZN(n1187) );
  INV_X1 U3622 ( .A(n1188), .ZN(n4051) );
  AOI22_X1 U3623 ( .A1(n794), .A2(n3526), .B1(n3527), .B2(\registers[24][8] ), 
        .ZN(n1188) );
  INV_X1 U3624 ( .A(n1189), .ZN(n4052) );
  AOI22_X1 U3625 ( .A1(n879), .A2(n17), .B1(n3530), .B2(\registers[24][9] ), 
        .ZN(n1189) );
  INV_X1 U3626 ( .A(n1211), .ZN(n4074) );
  AOI22_X1 U3627 ( .A1(n878), .A2(n603), .B1(n3527), .B2(\registers[24][31] ), 
        .ZN(n1211) );
  AND2_X1 U3628 ( .A1(RD2), .A2(ENABLE), .ZN(N218) );
  AND2_X1 U3629 ( .A1(RD1), .A2(ENABLE), .ZN(N83) );
  INV_X1 U3630 ( .A(n164), .ZN(n3345) );
  INV_X1 U3631 ( .A(n20), .ZN(n3355) );
  INV_X1 U3632 ( .A(n3371), .ZN(n3364) );
  INV_X1 U3633 ( .A(n3381), .ZN(n3374) );
  INV_X1 U3634 ( .A(n3387), .ZN(n3384) );
  INV_X1 U3635 ( .A(n3407), .ZN(n3400) );
  INV_X1 U3636 ( .A(n3422), .ZN(n3415) );
  INV_X1 U3637 ( .A(n3432), .ZN(n3425) );
  INV_X1 U3638 ( .A(n3458), .ZN(n3451) );
  INV_X1 U3639 ( .A(n3467), .ZN(n3460) );
  INV_X1 U3640 ( .A(n3471), .ZN(n3469) );
  INV_X1 U3641 ( .A(n3484), .ZN(n3479) );
  INV_X1 U3642 ( .A(n3491), .ZN(n3487) );
  INV_X1 U3643 ( .A(n3501), .ZN(n3494) );
  INV_X1 U3644 ( .A(n3511), .ZN(n3504) );
  INV_X1 U3645 ( .A(n3547), .ZN(n3540) );
  INV_X1 U3646 ( .A(n3557), .ZN(n3550) );
  INV_X1 U3647 ( .A(n3578), .ZN(n3575) );
  CLKBUF_X1 U3648 ( .A(N218), .Z(n3585) );
  CLKBUF_X1 U3649 ( .A(N218), .Z(n3586) );
  CLKBUF_X1 U3650 ( .A(N218), .Z(n3587) );
  CLKBUF_X1 U3651 ( .A(N218), .Z(n3588) );
  CLKBUF_X1 U3652 ( .A(N83), .Z(n3589) );
  CLKBUF_X1 U3653 ( .A(N83), .Z(n3590) );
  CLKBUF_X1 U3654 ( .A(N83), .Z(n3591) );
  CLKBUF_X1 U3655 ( .A(N83), .Z(n3592) );
  CLKBUF_X1 U3656 ( .A(n3710), .Z(n3604) );
  CLKBUF_X1 U3657 ( .A(n3709), .Z(n3605) );
  CLKBUF_X1 U3658 ( .A(n3709), .Z(n3606) );
  CLKBUF_X1 U3659 ( .A(n3709), .Z(n3607) );
  CLKBUF_X1 U3660 ( .A(n3709), .Z(n3608) );
  CLKBUF_X1 U3661 ( .A(n3709), .Z(n3609) );
  CLKBUF_X1 U3662 ( .A(n3709), .Z(n3610) );
  CLKBUF_X1 U3663 ( .A(n3708), .Z(n3611) );
  CLKBUF_X1 U3664 ( .A(n3708), .Z(n3612) );
  CLKBUF_X1 U3665 ( .A(n3708), .Z(n3613) );
  CLKBUF_X1 U3666 ( .A(n3708), .Z(n3614) );
  CLKBUF_X1 U3667 ( .A(n3708), .Z(n3615) );
  CLKBUF_X1 U3668 ( .A(n3708), .Z(n3616) );
  CLKBUF_X1 U3669 ( .A(n3707), .Z(n3617) );
  CLKBUF_X1 U3670 ( .A(n3707), .Z(n3618) );
  CLKBUF_X1 U3671 ( .A(n3707), .Z(n3619) );
  CLKBUF_X1 U3672 ( .A(n3707), .Z(n3620) );
  CLKBUF_X1 U3673 ( .A(n3707), .Z(n3621) );
  CLKBUF_X1 U3674 ( .A(n3707), .Z(n3622) );
  CLKBUF_X1 U3675 ( .A(n3706), .Z(n3623) );
  CLKBUF_X1 U3676 ( .A(n3706), .Z(n3624) );
  CLKBUF_X1 U3677 ( .A(n3706), .Z(n3625) );
  CLKBUF_X1 U3678 ( .A(n3706), .Z(n3626) );
  CLKBUF_X1 U3679 ( .A(n3706), .Z(n3627) );
  CLKBUF_X1 U3680 ( .A(n3706), .Z(n3628) );
  CLKBUF_X1 U3681 ( .A(n3705), .Z(n3629) );
  CLKBUF_X1 U3682 ( .A(n3705), .Z(n3630) );
  CLKBUF_X1 U3683 ( .A(n3705), .Z(n3631) );
  CLKBUF_X1 U3684 ( .A(n3705), .Z(n3632) );
  CLKBUF_X1 U3685 ( .A(n3705), .Z(n3633) );
  CLKBUF_X1 U3686 ( .A(n3705), .Z(n3634) );
  CLKBUF_X1 U3687 ( .A(n3704), .Z(n3635) );
  CLKBUF_X1 U3688 ( .A(n3704), .Z(n3636) );
  CLKBUF_X1 U3689 ( .A(n3704), .Z(n3637) );
  CLKBUF_X1 U3690 ( .A(n3704), .Z(n3638) );
  CLKBUF_X1 U3691 ( .A(n3704), .Z(n3639) );
  CLKBUF_X1 U3692 ( .A(n3704), .Z(n3640) );
  CLKBUF_X1 U3693 ( .A(n3703), .Z(n3641) );
  CLKBUF_X1 U3694 ( .A(n3703), .Z(n3642) );
  CLKBUF_X1 U3695 ( .A(n3703), .Z(n3643) );
  CLKBUF_X1 U3696 ( .A(n3703), .Z(n3644) );
  CLKBUF_X1 U3697 ( .A(n3703), .Z(n3645) );
  CLKBUF_X1 U3698 ( .A(n3703), .Z(n3646) );
  CLKBUF_X1 U3699 ( .A(n3702), .Z(n3647) );
  CLKBUF_X1 U3700 ( .A(n3702), .Z(n3648) );
  CLKBUF_X1 U3701 ( .A(n3702), .Z(n3649) );
  CLKBUF_X1 U3702 ( .A(n3702), .Z(n3650) );
  CLKBUF_X1 U3703 ( .A(n3702), .Z(n3651) );
  CLKBUF_X1 U3704 ( .A(n3702), .Z(n3652) );
  CLKBUF_X1 U3705 ( .A(n3701), .Z(n3653) );
  CLKBUF_X1 U3706 ( .A(n3701), .Z(n3654) );
  CLKBUF_X1 U3707 ( .A(n3701), .Z(n3655) );
  CLKBUF_X1 U3708 ( .A(n3701), .Z(n3656) );
  CLKBUF_X1 U3709 ( .A(n3701), .Z(n3657) );
  CLKBUF_X1 U3710 ( .A(n3701), .Z(n3658) );
  CLKBUF_X1 U3711 ( .A(n3700), .Z(n3659) );
  CLKBUF_X1 U3712 ( .A(n3700), .Z(n3660) );
  CLKBUF_X1 U3713 ( .A(n3700), .Z(n3661) );
  CLKBUF_X1 U3714 ( .A(n3700), .Z(n3662) );
  CLKBUF_X1 U3715 ( .A(n3700), .Z(n3663) );
  CLKBUF_X1 U3716 ( .A(n3700), .Z(n3664) );
  CLKBUF_X1 U3717 ( .A(n3699), .Z(n3665) );
  CLKBUF_X1 U3718 ( .A(n3699), .Z(n3666) );
  CLKBUF_X1 U3719 ( .A(n3699), .Z(n3667) );
  CLKBUF_X1 U3720 ( .A(n3699), .Z(n3668) );
  CLKBUF_X1 U3721 ( .A(n3699), .Z(n3669) );
  CLKBUF_X1 U3722 ( .A(n3699), .Z(n3670) );
  CLKBUF_X1 U3723 ( .A(n3698), .Z(n3671) );
  CLKBUF_X1 U3724 ( .A(n3698), .Z(n3672) );
  CLKBUF_X1 U3725 ( .A(n3698), .Z(n3673) );
  CLKBUF_X1 U3726 ( .A(n3698), .Z(n3674) );
  CLKBUF_X1 U3727 ( .A(n3698), .Z(n3675) );
  CLKBUF_X1 U3728 ( .A(n3698), .Z(n3676) );
  CLKBUF_X1 U3729 ( .A(n3697), .Z(n3677) );
  CLKBUF_X1 U3730 ( .A(n3697), .Z(n3678) );
  CLKBUF_X1 U3731 ( .A(n3697), .Z(n3679) );
  CLKBUF_X1 U3732 ( .A(n3697), .Z(n3680) );
  CLKBUF_X1 U3733 ( .A(n3697), .Z(n3681) );
  CLKBUF_X1 U3734 ( .A(n3697), .Z(n3682) );
  CLKBUF_X1 U3735 ( .A(n3696), .Z(n3683) );
  CLKBUF_X1 U3736 ( .A(n3696), .Z(n3684) );
  CLKBUF_X1 U3737 ( .A(n3696), .Z(n3685) );
  CLKBUF_X1 U3738 ( .A(n3696), .Z(n3686) );
  CLKBUF_X1 U3739 ( .A(n3696), .Z(n3687) );
  CLKBUF_X1 U3740 ( .A(n3696), .Z(n3688) );
  CLKBUF_X1 U3741 ( .A(n3695), .Z(n3689) );
  CLKBUF_X1 U3742 ( .A(n3695), .Z(n3690) );
  CLKBUF_X1 U3743 ( .A(n3695), .Z(n3691) );
  CLKBUF_X1 U3744 ( .A(n3695), .Z(n3692) );
  CLKBUF_X1 U3745 ( .A(n3695), .Z(n3693) );
  CLKBUF_X1 U3746 ( .A(n3695), .Z(n3694) );
  INV_X2 U3747 ( .A(CLK), .ZN(n4212) );
endmodule


module REG_PIPO_6_00_00_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n4, n5, n6, n7, n8, n3, n9, n10, n11, n12, n13, n14;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n14), .ZN(n2) );
  INV_X1 U3 ( .A(n1), .ZN(n13) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n2), .B1(n14), .B2(DOUT[0]), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(n12) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n2), .B1(n14), .B2(DOUT[1]), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n11) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n2), .B1(n14), .B2(DOUT[2]), .ZN(n5) );
  INV_X1 U9 ( .A(n6), .ZN(n10) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n2), .B1(n14), .B2(DOUT[3]), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n9) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n2), .B1(n14), .B2(DOUT[4]), .ZN(n7) );
  INV_X1 U13 ( .A(n8), .ZN(n3) );
  AOI22_X1 U14 ( .A1(DIN[5]), .A2(n2), .B1(n14), .B2(DOUT[5]), .ZN(n8) );
  INV_X1 U15 ( .A(EN), .ZN(n14) );
endmodule


module REG_PIPO_32_00000000_00000000_10 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_9 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_8 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_7 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n9), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n9) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n10), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n10) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n11), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n11) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n13), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n13) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n14), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n14) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n15), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_5_00_00_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n4, n5, n6, n7, n3, n8, n9, n10, n11, n12;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n12), .ZN(n2) );
  INV_X1 U3 ( .A(n1), .ZN(n11) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n2), .B1(n12), .B2(DOUT[0]), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(n10) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n2), .B1(n12), .B2(DOUT[1]), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n2), .B1(n12), .B2(DOUT[2]), .ZN(n5) );
  INV_X1 U9 ( .A(n6), .ZN(n8) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n2), .B1(n12), .B2(DOUT[3]), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n3) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n2), .B1(n12), .B2(DOUT[4]), .ZN(n7) );
  INV_X1 U13 ( .A(EN), .ZN(n12) );
endmodule


module REG_PIPO_5_00_00_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(n11) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  INV_X1 U5 ( .A(n16), .ZN(n10) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  INV_X1 U9 ( .A(n14), .ZN(n8) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  INV_X1 U11 ( .A(n13), .ZN(n3) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  INV_X1 U13 ( .A(EN), .ZN(n12) );
endmodule


module ALU_DATA_W32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n214, net17647, net17644, net17641, net17624, net17612, net17555,
         net17554, net17553, net17552, net17551, net17550, net17549, net17548,
         net17547, net17546, net17545, net17544, net17543, net17530, net17529,
         net17528, net17525, net17521, net17520, net17519, net17518, net17515,
         net17511, net17510, net17509, net17508, net17505, net17504, net17501,
         net17500, net17499, net17498, net17495, net17494, net17491, net17490,
         net17489, net17488, net17485, net17484, net17481, net17480, net17479,
         net17478, net17469, net17468, net17467, net17465, net18938, net18952,
         net18953, net18959, net18961, net18965, net18967, net18971, net18973,
         net26762, net26771, net26785, net32861, net32902, net32940, net33002,
         net32999, net17542, net17531, net34081, net34413, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n73, n74, n75, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213;

  AND2_X1 U1 ( .A1(n200), .A2(net17554), .ZN(net17479) );
  INV_X1 U2 ( .A(net17510), .ZN(n103) );
  AND2_X1 U3 ( .A1(n207), .A2(net17548), .ZN(net17509) );
  INV_X1 U4 ( .A(n41), .ZN(n65) );
  NOR2_X1 U5 ( .A1(n40), .A2(n42), .ZN(n44) );
  NOR2_X1 U6 ( .A1(net17500), .A2(n41), .ZN(n40) );
  AND2_X1 U7 ( .A1(net17550), .A2(net17551), .ZN(n43) );
  AND2_X1 U8 ( .A1(n9), .A2(n161), .ZN(n154) );
  NAND2_X1 U9 ( .A1(net17530), .A2(net17531), .ZN(n134) );
  INV_X1 U10 ( .A(net17624), .ZN(n89) );
  AND2_X1 U11 ( .A1(net17549), .A2(net17548), .ZN(n100) );
  NAND2_X1 U12 ( .A1(net17499), .A2(net17498), .ZN(n41) );
  AND2_X1 U13 ( .A1(n147), .A2(n122), .ZN(n73) );
  AND2_X1 U14 ( .A1(net17554), .A2(net17555), .ZN(n54) );
  INV_X1 U15 ( .A(net17481), .ZN(n59) );
  NAND2_X1 U16 ( .A1(n46), .A2(n2), .ZN(n47) );
  OAI21_X1 U17 ( .B1(net17489), .B2(n45), .A(n1), .ZN(n48) );
  NOR2_X1 U18 ( .A1(net17484), .A2(net17485), .ZN(n46) );
  AND2_X1 U19 ( .A1(net17478), .A2(net17479), .ZN(n52) );
  INV_X1 U20 ( .A(net17488), .ZN(n57) );
  NOR2_X1 U21 ( .A1(net17495), .A2(net17494), .ZN(n37) );
  AND2_X1 U22 ( .A1(n3), .A2(n7), .ZN(n116) );
  AND2_X1 U23 ( .A1(n8), .A2(n154), .ZN(n153) );
  OR2_X1 U24 ( .A1(n170), .A2(A[27]), .ZN(n1) );
  AND2_X1 U25 ( .A1(n199), .A2(n197), .ZN(n2) );
  AND2_X1 U26 ( .A1(n1), .A2(n200), .ZN(n3) );
  OR2_X1 U27 ( .A1(A[3]), .A2(n138), .ZN(n4) );
  AND2_X1 U28 ( .A1(net17518), .A2(net17624), .ZN(n5) );
  AND2_X1 U29 ( .A1(net18961), .A2(net17549), .ZN(n6) );
  AND2_X1 U30 ( .A1(net17468), .A2(n199), .ZN(n7) );
  AND2_X1 U31 ( .A1(net17489), .A2(net17490), .ZN(n8) );
  AND2_X1 U32 ( .A1(net18973), .A2(net17553), .ZN(n9) );
  AND2_X1 U33 ( .A1(net17529), .A2(net17530), .ZN(n10) );
  AND2_X1 U34 ( .A1(n2), .A2(net17555), .ZN(n11) );
  AND2_X1 U35 ( .A1(net18959), .A2(n207), .ZN(n12) );
  AND2_X1 U36 ( .A1(net17478), .A2(n201), .ZN(n13) );
  AND2_X1 U37 ( .A1(net17488), .A2(n204), .ZN(n14) );
  AND2_X1 U38 ( .A1(n93), .A2(net17520), .ZN(n15) );
  AND2_X1 U39 ( .A1(net18965), .A2(n205), .ZN(n16) );
  OR2_X1 U40 ( .A1(net17505), .A2(net17504), .ZN(n17) );
  AND2_X1 U41 ( .A1(n101), .A2(n210), .ZN(n18) );
  CLKBUF_X1 U42 ( .A(A[6]), .Z(n19) );
  AND2_X1 U43 ( .A1(n20), .A2(n21), .ZN(n144) );
  NAND2_X1 U44 ( .A1(n154), .A2(n157), .ZN(n20) );
  OR2_X1 U45 ( .A1(n160), .A2(n13), .ZN(n21) );
  CLKBUF_X1 U46 ( .A(net17553), .Z(n22) );
  AND2_X1 U47 ( .A1(n31), .A2(n142), .ZN(n23) );
  AND2_X1 U48 ( .A1(n149), .A2(net17612), .ZN(n24) );
  CLKBUF_X1 U49 ( .A(net17511), .Z(n25) );
  INV_X1 U50 ( .A(net17480), .ZN(n58) );
  CLKBUF_X1 U51 ( .A(n125), .Z(n118) );
  NOR2_X1 U52 ( .A1(net17501), .A2(n41), .ZN(n42) );
  AND2_X1 U53 ( .A1(net17519), .A2(net17520), .ZN(n26) );
  NOR2_X1 U54 ( .A1(net17544), .A2(n89), .ZN(n90) );
  OR2_X2 U55 ( .A1(n188), .A2(A[8]), .ZN(net17624) );
  NOR2_X1 U56 ( .A1(n27), .A2(n28), .ZN(n79) );
  NOR2_X1 U57 ( .A1(n158), .A2(n150), .ZN(n27) );
  NAND2_X1 U58 ( .A1(n12), .A2(n164), .ZN(n28) );
  NAND4_X1 U59 ( .A1(net17552), .A2(n22), .A3(net17491), .A4(net17490), .ZN(
        n39) );
  NAND2_X1 U60 ( .A1(net17553), .A2(net17552), .ZN(n45) );
  AND2_X1 U61 ( .A1(n208), .A2(net17546), .ZN(n29) );
  AND2_X1 U62 ( .A1(net32861), .A2(n117), .ZN(n30) );
  INV_X1 U63 ( .A(n25), .ZN(n104) );
  CLKBUF_X1 U64 ( .A(net32902), .Z(net26762) );
  INV_X1 U65 ( .A(n29), .ZN(n102) );
  NOR2_X1 U66 ( .A1(net17518), .A2(n92), .ZN(n94) );
  NAND2_X1 U67 ( .A1(n23), .A2(n141), .ZN(n139) );
  NOR2_X1 U68 ( .A1(n162), .A2(n143), .ZN(n31) );
  NOR2_X1 U69 ( .A1(n47), .A2(n48), .ZN(n49) );
  AND3_X1 U70 ( .A1(n52), .A2(n53), .A3(net17469), .ZN(n51) );
  XNOR2_X1 U71 ( .A(A[30]), .B(B[30]), .ZN(net17469) );
  AND2_X1 U72 ( .A1(n88), .A2(n87), .ZN(n86) );
  NAND2_X1 U73 ( .A1(n213), .A2(n30), .ZN(n212) );
  OAI21_X1 U74 ( .B1(n33), .B2(n34), .A(n35), .ZN(n32) );
  AND3_X1 U75 ( .A1(net34081), .A2(n105), .A3(n15), .ZN(n33) );
  NAND3_X1 U76 ( .A1(n95), .A2(n96), .A3(n97), .ZN(n34) );
  AND3_X1 U77 ( .A1(n98), .A2(n99), .A3(n100), .ZN(n35) );
  NAND3_X1 U78 ( .A1(n51), .A2(n69), .A3(n49), .ZN(n50) );
  NAND3_X1 U79 ( .A1(net17500), .A2(net17501), .A3(n17), .ZN(n61) );
  NAND3_X1 U80 ( .A1(net17552), .A2(n57), .A3(n22), .ZN(n53) );
  NAND3_X1 U81 ( .A1(net17479), .A2(n59), .A3(net17478), .ZN(n62) );
  NAND3_X1 U82 ( .A1(net17479), .A2(n58), .A3(net17478), .ZN(n63) );
  NAND3_X1 U83 ( .A1(n32), .A2(n61), .A3(n65), .ZN(n64) );
  NAND3_X1 U84 ( .A1(n69), .A2(net17469), .A3(net17467), .ZN(n66) );
  NAND3_X1 U85 ( .A1(n63), .A2(n62), .A3(n54), .ZN(n67) );
  NAND3_X1 U86 ( .A1(n55), .A2(n69), .A3(n67), .ZN(n68) );
  NAND3_X1 U87 ( .A1(n64), .A2(n44), .A3(n43), .ZN(n38) );
  AND3_X1 U88 ( .A1(net17469), .A2(n2), .A3(n1), .ZN(n55) );
  OAI21_X1 U89 ( .B1(n36), .B2(n50), .A(n56), .ZN(n60) );
  INV_X1 U90 ( .A(n60), .ZN(net17465) );
  AND2_X1 U91 ( .A1(n68), .A2(n66), .ZN(n56) );
  BUF_X1 U92 ( .A(net17468), .Z(n69) );
  AOI21_X1 U93 ( .B1(n38), .B2(n37), .A(n39), .ZN(n36) );
  NAND2_X1 U94 ( .A1(n139), .A2(n70), .ZN(n203) );
  AND2_X1 U95 ( .A1(n140), .A2(n14), .ZN(n70) );
  INV_X1 U96 ( .A(net17546), .ZN(n92) );
  AND2_X1 U97 ( .A1(n208), .A2(net17546), .ZN(net17519) );
  AND2_X1 U98 ( .A1(net17508), .A2(net17612), .ZN(n71) );
  OAI21_X1 U99 ( .B1(n90), .B2(n91), .A(n101), .ZN(n105) );
  AND3_X1 U100 ( .A1(net17546), .A2(net17521), .A3(net17547), .ZN(n93) );
  AOI21_X1 U101 ( .B1(n94), .B2(net17547), .A(net17515), .ZN(n95) );
  AND2_X1 U102 ( .A1(n198), .A2(n165), .ZN(GE) );
  NOR2_X1 U103 ( .A1(net17545), .A2(net34413), .ZN(n91) );
  CLKBUF_X1 U104 ( .A(B[1]), .Z(n74) );
  NOR2_X1 U105 ( .A1(net26771), .A2(A[0]), .ZN(n75) );
  AOI21_X1 U106 ( .B1(n194), .B2(A[31]), .A(n195), .ZN(LE) );
  OR2_X1 U107 ( .A1(n184), .A2(A[13]), .ZN(n77) );
  OR2_X1 U108 ( .A1(n184), .A2(A[13]), .ZN(net17508) );
  AND2_X1 U109 ( .A1(net17528), .A2(net26762), .ZN(n78) );
  NAND2_X1 U110 ( .A1(n146), .A2(n79), .ZN(n141) );
  INV_X1 U111 ( .A(net17525), .ZN(n101) );
  AND3_X1 U112 ( .A1(net17508), .A2(net17612), .A3(net17509), .ZN(n97) );
  AND2_X1 U113 ( .A1(n111), .A2(n4), .ZN(n80) );
  AND2_X1 U114 ( .A1(n114), .A2(n83), .ZN(n81) );
  NOR2_X1 U115 ( .A1(n81), .A2(n82), .ZN(n165) );
  AND2_X1 U116 ( .A1(n192), .A2(n167), .ZN(n82) );
  AND2_X1 U117 ( .A1(n107), .A2(n192), .ZN(n83) );
  NAND2_X1 U118 ( .A1(n152), .A2(n86), .ZN(n84) );
  AND2_X1 U119 ( .A1(n84), .A2(n85), .ZN(n166) );
  OR2_X1 U120 ( .A1(n167), .A2(n107), .ZN(n85) );
  INV_X1 U121 ( .A(n167), .ZN(n87) );
  AND2_X1 U122 ( .A1(n116), .A2(n144), .ZN(n88) );
  NAND2_X1 U123 ( .A1(net17641), .A2(n80), .ZN(n213) );
  NAND3_X1 U124 ( .A1(net17546), .A2(net17547), .A3(n102), .ZN(n96) );
  NAND3_X1 U125 ( .A1(n77), .A2(n104), .A3(net17509), .ZN(n98) );
  NAND3_X1 U126 ( .A1(n77), .A2(n103), .A3(net17509), .ZN(n99) );
  NAND2_X1 U127 ( .A1(n110), .A2(A[2]), .ZN(n106) );
  NOR2_X1 U128 ( .A1(n108), .A2(n124), .ZN(n107) );
  NOR2_X1 U129 ( .A1(n115), .A2(n11), .ZN(n108) );
  NAND2_X1 U130 ( .A1(net17624), .A2(net17521), .ZN(net34413) );
  NOR2_X1 U131 ( .A1(n110), .A2(A[2]), .ZN(n109) );
  INV_X1 U132 ( .A(B[2]), .ZN(n110) );
  OR2_X1 U133 ( .A1(A[2]), .A2(net26785), .ZN(n111) );
  AND2_X1 U134 ( .A1(net17624), .A2(net17521), .ZN(n112) );
  NAND2_X1 U135 ( .A1(A[3]), .A2(n138), .ZN(n113) );
  NAND2_X1 U136 ( .A1(n152), .A2(n88), .ZN(n114) );
  INV_X1 U137 ( .A(n7), .ZN(n115) );
  CLKBUF_X1 U138 ( .A(net17543), .Z(n117) );
  NAND2_X1 U139 ( .A1(A[0]), .A2(net26771), .ZN(n130) );
  NOR2_X1 U140 ( .A1(n189), .A2(A[7]), .ZN(net17525) );
  NAND2_X1 U141 ( .A1(n132), .A2(n4), .ZN(n128) );
  AND2_X1 U142 ( .A1(n156), .A2(n159), .ZN(n147) );
  NAND2_X1 U143 ( .A1(n24), .A2(n119), .ZN(n155) );
  NAND2_X1 U144 ( .A1(net18953), .A2(n208), .ZN(n119) );
  NAND2_X1 U145 ( .A1(n5), .A2(n120), .ZN(n122) );
  NAND2_X1 U146 ( .A1(n112), .A2(net17545), .ZN(n120) );
  NAND2_X1 U147 ( .A1(n130), .A2(n125), .ZN(n129) );
  INV_X1 U148 ( .A(A[1]), .ZN(n125) );
  AND2_X1 U149 ( .A1(n148), .A2(n26), .ZN(n156) );
  AND2_X1 U150 ( .A1(net17529), .A2(net17528), .ZN(n136) );
  NOR2_X1 U151 ( .A1(n127), .A2(n128), .ZN(n126) );
  NAND2_X1 U152 ( .A1(n209), .A2(n123), .ZN(n121) );
  AND2_X1 U153 ( .A1(n18), .A2(n5), .ZN(n123) );
  NAND2_X1 U154 ( .A1(net17469), .A2(n196), .ZN(n124) );
  NAND3_X1 U155 ( .A1(A[1]), .A2(net26771), .A3(A[0]), .ZN(n137) );
  NAND3_X1 U156 ( .A1(n109), .A2(n113), .A3(net17542), .ZN(n133) );
  NOR2_X1 U157 ( .A1(net34413), .A2(net17525), .ZN(n135) );
  NAND2_X1 U158 ( .A1(net17543), .A2(n106), .ZN(n131) );
  OAI221_X1 U159 ( .B1(net32999), .B2(A[4]), .C1(n129), .C2(n131), .A(n133), 
        .ZN(n127) );
  AOI21_X1 U160 ( .B1(net17644), .B2(n125), .A(B[1]), .ZN(net17647) );
  OAI211_X1 U161 ( .C1(n126), .C2(n134), .A(n135), .B(n136), .ZN(net34081) );
  OAI211_X1 U162 ( .C1(n75), .C2(n118), .A(net33002), .B(net18938), .ZN(
        net17641) );
  NAND4_X1 U163 ( .A1(n113), .A2(net17542), .A3(n74), .A4(n137), .ZN(n132) );
  INV_X1 U164 ( .A(B[0]), .ZN(net26771) );
  NOR2_X1 U165 ( .A1(net18952), .A2(A[11]), .ZN(net17515) );
  INV_X1 U166 ( .A(B[3]), .ZN(n138) );
  NAND2_X1 U167 ( .A1(A[3]), .A2(n138), .ZN(net17543) );
  NAND2_X1 U168 ( .A1(net32999), .A2(A[4]), .ZN(net17531) );
  AND2_X1 U169 ( .A1(net17531), .A2(net32902), .ZN(net32861) );
  INV_X1 U170 ( .A(B[4]), .ZN(net32999) );
  OR2_X1 U171 ( .A1(net32999), .A2(A[4]), .ZN(net32902) );
  NAND2_X1 U172 ( .A1(net26785), .A2(A[2]), .ZN(net17542) );
  AND2_X1 U173 ( .A1(n111), .A2(net17542), .ZN(net33002) );
  OR2_X1 U174 ( .A1(n143), .A2(n16), .ZN(n140) );
  OR2_X1 U175 ( .A1(n163), .A2(n6), .ZN(n142) );
  NAND2_X1 U176 ( .A1(n211), .A2(n10), .ZN(n209) );
  CLKBUF_X1 U177 ( .A(net17465), .Z(net32940) );
  NAND2_X1 U178 ( .A1(net18967), .A2(net17551), .ZN(n143) );
  NAND2_X1 U179 ( .A1(n212), .A2(n78), .ZN(n211) );
  AND2_X1 U180 ( .A1(net17465), .A2(n151), .ZN(n145) );
  NAND2_X1 U181 ( .A1(n121), .A2(n73), .ZN(n146) );
  AND2_X1 U182 ( .A1(n149), .A2(net17612), .ZN(n148) );
  AND2_X1 U183 ( .A1(net17511), .A2(net17547), .ZN(n149) );
  AND2_X1 U184 ( .A1(n155), .A2(n71), .ZN(n150) );
  OR2_X1 U185 ( .A1(B[30]), .A2(n193), .ZN(n151) );
  NAND2_X1 U186 ( .A1(net32940), .A2(n151), .ZN(n194) );
  NAND2_X1 U187 ( .A1(n203), .A2(n153), .ZN(n152) );
  NAND2_X1 U188 ( .A1(net18971), .A2(n202), .ZN(n157) );
  NAND2_X1 U189 ( .A1(net17509), .A2(net17510), .ZN(n158) );
  INV_X1 U190 ( .A(n158), .ZN(n159) );
  NAND2_X1 U191 ( .A1(net17479), .A2(net17480), .ZN(n160) );
  INV_X1 U192 ( .A(n160), .ZN(n161) );
  NAND2_X1 U193 ( .A1(net17499), .A2(net17500), .ZN(n162) );
  NAND2_X1 U194 ( .A1(net17498), .A2(n206), .ZN(n163) );
  INV_X1 U195 ( .A(n163), .ZN(n164) );
  AND2_X1 U196 ( .A1(n193), .A2(B[30]), .ZN(n167) );
  INV_X1 U197 ( .A(net17484), .ZN(net18973) );
  INV_X1 U198 ( .A(net17485), .ZN(net18971) );
  INV_X1 U199 ( .A(net17504), .ZN(net18961) );
  INV_X1 U200 ( .A(net17505), .ZN(net18959) );
  INV_X1 U201 ( .A(net17494), .ZN(net18967) );
  INV_X1 U202 ( .A(net17495), .ZN(net18965) );
  INV_X1 U203 ( .A(B[11]), .ZN(net18952) );
  INV_X1 U204 ( .A(B[7]), .ZN(n189) );
  INV_X1 U205 ( .A(B[26]), .ZN(n171) );
  INV_X1 U206 ( .A(B[27]), .ZN(n170) );
  INV_X1 U207 ( .A(B[19]), .ZN(n178) );
  INV_X1 U208 ( .A(B[25]), .ZN(n172) );
  INV_X1 U209 ( .A(B[24]), .ZN(n173) );
  INV_X1 U210 ( .A(B[20]), .ZN(n177) );
  INV_X1 U211 ( .A(B[23]), .ZN(n174) );
  INV_X1 U212 ( .A(B[13]), .ZN(n184) );
  INV_X1 U213 ( .A(B[15]), .ZN(n182) );
  INV_X1 U214 ( .A(B[14]), .ZN(n183) );
  INV_X1 U215 ( .A(B[22]), .ZN(n175) );
  INV_X1 U216 ( .A(B[21]), .ZN(n176) );
  INV_X1 U217 ( .A(B[8]), .ZN(n188) );
  INV_X1 U218 ( .A(B[12]), .ZN(n185) );
  INV_X1 U219 ( .A(B[18]), .ZN(n179) );
  INV_X1 U220 ( .A(B[16]), .ZN(n181) );
  INV_X1 U221 ( .A(B[17]), .ZN(n180) );
  INV_X1 U222 ( .A(B[10]), .ZN(n186) );
  INV_X1 U223 ( .A(B[5]), .ZN(n191) );
  INV_X1 U224 ( .A(B[28]), .ZN(n169) );
  INV_X1 U225 ( .A(B[29]), .ZN(n168) );
  INV_X1 U226 ( .A(B[9]), .ZN(n187) );
  INV_X1 U227 ( .A(A[30]), .ZN(n193) );
  INV_X1 U228 ( .A(A[31]), .ZN(n192) );
  INV_X1 U229 ( .A(B[6]), .ZN(n190) );
  INV_X1 U230 ( .A(B[2]), .ZN(net26785) );
  INV_X1 U231 ( .A(net17515), .ZN(net18953) );
  INV_X1 U232 ( .A(net17647), .ZN(net18938) );
  NAND2_X1 U233 ( .A1(n214), .A2(GE), .ZN(NE) );
  AOI21_X1 U234 ( .B1(n194), .B2(A[31]), .A(n195), .ZN(n214) );
  AOI21_X1 U235 ( .B1(n145), .B2(n192), .A(B[31]), .ZN(n195) );
  NAND2_X1 U236 ( .A1(n196), .A2(n197), .ZN(net17467) );
  OAI21_X1 U237 ( .B1(n166), .B2(n192), .A(B[31]), .ZN(n198) );
  NAND2_X1 U238 ( .A1(A[29]), .A2(n168), .ZN(n196) );
  OR2_X1 U239 ( .A1(n168), .A2(A[29]), .ZN(net17468) );
  NAND2_X1 U240 ( .A1(A[28]), .A2(n169), .ZN(n197) );
  OR2_X1 U241 ( .A1(n169), .A2(A[28]), .ZN(n199) );
  NAND2_X1 U242 ( .A1(A[27]), .A2(n170), .ZN(net17555) );
  NAND2_X1 U243 ( .A1(A[26]), .A2(n171), .ZN(net17554) );
  OR2_X1 U244 ( .A1(A[26]), .A2(n171), .ZN(n200) );
  NAND2_X1 U245 ( .A1(n172), .A2(A[25]), .ZN(net17480) );
  OR2_X1 U246 ( .A1(n172), .A2(A[25]), .ZN(net17478) );
  NAND2_X1 U247 ( .A1(n201), .A2(net17481), .ZN(net17484) );
  NAND2_X1 U248 ( .A1(A[24]), .A2(n173), .ZN(net17481) );
  OR2_X1 U249 ( .A1(n173), .A2(A[24]), .ZN(n201) );
  NAND2_X1 U250 ( .A1(A[23]), .A2(n174), .ZN(net17553) );
  NOR2_X1 U251 ( .A1(n174), .A2(A[23]), .ZN(net17485) );
  AND2_X1 U252 ( .A1(n202), .A2(net17552), .ZN(net17489) );
  NAND2_X1 U253 ( .A1(A[22]), .A2(n175), .ZN(net17552) );
  OR2_X1 U254 ( .A1(n175), .A2(A[22]), .ZN(n202) );
  NAND2_X1 U255 ( .A1(n176), .A2(A[21]), .ZN(net17490) );
  OR2_X1 U256 ( .A1(n176), .A2(A[21]), .ZN(net17488) );
  NAND2_X1 U257 ( .A1(n204), .A2(net17491), .ZN(net17494) );
  NAND2_X1 U258 ( .A1(A[20]), .A2(n177), .ZN(net17491) );
  OR2_X1 U259 ( .A1(n177), .A2(A[20]), .ZN(n204) );
  NAND2_X1 U260 ( .A1(A[19]), .A2(n178), .ZN(net17551) );
  NOR2_X1 U261 ( .A1(n178), .A2(A[19]), .ZN(net17495) );
  AND2_X1 U262 ( .A1(n205), .A2(net17550), .ZN(net17499) );
  NAND2_X1 U263 ( .A1(A[18]), .A2(n179), .ZN(net17550) );
  OR2_X1 U264 ( .A1(n179), .A2(A[18]), .ZN(n205) );
  NAND2_X1 U265 ( .A1(A[17]), .A2(n180), .ZN(net17500) );
  OR2_X1 U266 ( .A1(n180), .A2(A[17]), .ZN(net17498) );
  NAND2_X1 U267 ( .A1(n206), .A2(net17501), .ZN(net17504) );
  NAND2_X1 U268 ( .A1(A[16]), .A2(n181), .ZN(net17501) );
  OR2_X1 U269 ( .A1(n181), .A2(A[16]), .ZN(n206) );
  NAND2_X1 U270 ( .A1(A[15]), .A2(n182), .ZN(net17549) );
  NOR2_X1 U271 ( .A1(n182), .A2(A[15]), .ZN(net17505) );
  NAND2_X1 U272 ( .A1(A[14]), .A2(n183), .ZN(net17548) );
  OR2_X1 U273 ( .A1(n183), .A2(A[14]), .ZN(n207) );
  NAND2_X1 U274 ( .A1(A[13]), .A2(n184), .ZN(net17510) );
  NAND2_X1 U275 ( .A1(A[12]), .A2(n185), .ZN(net17511) );
  OR2_X1 U276 ( .A1(n185), .A2(A[12]), .ZN(net17612) );
  NAND2_X1 U277 ( .A1(A[11]), .A2(net18952), .ZN(net17547) );
  NAND2_X1 U278 ( .A1(A[10]), .A2(n186), .ZN(net17546) );
  OR2_X1 U279 ( .A1(n186), .A2(A[10]), .ZN(n208) );
  NAND2_X1 U280 ( .A1(A[9]), .A2(n187), .ZN(net17520) );
  OR2_X1 U281 ( .A1(n187), .A2(A[9]), .ZN(net17518) );
  NAND2_X1 U282 ( .A1(A[8]), .A2(n188), .ZN(net17521) );
  NAND2_X1 U283 ( .A1(A[7]), .A2(n189), .ZN(net17545) );
  AND2_X1 U284 ( .A1(n210), .A2(net17544), .ZN(net17529) );
  NAND2_X1 U285 ( .A1(n19), .A2(n190), .ZN(net17544) );
  OR2_X1 U286 ( .A1(n190), .A2(A[6]), .ZN(n210) );
  NAND2_X1 U287 ( .A1(A[5]), .A2(n191), .ZN(net17530) );
  OR2_X1 U288 ( .A1(n191), .A2(A[5]), .ZN(net17528) );
  NOR2_X1 U289 ( .A1(net26771), .A2(A[0]), .ZN(net17644) );
endmodule


module ALU_DATA_W32_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   net21689, net21679, net21667, net21664, net21662, net21661, net21655,
         net21654, net21653, net21652, net21650, net21649, net21645, net21644,
         net21638, net21634, net21633, net21632, net21622, net21620, net21618,
         net21617, net21615, net21614, net21609, net21607, net21605, net21601,
         net21598, net21584, net21582, net21577, net21574, net21572, net21569,
         net21568, net21567, net21566, net21565, net21563, net21561, net21558,
         net21557, net21556, net21554, net21552, net21549, net21546, net21542,
         net21537, net21536, net21535, net21532, net21530, net21525, net21524,
         net21523, net21522, net21520, net21518, net21517, net21508, net21504,
         net21500, net21493, net21491, net21488, net21487, net21485, net21484,
         net21482, net21480, net21479, net21474, net21466, net21465, net21461,
         net21457, net21456, net21455, net21454, net21453, net21436, net21433,
         net21432, net21431, net21426, net21423, net21421, net21420, net21416,
         net21413, net21409, net21406, net21405, net21404, net21402, net21401,
         net32548, net32593, net34370, net34369, net34389, net34445, net34781,
         net34842, net34844, net34856, net34876, net34879, net34885, net34890,
         net34928, net34935, net34937, net35044, net35060, net35207, net35233,
         net35301, net35338, net35362, net36879, net36888, net38259, net38387,
         net38531, net39646, net39733, net39805, net39821, net39823, net39968,
         net39744, net37566, net31997, net21647, net21643, net21642, net21641,
         net21640, net21507, net21501, net21481, net21473, net21472, net21526,
         net21519, net21516, net21513, net21512, net21511, net21510, net37701,
         net34283, net38388, net34902, net21687, net21686, net35331, net34940,
         net21553, net21545, net21544, net21539, net21538, net21509, net37698,
         net37697, net37683, net37682, net37681, net37679, net37647, net21470,
         net21579, net21543, net34887, net21677, net21670, net21594, net21425,
         net21419, net21418, net21417, net21412, net37662, net37657, net39836,
         net34941, net34780, net21611, net21610, net21603, net21593, net21590,
         net21588, net21587, net21586, net21585, net21578, net39642, net38206,
         net34905, net21674, net21669, net21668, net21411, net21410, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130;

  NAND2_X1 U3 ( .A1(n74), .A2(n1), .ZN(n73) );
  AND2_X1 U4 ( .A1(n75), .A2(net21484), .ZN(n1) );
  CLKBUF_X1 U5 ( .A(net21418), .Z(n2) );
  AND4_X1 U6 ( .A1(net21605), .A2(net21614), .A3(net21615), .A4(net21601), 
        .ZN(net31997) );
  AND2_X1 U7 ( .A1(A[17]), .A2(n108), .ZN(n3) );
  INV_X4 U8 ( .A(n3), .ZN(net21556) );
  AOI21_X2 U9 ( .B1(net21546), .B2(n47), .A(n48), .ZN(net21545) );
  NOR2_X1 U10 ( .A1(net21472), .A2(n45), .ZN(net37682) );
  INV_X1 U11 ( .A(net21473), .ZN(net37679) );
  INV_X1 U12 ( .A(A[29]), .ZN(n40) );
  OR2_X1 U13 ( .A1(A[3]), .A2(n71), .ZN(net21431) );
  INV_X1 U14 ( .A(A[30]), .ZN(n58) );
  INV_X1 U15 ( .A(net21501), .ZN(n45) );
  NAND2_X1 U16 ( .A1(A[29]), .A2(n41), .ZN(n39) );
  OAI21_X1 U17 ( .B1(net35044), .B2(net21472), .A(net21473), .ZN(net21461) );
  NOR2_X1 U18 ( .A1(net37647), .A2(n4), .ZN(net21466) );
  INV_X1 U19 ( .A(net37698), .ZN(net37647) );
  INV_X1 U20 ( .A(net34935), .ZN(net21421) );
  NAND2_X1 U21 ( .A1(net37657), .A2(n38), .ZN(net21457) );
  NAND2_X1 U22 ( .A1(A[29]), .A2(n41), .ZN(n38) );
  AND2_X1 U23 ( .A1(B[28]), .A2(net21470), .ZN(n4) );
  AND2_X1 U24 ( .A1(A[27]), .A2(n68), .ZN(n5) );
  AND2_X1 U25 ( .A1(A[23]), .A2(n61), .ZN(n6) );
  AND4_X1 U26 ( .A1(net21401), .A2(net21406), .A3(net21644), .A4(net21649), 
        .ZN(n7) );
  XOR2_X1 U27 ( .A(A[30]), .B(B[30]), .Z(n8) );
  OR2_X1 U28 ( .A1(B[30]), .A2(n58), .ZN(n9) );
  AND2_X1 U29 ( .A1(net21485), .A2(net21501), .ZN(n10) );
  AND2_X1 U30 ( .A1(net21501), .A2(net21482), .ZN(n11) );
  INV_X1 U31 ( .A(net35362), .ZN(net21405) );
  AND2_X1 U32 ( .A1(A[8]), .A2(n124), .ZN(net35362) );
  AND2_X2 U33 ( .A1(B[0]), .A2(n129), .ZN(net34885) );
  INV_X1 U34 ( .A(net21633), .ZN(n12) );
  OAI21_X1 U35 ( .B1(net21632), .B2(net21633), .A(n109), .ZN(n13) );
  INV_X1 U36 ( .A(net21417), .ZN(n14) );
  XNOR2_X1 U37 ( .A(n15), .B(n16), .ZN(DIFF[31]) );
  NAND2_X1 U38 ( .A1(n19), .A2(n20), .ZN(n15) );
  XOR2_X1 U39 ( .A(B[31]), .B(A[31]), .Z(n16) );
  BUF_X1 U40 ( .A(net21410), .Z(n17) );
  CLKBUF_X1 U41 ( .A(net21574), .Z(n18) );
  NAND2_X1 U42 ( .A1(net37697), .A2(n22), .ZN(n19) );
  OR2_X1 U43 ( .A1(n21), .A2(n26), .ZN(n20) );
  INV_X1 U44 ( .A(net37701), .ZN(n21) );
  AND2_X1 U45 ( .A1(net37657), .A2(net37701), .ZN(n22) );
  CLKBUF_X1 U46 ( .A(n17), .Z(n23) );
  CLKBUF_X1 U47 ( .A(net21585), .Z(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(net37681), .A(net37698), .ZN(n25) );
  NAND2_X1 U49 ( .A1(n46), .A2(A[28]), .ZN(net37698) );
  AND2_X1 U50 ( .A1(n39), .A2(n9), .ZN(n26) );
  NAND2_X1 U51 ( .A1(B[30]), .A2(n58), .ZN(net37701) );
  AND2_X1 U52 ( .A1(net39642), .A2(net21411), .ZN(net21668) );
  NAND2_X1 U53 ( .A1(net21669), .A2(net21668), .ZN(net21594) );
  NAND2_X1 U54 ( .A1(net34905), .A2(net21410), .ZN(net39642) );
  NAND2_X1 U55 ( .A1(net38206), .A2(net21674), .ZN(net21411) );
  NAND2_X1 U56 ( .A1(n23), .A2(net21411), .ZN(net21409) );
  INV_X1 U57 ( .A(B[7]), .ZN(net21674) );
  CLKBUF_X1 U58 ( .A(A[7]), .Z(net38206) );
  AND2_X1 U59 ( .A1(n27), .A2(A[6]), .ZN(net34905) );
  CLKBUF_X1 U60 ( .A(net34905), .Z(net34935) );
  INV_X1 U61 ( .A(B[6]), .ZN(n27) );
  NAND2_X1 U62 ( .A1(n28), .A2(B[7]), .ZN(net21410) );
  NAND4_X1 U63 ( .A1(net21670), .A2(net21419), .A3(net21412), .A4(n17), .ZN(
        net21669) );
  AND4_X1 U64 ( .A1(net21410), .A2(net21419), .A3(net21412), .A4(net21426), 
        .ZN(net34902) );
  INV_X1 U65 ( .A(A[7]), .ZN(n28) );
  INV_X1 U66 ( .A(A[6]), .ZN(net21677) );
  CLKBUF_X1 U67 ( .A(B[6]), .Z(net34887) );
  NAND2_X1 U68 ( .A1(net21586), .A2(net21585), .ZN(net21578) );
  NAND2_X1 U69 ( .A1(net21578), .A2(net21579), .ZN(net21543) );
  OAI21_X1 U70 ( .B1(net21587), .B2(net21588), .A(net31997), .ZN(net21586) );
  CLKBUF_X1 U71 ( .A(net21586), .Z(net34941) );
  NAND2_X1 U72 ( .A1(net21640), .A2(net21641), .ZN(net21588) );
  NOR2_X1 U73 ( .A1(net21590), .A2(net38388), .ZN(net21587) );
  AOI21_X1 U74 ( .B1(net21593), .B2(net34902), .A(net21594), .ZN(net21590) );
  NAND2_X1 U75 ( .A1(net21687), .A2(net21686), .ZN(net21593) );
  NOR2_X1 U76 ( .A1(n29), .A2(n30), .ZN(net21585) );
  NAND2_X1 U77 ( .A1(n24), .A2(net34941), .ZN(net34781) );
  NAND2_X1 U78 ( .A1(n31), .A2(net21598), .ZN(n30) );
  OAI21_X1 U79 ( .B1(n33), .B2(n32), .A(net21601), .ZN(n31) );
  INV_X1 U80 ( .A(net21609), .ZN(n32) );
  NOR2_X1 U81 ( .A1(n34), .A2(net21603), .ZN(n33) );
  INV_X1 U82 ( .A(net21615), .ZN(net21603) );
  OAI21_X1 U83 ( .B1(net36888), .B2(net21603), .A(net21609), .ZN(net21620) );
  AOI21_X1 U84 ( .B1(n37), .B2(net21605), .A(net34389), .ZN(n34) );
  AND2_X1 U85 ( .A1(n35), .A2(A[12]), .ZN(n37) );
  INV_X1 U86 ( .A(B[12]), .ZN(n35) );
  CLKBUF_X1 U87 ( .A(n35), .Z(net39968) );
  NOR2_X1 U88 ( .A1(net21610), .A2(net21611), .ZN(n29) );
  NAND2_X1 U89 ( .A1(n7), .A2(net31997), .ZN(net21611) );
  NAND2_X1 U90 ( .A1(net34902), .A2(net34780), .ZN(net21610) );
  AND3_X1 U91 ( .A1(net39733), .A2(net39836), .A3(n36), .ZN(net34780) );
  NOR2_X1 U92 ( .A1(net34445), .A2(net34885), .ZN(n36) );
  BUF_X1 U93 ( .A(net21436), .Z(net39836) );
  NAND3_X1 U94 ( .A1(net39733), .A2(net39836), .A3(net34937), .ZN(net21618) );
  CLKBUF_X1 U95 ( .A(net39836), .Z(net35060) );
  NAND2_X1 U96 ( .A1(net37697), .A2(net37657), .ZN(net37662) );
  NAND2_X1 U97 ( .A1(net37662), .A2(n39), .ZN(net38531) );
  INV_X1 U98 ( .A(B[29]), .ZN(n41) );
  NAND2_X1 U99 ( .A1(n40), .A2(B[29]), .ZN(net37657) );
  CLKBUF_X1 U100 ( .A(net21594), .Z(net35233) );
  NAND2_X1 U101 ( .A1(net21425), .A2(net21418), .ZN(net21670) );
  OR2_X1 U102 ( .A1(A[5]), .A2(n43), .ZN(net21419) );
  INV_X1 U103 ( .A(net21419), .ZN(net21417) );
  AND2_X1 U104 ( .A1(n14), .A2(n2), .ZN(net32593) );
  INV_X1 U105 ( .A(B[5]), .ZN(n43) );
  NAND2_X1 U106 ( .A1(A[5]), .A2(n43), .ZN(net21418) );
  NAND2_X1 U107 ( .A1(net34887), .A2(net21677), .ZN(net21412) );
  CLKBUF_X1 U108 ( .A(net21412), .Z(net39646) );
  OAI21_X1 U109 ( .B1(net21416), .B2(net21417), .A(n2), .ZN(net21413) );
  NAND2_X1 U110 ( .A1(A[4]), .A2(n42), .ZN(net21425) );
  CLKBUF_X1 U111 ( .A(net21425), .Z(net34844) );
  INV_X1 U112 ( .A(B[4]), .ZN(n42) );
  OAI21_X1 U113 ( .B1(net21543), .B2(net21544), .A(net21545), .ZN(net21538) );
  CLKBUF_X1 U114 ( .A(net21543), .Z(net35331) );
  NAND2_X1 U115 ( .A1(B[16]), .A2(n44), .ZN(net21579) );
  NAND2_X1 U116 ( .A1(net34781), .A2(net21579), .ZN(net34283) );
  NAND2_X1 U117 ( .A1(net21557), .A2(net21579), .ZN(net21582) );
  INV_X1 U118 ( .A(A[16]), .ZN(n44) );
  OAI21_X1 U119 ( .B1(net37681), .B2(n4), .A(net37698), .ZN(net37697) );
  INV_X1 U120 ( .A(A[28]), .ZN(net21470) );
  AOI21_X1 U121 ( .B1(net37683), .B2(net37682), .A(net37679), .ZN(net37681) );
  OAI21_X1 U122 ( .B1(net21509), .B2(net21510), .A(net21511), .ZN(net37683) );
  INV_X1 U123 ( .A(B[28]), .ZN(n46) );
  NAND2_X1 U124 ( .A1(net35301), .A2(net21501), .ZN(net35044) );
  OAI21_X1 U125 ( .B1(net21509), .B2(net21510), .A(net21511), .ZN(net35301) );
  OAI21_X1 U126 ( .B1(net21510), .B2(net34876), .A(net21511), .ZN(net21500) );
  NAND2_X1 U127 ( .A1(net21538), .A2(net21539), .ZN(net21509) );
  NAND2_X1 U128 ( .A1(B[20]), .A2(n51), .ZN(net21539) );
  NAND2_X1 U129 ( .A1(net21523), .A2(net21539), .ZN(net21542) );
  NAND2_X1 U130 ( .A1(net34940), .A2(net21539), .ZN(net34876) );
  INV_X1 U131 ( .A(A[20]), .ZN(n51) );
  NAND3_X1 U132 ( .A1(net21558), .A2(net21546), .A3(net21554), .ZN(net21544)
         );
  OAI21_X1 U133 ( .B1(net34283), .B2(net21544), .A(net21545), .ZN(net32548) );
  OAI21_X1 U134 ( .B1(net35331), .B2(net21544), .A(net21545), .ZN(net34940) );
  INV_X1 U135 ( .A(net21549), .ZN(n48) );
  OAI21_X1 U136 ( .B1(n49), .B2(n50), .A(net21552), .ZN(n47) );
  INV_X1 U137 ( .A(net21558), .ZN(n50) );
  OAI21_X1 U138 ( .B1(net21568), .B2(n50), .A(net21552), .ZN(net21567) );
  AOI21_X1 U139 ( .B1(net21553), .B2(net21554), .A(n3), .ZN(n49) );
  INV_X1 U140 ( .A(net21557), .ZN(net21553) );
  INV_X1 U141 ( .A(B[20]), .ZN(n52) );
  NAND2_X1 U142 ( .A1(A[20]), .A2(n52), .ZN(net21523) );
  NAND2_X1 U143 ( .A1(net21552), .A2(net21558), .ZN(net21572) );
  NAND2_X1 U144 ( .A1(net21549), .A2(net21546), .ZN(net21566) );
  NAND4_X1 U145 ( .A1(net21401), .A2(net21649), .A3(net21644), .A4(net21406), 
        .ZN(net38388) );
  OAI21_X1 U146 ( .B1(net21638), .B2(net38388), .A(net37566), .ZN(net21634) );
  INV_X1 U147 ( .A(net34902), .ZN(net21617) );
  NAND4_X1 U148 ( .A1(net21455), .A2(n53), .A3(net21436), .A4(net21431), .ZN(
        net21687) );
  AND2_X1 U149 ( .A1(net21686), .A2(net21687), .ZN(net34928) );
  NAND2_X1 U150 ( .A1(net21454), .A2(net21563), .ZN(n53) );
  AOI21_X1 U151 ( .B1(n56), .B2(net21431), .A(n54), .ZN(net21686) );
  INV_X1 U152 ( .A(net21432), .ZN(n54) );
  AND2_X1 U153 ( .A1(A[2]), .A2(n55), .ZN(n56) );
  INV_X1 U154 ( .A(B[2]), .ZN(n55) );
  NAND2_X1 U155 ( .A1(A[2]), .A2(n55), .ZN(net21433) );
  INV_X1 U156 ( .A(net21649), .ZN(net21647) );
  OAI21_X1 U157 ( .B1(net21642), .B2(net21643), .A(net21644), .ZN(net21640) );
  NAND2_X1 U158 ( .A1(net21641), .A2(net21644), .ZN(net21652) );
  CLKBUF_X1 U159 ( .A(net21406), .Z(net35338) );
  NAND2_X1 U160 ( .A1(net21404), .A2(net21406), .ZN(net21664) );
  CLKBUF_X1 U161 ( .A(net21426), .Z(net34842) );
  NAND2_X1 U162 ( .A1(net21554), .A2(net21574), .ZN(n57) );
  NAND2_X1 U163 ( .A1(net21556), .A2(net21554), .ZN(net21577) );
  NAND2_X1 U164 ( .A1(n57), .A2(net21556), .ZN(net21569) );
  NAND2_X1 U165 ( .A1(net34283), .A2(net21557), .ZN(net21574) );
  NAND3_X1 U166 ( .A1(net21518), .A2(net21512), .A3(net21520), .ZN(net21510)
         );
  AOI21_X1 U167 ( .B1(net21512), .B2(net21513), .A(n6), .ZN(net21511) );
  NOR2_X1 U168 ( .A1(net21526), .A2(n6), .ZN(net21525) );
  INV_X1 U169 ( .A(B[23]), .ZN(n61) );
  OAI21_X1 U170 ( .B1(n59), .B2(net21516), .A(net21517), .ZN(net21513) );
  INV_X1 U171 ( .A(net21518), .ZN(net21516) );
  AOI21_X1 U172 ( .B1(net21519), .B2(net21520), .A(n60), .ZN(n59) );
  INV_X1 U173 ( .A(net21522), .ZN(n60) );
  INV_X1 U174 ( .A(net21523), .ZN(net21519) );
  AOI21_X1 U175 ( .B1(net21518), .B2(net21530), .A(n63), .ZN(net21524) );
  NAND2_X1 U176 ( .A1(net21517), .A2(net21518), .ZN(net21532) );
  INV_X1 U177 ( .A(net21512), .ZN(net21526) );
  NAND2_X1 U178 ( .A1(net21520), .A2(net21536), .ZN(net21535) );
  NAND2_X1 U179 ( .A1(net21522), .A2(net21520), .ZN(net21537) );
  INV_X1 U180 ( .A(A[23]), .ZN(n62) );
  NAND2_X1 U181 ( .A1(B[23]), .A2(n62), .ZN(net21512) );
  INV_X1 U182 ( .A(net21517), .ZN(n63) );
  AOI21_X1 U183 ( .B1(net21474), .B2(n64), .A(n5), .ZN(net21473) );
  NOR2_X1 U184 ( .A1(net21488), .A2(n5), .ZN(net21487) );
  INV_X1 U185 ( .A(B[27]), .ZN(n68) );
  OAI21_X1 U186 ( .B1(n65), .B2(n66), .A(net21479), .ZN(n64) );
  INV_X1 U187 ( .A(net21480), .ZN(n66) );
  AOI21_X1 U188 ( .B1(net21481), .B2(net21482), .A(n67), .ZN(n65) );
  INV_X1 U189 ( .A(net21484), .ZN(n67) );
  INV_X1 U190 ( .A(net21485), .ZN(net21481) );
  NAND3_X1 U191 ( .A1(net21480), .A2(net21474), .A3(net21482), .ZN(net21472)
         );
  NAND2_X1 U192 ( .A1(B[24]), .A2(net21507), .ZN(net21501) );
  INV_X1 U193 ( .A(A[24]), .ZN(net21507) );
  NAND2_X1 U194 ( .A1(net21455), .A2(net34879), .ZN(net21561) );
  NAND2_X1 U195 ( .A1(net21455), .A2(net21456), .ZN(net21453) );
  CLKBUF_X1 U196 ( .A(net21640), .Z(net39744) );
  INV_X1 U197 ( .A(net21645), .ZN(net21643) );
  AOI21_X1 U198 ( .B1(net21402), .B2(n69), .A(net21647), .ZN(net21642) );
  INV_X1 U199 ( .A(net21647), .ZN(net39821) );
  OAI21_X1 U200 ( .B1(net21654), .B2(net21647), .A(net21645), .ZN(net21653) );
  NAND2_X1 U201 ( .A1(net38387), .A2(net35362), .ZN(n69) );
  NAND2_X1 U202 ( .A1(A[11]), .A2(n70), .ZN(net21641) );
  AND2_X1 U203 ( .A1(net39744), .A2(net21641), .ZN(net37566) );
  INV_X1 U204 ( .A(B[11]), .ZN(n70) );
  INV_X1 U205 ( .A(net21632), .ZN(net39823) );
  NOR2_X1 U206 ( .A1(n118), .A2(B[13]), .ZN(net34389) );
  CLKBUF_X1 U207 ( .A(net21402), .Z(net39805) );
  BUF_X1 U208 ( .A(net21431), .Z(net39733) );
  INV_X1 U209 ( .A(net36888), .ZN(net21622) );
  INV_X1 U210 ( .A(B[3]), .ZN(n71) );
  NAND2_X1 U211 ( .A1(n74), .A2(n72), .ZN(n91) );
  AND2_X1 U212 ( .A1(n75), .A2(net21484), .ZN(n72) );
  NAND2_X1 U213 ( .A1(B[9]), .A2(n128), .ZN(net38387) );
  CLKBUF_X1 U214 ( .A(net34389), .Z(net38259) );
  AOI21_X1 U215 ( .B1(n114), .B2(net34370), .A(net38259), .ZN(net36888) );
  INV_X1 U216 ( .A(net38259), .ZN(net21607) );
  NAND2_X1 U217 ( .A1(net35301), .A2(n11), .ZN(n74) );
  OR2_X1 U218 ( .A1(net36879), .A2(net21485), .ZN(n75) );
  INV_X1 U219 ( .A(net21482), .ZN(net36879) );
  OAI21_X2 U220 ( .B1(n82), .B2(net21617), .A(net21667), .ZN(net21404) );
  CLKBUF_X1 U221 ( .A(net21563), .Z(net35207) );
  CLKBUF_X1 U222 ( .A(B[1]), .Z(n76) );
  INV_X1 U223 ( .A(net34885), .ZN(net21565) );
  NOR2_X1 U224 ( .A1(net34885), .A2(net34445), .ZN(net34937) );
  XNOR2_X1 U225 ( .A(net38531), .B(n8), .ZN(DIFF[30]) );
  CLKBUF_X1 U226 ( .A(B[4]), .Z(net34890) );
  CLKBUF_X1 U227 ( .A(net21454), .Z(net34879) );
  CLKBUF_X1 U228 ( .A(net38387), .Z(net34856) );
  AND2_X1 U229 ( .A1(n76), .A2(n126), .ZN(net34445) );
  CLKBUF_X1 U230 ( .A(net34781), .Z(net34369) );
  CLKBUF_X1 U231 ( .A(net21605), .Z(net34370) );
  XOR2_X1 U232 ( .A(net32593), .B(net21420), .Z(DIFF[5]) );
  XOR2_X1 U233 ( .A(n80), .B(net21409), .Z(DIFF[7]) );
  XNOR2_X1 U234 ( .A(net34369), .B(net21582), .ZN(DIFF[16]) );
  NAND2_X1 U235 ( .A1(net34928), .A2(net21618), .ZN(n84) );
  XNOR2_X1 U236 ( .A(net21577), .B(n18), .ZN(DIFF[17]) );
  XNOR2_X1 U237 ( .A(n95), .B(n96), .ZN(DIFF[25]) );
  XNOR2_X1 U238 ( .A(net21537), .B(net21536), .ZN(DIFF[21]) );
  XNOR2_X1 U239 ( .A(n73), .B(n92), .ZN(DIFF[26]) );
  XNOR2_X1 U240 ( .A(net21572), .B(net21569), .ZN(DIFF[18]) );
  XNOR2_X1 U241 ( .A(net21567), .B(net21566), .ZN(DIFF[19]) );
  XNOR2_X1 U242 ( .A(net21504), .B(n10), .ZN(DIFF[24]) );
  XNOR2_X1 U243 ( .A(n110), .B(net21620), .ZN(DIFF[15]) );
  XNOR2_X1 U244 ( .A(n83), .B(n84), .ZN(DIFF[4]) );
  NAND2_X1 U245 ( .A1(net34844), .A2(net34842), .ZN(n83) );
  XOR2_X1 U246 ( .A(n77), .B(n78), .Z(DIFF[9]) );
  NAND2_X1 U247 ( .A1(net34856), .A2(net39805), .ZN(n78) );
  XNOR2_X1 U248 ( .A(n81), .B(net21413), .ZN(DIFF[6]) );
  NAND2_X1 U249 ( .A1(net39646), .A2(net21421), .ZN(n81) );
  AOI21_X1 U250 ( .B1(net39646), .B2(net21413), .A(net34935), .ZN(n80) );
  XOR2_X1 U251 ( .A(net21654), .B(n120), .Z(DIFF[10]) );
  NAND2_X1 U252 ( .A1(net21405), .A2(net35338), .ZN(n79) );
  NAND2_X1 U253 ( .A1(net35207), .A2(net21565), .ZN(DIFF[0]) );
  XNOR2_X1 U254 ( .A(net21561), .B(net21456), .ZN(DIFF[1]) );
  AOI21_X1 U255 ( .B1(n91), .B2(net21480), .A(net21493), .ZN(n90) );
  OAI21_X1 U256 ( .B1(net21632), .B2(net21633), .A(n109), .ZN(n114) );
  OAI21_X1 U257 ( .B1(net21423), .B2(n82), .A(net34844), .ZN(net21420) );
  NAND2_X1 U258 ( .A1(net21607), .A2(net34370), .ZN(n117) );
  NAND2_X1 U259 ( .A1(net35044), .A2(net21485), .ZN(n95) );
  NAND2_X1 U260 ( .A1(net34876), .A2(net21523), .ZN(net21536) );
  NAND2_X1 U261 ( .A1(net21535), .A2(net21522), .ZN(net21530) );
  OAI21_X1 U262 ( .B1(net21662), .B2(n77), .A(net21402), .ZN(net21661) );
  XNOR2_X1 U263 ( .A(net21465), .B(net21466), .ZN(DIFF[28]) );
  XNOR2_X1 U264 ( .A(n89), .B(n88), .ZN(DIFF[2]) );
  NAND2_X1 U265 ( .A1(net35060), .A2(net21433), .ZN(n89) );
  XNOR2_X1 U266 ( .A(n85), .B(n86), .ZN(DIFF[3]) );
  NAND2_X1 U267 ( .A1(net39733), .A2(net21432), .ZN(n86) );
  XNOR2_X1 U268 ( .A(net21457), .B(n25), .ZN(DIFF[29]) );
  XNOR2_X1 U269 ( .A(net21530), .B(net21532), .ZN(DIFF[22]) );
  XNOR2_X1 U270 ( .A(n90), .B(net21487), .ZN(DIFF[27]) );
  XNOR2_X1 U271 ( .A(net21524), .B(net21525), .ZN(DIFF[23]) );
  XNOR2_X1 U272 ( .A(n113), .B(net21622), .ZN(DIFF[14]) );
  NAND2_X1 U273 ( .A1(net21609), .A2(net21615), .ZN(n113) );
  XNOR2_X1 U274 ( .A(n119), .B(n12), .ZN(DIFF[12]) );
  NAND2_X1 U275 ( .A1(n109), .A2(net39823), .ZN(n119) );
  NAND2_X1 U276 ( .A1(net21479), .A2(net21480), .ZN(n92) );
  NAND2_X1 U277 ( .A1(net21484), .A2(net21482), .ZN(n96) );
  NAND2_X1 U278 ( .A1(net21453), .A2(net34879), .ZN(n88) );
  NAND2_X1 U279 ( .A1(net21598), .A2(net21601), .ZN(n110) );
  NAND2_X1 U280 ( .A1(net21645), .A2(net39821), .ZN(n120) );
  NAND2_X1 U281 ( .A1(net21433), .A2(n87), .ZN(n85) );
  NAND2_X1 U282 ( .A1(n88), .A2(net35060), .ZN(n87) );
  AND2_X1 U283 ( .A1(net21664), .A2(net21405), .ZN(n77) );
  NAND2_X1 U284 ( .A1(net34885), .A2(net35207), .ZN(net21456) );
  INV_X1 U285 ( .A(A[1]), .ZN(n126) );
  NAND2_X1 U286 ( .A1(A[26]), .A2(n94), .ZN(net21479) );
  INV_X1 U287 ( .A(B[26]), .ZN(n94) );
  NAND2_X1 U288 ( .A1(A[25]), .A2(n98), .ZN(net21484) );
  INV_X1 U289 ( .A(B[25]), .ZN(n98) );
  NAND2_X1 U290 ( .A1(A[24]), .A2(net21508), .ZN(net21485) );
  INV_X1 U291 ( .A(B[24]), .ZN(net21508) );
  NAND2_X1 U292 ( .A1(A[18]), .A2(n106), .ZN(net21552) );
  INV_X1 U293 ( .A(B[18]), .ZN(n106) );
  NAND2_X1 U294 ( .A1(A[21]), .A2(n102), .ZN(net21522) );
  INV_X1 U295 ( .A(B[21]), .ZN(n102) );
  NAND2_X1 U296 ( .A1(A[22]), .A2(n100), .ZN(net21517) );
  INV_X1 U297 ( .A(B[22]), .ZN(n100) );
  INV_X1 U298 ( .A(B[8]), .ZN(n124) );
  NAND2_X1 U299 ( .A1(A[16]), .A2(net21584), .ZN(net21557) );
  INV_X1 U300 ( .A(B[16]), .ZN(net21584) );
  INV_X1 U301 ( .A(B[17]), .ZN(n108) );
  NAND2_X1 U302 ( .A1(A[12]), .A2(net39968), .ZN(n109) );
  NAND2_X1 U303 ( .A1(A[9]), .A2(n123), .ZN(net21402) );
  INV_X1 U304 ( .A(B[9]), .ZN(n123) );
  NAND2_X1 U305 ( .A1(A[15]), .A2(n112), .ZN(net21598) );
  INV_X1 U306 ( .A(B[15]), .ZN(n112) );
  NAND2_X1 U307 ( .A1(A[19]), .A2(n104), .ZN(net21549) );
  INV_X1 U308 ( .A(B[19]), .ZN(n104) );
  NAND2_X1 U309 ( .A1(B[9]), .A2(n128), .ZN(net21401) );
  INV_X1 U310 ( .A(A[9]), .ZN(n128) );
  NAND2_X1 U311 ( .A1(B[25]), .A2(n97), .ZN(net21482) );
  INV_X1 U312 ( .A(A[25]), .ZN(n97) );
  NAND2_X1 U313 ( .A1(B[21]), .A2(n101), .ZN(net21520) );
  INV_X1 U314 ( .A(A[21]), .ZN(n101) );
  NAND2_X1 U315 ( .A1(B[8]), .A2(n125), .ZN(net21406) );
  INV_X1 U316 ( .A(A[8]), .ZN(n125) );
  NAND2_X1 U317 ( .A1(B[11]), .A2(net21655), .ZN(net21644) );
  INV_X1 U318 ( .A(A[11]), .ZN(net21655) );
  NAND2_X1 U319 ( .A1(B[22]), .A2(n99), .ZN(net21518) );
  INV_X1 U320 ( .A(A[22]), .ZN(n99) );
  NAND2_X1 U321 ( .A1(B[26]), .A2(n93), .ZN(net21480) );
  INV_X1 U322 ( .A(A[26]), .ZN(n93) );
  NAND2_X1 U323 ( .A1(net34890), .A2(net21679), .ZN(net21426) );
  NAND2_X1 U324 ( .A1(B[19]), .A2(n103), .ZN(net21546) );
  INV_X1 U325 ( .A(A[19]), .ZN(n103) );
  NAND2_X1 U326 ( .A1(B[27]), .A2(net21491), .ZN(net21474) );
  INV_X1 U327 ( .A(A[27]), .ZN(net21491) );
  NAND2_X1 U328 ( .A1(B[13]), .A2(n118), .ZN(net21605) );
  INV_X1 U329 ( .A(A[13]), .ZN(n118) );
  NAND2_X1 U330 ( .A1(B[14]), .A2(n115), .ZN(net21615) );
  INV_X1 U331 ( .A(A[14]), .ZN(n115) );
  NAND2_X1 U332 ( .A1(B[12]), .A2(net21650), .ZN(net21614) );
  INV_X1 U333 ( .A(A[12]), .ZN(net21650) );
  NAND2_X1 U334 ( .A1(B[17]), .A2(n107), .ZN(net21554) );
  INV_X1 U335 ( .A(A[17]), .ZN(n107) );
  NAND2_X1 U336 ( .A1(B[18]), .A2(n105), .ZN(net21558) );
  INV_X1 U337 ( .A(A[18]), .ZN(n105) );
  NAND2_X1 U338 ( .A1(B[15]), .A2(n111), .ZN(net21601) );
  INV_X1 U339 ( .A(A[15]), .ZN(n111) );
  NAND2_X1 U340 ( .A1(B[10]), .A2(n121), .ZN(net21649) );
  INV_X1 U341 ( .A(A[10]), .ZN(n121) );
  NAND2_X1 U342 ( .A1(A[1]), .A2(n127), .ZN(net21454) );
  NAND2_X1 U343 ( .A1(A[10]), .A2(n122), .ZN(net21645) );
  INV_X1 U344 ( .A(B[10]), .ZN(n122) );
  NAND2_X1 U345 ( .A1(A[14]), .A2(n116), .ZN(net21609) );
  INV_X1 U346 ( .A(B[14]), .ZN(n116) );
  NAND2_X1 U347 ( .A1(B[2]), .A2(net21689), .ZN(net21436) );
  NAND2_X1 U348 ( .A1(A[3]), .A2(n71), .ZN(net21432) );
  INV_X1 U349 ( .A(A[4]), .ZN(net21679) );
  INV_X1 U350 ( .A(B[0]), .ZN(n130) );
  NAND2_X1 U351 ( .A1(n76), .A2(n126), .ZN(net21455) );
  INV_X1 U352 ( .A(B[1]), .ZN(n127) );
  NAND2_X1 U353 ( .A1(A[0]), .A2(n130), .ZN(net21563) );
  INV_X1 U354 ( .A(A[0]), .ZN(n129) );
  INV_X1 U355 ( .A(A[2]), .ZN(net21689) );
  XNOR2_X1 U356 ( .A(n79), .B(net21404), .ZN(DIFF[8]) );
  INV_X1 U357 ( .A(net21420), .ZN(net21416) );
  INV_X1 U358 ( .A(net34842), .ZN(net21423) );
  INV_X1 U359 ( .A(net21461), .ZN(net21465) );
  INV_X1 U360 ( .A(net21474), .ZN(net21488) );
  INV_X1 U361 ( .A(net21479), .ZN(net21493) );
  INV_X1 U362 ( .A(net21500), .ZN(net21504) );
  XNOR2_X1 U363 ( .A(net21542), .B(net32548), .ZN(DIFF[20]) );
  INV_X1 U364 ( .A(net21569), .ZN(net21568) );
  XNOR2_X1 U365 ( .A(n117), .B(n13), .ZN(DIFF[13]) );
  INV_X1 U366 ( .A(net21634), .ZN(net21633) );
  INV_X1 U367 ( .A(net21614), .ZN(net21632) );
  INV_X1 U368 ( .A(net21404), .ZN(net21638) );
  XNOR2_X1 U369 ( .A(net21652), .B(net21653), .ZN(DIFF[11]) );
  INV_X1 U370 ( .A(net21661), .ZN(net21654) );
  INV_X1 U371 ( .A(net35233), .ZN(net21667) );
  INV_X1 U372 ( .A(n84), .ZN(n82) );
  INV_X1 U373 ( .A(net34856), .ZN(net21662) );
endmodule


module ALU_DATA_W32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   net22706, net22684, net22682, net22678, net22673, net22670, net22665,
         net22664, net22658, net22655, net22654, net22653, net22651, net22647,
         net22646, net22643, net22636, net22627, net22626, net22610, net22593,
         net22577, net22542, net22541, net22537, net22535, net22532, net22530,
         net22529, net22525, net22523, net22519, net22518, net22517, net22516,
         net22515, net22514, net22511, net22509, net22491, net22490, net22488,
         net22485, net22484, net22465, net22463, net22462, net22461, net22460,
         net22458, net22457, net22456, net22452, net22451, net22450, net22447,
         net22446, net22444, net22443, net22440, net22439, net22438, net22437,
         net22435, net22434, net22433, net22432, net31820, net31956, net34346,
         net34345, net34383, net34452, net34451, net34775, net34787, net34831,
         net34874, net34908, net34951, net35051, net35056, net35151, net35302,
         net35304, net35340, net37487, net37442, net37430, net37898, net38135,
         net38162, net38298, net38371, net38443, net38489, net38589, net35345,
         net35293, net22669, net22668, net22666, net37569, net37480, net37469,
         net35350, net35187, net22634, net38577, net22640, net22639, net22618,
         net22616, net22615, net22614, net22609, net31791, net22474, net22473,
         net22472, net22468, net22495, net22492, n1, n2, n3, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149;

  INV_X1 U2 ( .A(net22541), .ZN(n27) );
  INV_X1 U3 ( .A(net22509), .ZN(n15) );
  INV_X1 U4 ( .A(net22532), .ZN(n19) );
  INV_X1 U5 ( .A(net22495), .ZN(n22) );
  NOR2_X1 U6 ( .A1(n23), .A2(n33), .ZN(n29) );
  OAI21_X1 U7 ( .B1(net22514), .B2(n38), .A(n32), .ZN(n33) );
  NAND2_X1 U8 ( .A1(n2), .A2(n27), .ZN(n26) );
  AOI21_X1 U9 ( .B1(n15), .B2(net22517), .A(net31820), .ZN(n32) );
  INV_X1 U10 ( .A(net22514), .ZN(n20) );
  NAND2_X1 U11 ( .A1(n28), .A2(net22495), .ZN(n35) );
  NAND2_X1 U12 ( .A1(n77), .A2(n78), .ZN(net22706) );
  OAI21_X1 U13 ( .B1(net22664), .B2(net22643), .A(net22665), .ZN(n144) );
  INV_X1 U14 ( .A(n58), .ZN(n52) );
  NOR2_X1 U15 ( .A1(net31820), .A2(n16), .ZN(net22519) );
  INV_X1 U16 ( .A(net22517), .ZN(n16) );
  NAND2_X1 U17 ( .A1(net22514), .A2(net22532), .ZN(net22537) );
  AND2_X1 U18 ( .A1(n3), .A2(n17), .ZN(n1) );
  AND2_X1 U19 ( .A1(n25), .A2(net22532), .ZN(n2) );
  AND2_X1 U20 ( .A1(n29), .A2(n30), .ZN(n3) );
  AND2_X1 U21 ( .A1(net38298), .A2(net22706), .ZN(SUM[0]) );
  AND2_X1 U22 ( .A1(n115), .A2(n116), .ZN(n5) );
  AND2_X1 U23 ( .A1(n115), .A2(n116), .ZN(n10) );
  CLKBUF_X1 U24 ( .A(n7), .Z(net34345) );
  OAI21_X1 U25 ( .B1(net34345), .B2(net22634), .A(net37569), .ZN(net22437) );
  NAND2_X1 U26 ( .A1(n40), .A2(n11), .ZN(n6) );
  NAND2_X1 U27 ( .A1(net22509), .A2(net22511), .ZN(net22525) );
  INV_X1 U28 ( .A(n26), .ZN(n37) );
  NOR2_X1 U29 ( .A1(n26), .A2(n22), .ZN(n34) );
  NOR2_X1 U30 ( .A1(n20), .A2(n31), .ZN(n13) );
  AOI21_X1 U31 ( .B1(net37480), .B2(n69), .A(n70), .ZN(n7) );
  CLKBUF_X1 U32 ( .A(net22639), .Z(n8) );
  INV_X1 U33 ( .A(n5), .ZN(net34951) );
  AOI21_X1 U34 ( .B1(n8), .B2(net35345), .A(net34831), .ZN(n9) );
  OR2_X1 U35 ( .A1(B[10]), .A2(A[10]), .ZN(net22670) );
  NAND3_X1 U36 ( .A1(net22532), .A2(n27), .A3(n10), .ZN(n14) );
  INV_X1 U37 ( .A(net22515), .ZN(n21) );
  OAI211_X1 U38 ( .C1(n21), .C2(net22516), .A(net22517), .B(net22511), .ZN(n24) );
  OAI211_X1 U39 ( .C1(n21), .C2(net22516), .A(net22517), .B(net22511), .ZN(n38) );
  NOR2_X1 U40 ( .A1(n40), .A2(n38), .ZN(n23) );
  NAND2_X1 U41 ( .A1(n40), .A2(net22516), .ZN(net22530) );
  NAND2_X1 U42 ( .A1(n11), .A2(n40), .ZN(net22523) );
  INV_X1 U43 ( .A(net22542), .ZN(n18) );
  NAND2_X1 U44 ( .A1(n34), .A2(n10), .ZN(n36) );
  NAND2_X1 U45 ( .A1(n37), .A2(n5), .ZN(n17) );
  INV_X1 U46 ( .A(n24), .ZN(n25) );
  NAND2_X1 U47 ( .A1(n2), .A2(n18), .ZN(n30) );
  NAND2_X1 U48 ( .A1(n29), .A2(n30), .ZN(n28) );
  NAND2_X1 U49 ( .A1(n12), .A2(net22516), .ZN(n11) );
  CLKBUF_X1 U50 ( .A(net22515), .Z(n40) );
  AOI21_X1 U51 ( .B1(net22523), .B2(net22511), .A(n15), .ZN(net22518) );
  NAND2_X1 U52 ( .A1(n14), .A2(n13), .ZN(n12) );
  AND2_X1 U53 ( .A1(n35), .A2(n36), .ZN(net22492) );
  BUF_X1 U54 ( .A(net22542), .Z(n39) );
  NOR2_X1 U55 ( .A1(n19), .A2(n39), .ZN(n31) );
  OAI21_X1 U56 ( .B1(net22541), .B2(net34951), .A(n39), .ZN(net34346) );
  CLKBUF_X1 U57 ( .A(n12), .Z(net22529) );
  OAI21_X1 U58 ( .B1(n43), .B2(n42), .A(n44), .ZN(n41) );
  AOI21_X1 U59 ( .B1(n41), .B2(net22472), .A(net22473), .ZN(net22468) );
  INV_X1 U60 ( .A(n45), .ZN(n42) );
  OAI21_X1 U61 ( .B1(n42), .B2(net34787), .A(n44), .ZN(net34383) );
  AND2_X1 U62 ( .A1(net22492), .A2(n46), .ZN(n43) );
  NAND2_X1 U63 ( .A1(B[29]), .A2(A[29]), .ZN(n44) );
  NAND2_X1 U64 ( .A1(n44), .A2(n45), .ZN(net22490) );
  OR2_X1 U65 ( .A1(B[29]), .A2(A[29]), .ZN(n45) );
  AND2_X1 U66 ( .A1(net22492), .A2(n46), .ZN(net34787) );
  NAND2_X1 U67 ( .A1(B[28]), .A2(A[28]), .ZN(n46) );
  AND2_X1 U68 ( .A1(n46), .A2(net22495), .ZN(net31956) );
  OR2_X1 U69 ( .A1(B[28]), .A2(A[28]), .ZN(net22495) );
  XNOR2_X1 U70 ( .A(net22468), .B(net31791), .ZN(SUM[31]) );
  XOR2_X1 U71 ( .A(B[31]), .B(A[31]), .Z(net31791) );
  INV_X1 U72 ( .A(net22474), .ZN(net22473) );
  OR2_X1 U73 ( .A1(B[30]), .A2(A[30]), .ZN(net22472) );
  NAND2_X1 U74 ( .A1(net22474), .A2(net22472), .ZN(net38371) );
  NAND2_X1 U75 ( .A1(B[30]), .A2(A[30]), .ZN(net22474) );
  OAI21_X1 U76 ( .B1(net22614), .B2(net22615), .A(net22616), .ZN(net22609) );
  NAND2_X1 U77 ( .A1(net22609), .A2(net22610), .ZN(net22577) );
  INV_X1 U78 ( .A(net22618), .ZN(net22616) );
  CLKBUF_X1 U79 ( .A(net22616), .Z(net38577) );
  OAI21_X1 U80 ( .B1(n47), .B2(n48), .A(n49), .ZN(net22618) );
  INV_X1 U81 ( .A(n53), .ZN(n48) );
  NOR2_X1 U82 ( .A1(n48), .A2(n54), .ZN(net22647) );
  AOI21_X1 U83 ( .B1(n51), .B2(n50), .A(n57), .ZN(n47) );
  OAI21_X1 U84 ( .B1(n58), .B2(net22626), .A(net22627), .ZN(n51) );
  AOI21_X1 U85 ( .B1(net22639), .B2(net35345), .A(net22640), .ZN(net22614) );
  OAI21_X1 U86 ( .B1(net22666), .B2(n56), .A(net22668), .ZN(net22640) );
  INV_X1 U87 ( .A(net22669), .ZN(n56) );
  OAI21_X1 U88 ( .B1(net35293), .B2(n56), .A(net22668), .ZN(net34831) );
  OAI21_X1 U89 ( .B1(n7), .B2(net22634), .A(net35350), .ZN(net22639) );
  NAND4_X1 U90 ( .A1(net22636), .A2(n52), .A3(n50), .A4(n53), .ZN(net22615) );
  OAI21_X1 U91 ( .B1(n9), .B2(net22615), .A(net38577), .ZN(net34452) );
  NAND2_X1 U92 ( .A1(net22627), .A2(n52), .ZN(net22658) );
  NAND2_X1 U93 ( .A1(B[15]), .A2(A[15]), .ZN(n49) );
  INV_X1 U94 ( .A(n49), .ZN(n54) );
  OR2_X1 U95 ( .A1(B[15]), .A2(A[15]), .ZN(n53) );
  OR2_X2 U96 ( .A1(B[14]), .A2(A[14]), .ZN(n50) );
  AOI21_X1 U97 ( .B1(n50), .B2(net22651), .A(n57), .ZN(net22646) );
  NAND2_X1 U98 ( .A1(n55), .A2(n50), .ZN(net22653) );
  AND2_X2 U99 ( .A1(B[14]), .A2(A[14]), .ZN(n57) );
  INV_X1 U100 ( .A(n57), .ZN(n55) );
  NOR2_X1 U101 ( .A1(A[13]), .A2(B[13]), .ZN(n58) );
  OAI21_X1 U102 ( .B1(net22654), .B2(n58), .A(net22627), .ZN(net22651) );
  NAND2_X1 U103 ( .A1(B[12]), .A2(A[12]), .ZN(net22626) );
  OR2_X1 U104 ( .A1(n67), .A2(n71), .ZN(n70) );
  NOR2_X1 U105 ( .A1(n65), .A2(n64), .ZN(n71) );
  INV_X1 U106 ( .A(A[3]), .ZN(n64) );
  NAND2_X1 U107 ( .A1(n64), .A2(n65), .ZN(n68) );
  INV_X1 U108 ( .A(B[3]), .ZN(n65) );
  INV_X1 U109 ( .A(n65), .ZN(net37898) );
  NOR2_X1 U110 ( .A1(net37442), .A2(n66), .ZN(n67) );
  NOR2_X1 U111 ( .A1(A[3]), .A2(B[3]), .ZN(n66) );
  AND2_X1 U112 ( .A1(net37469), .A2(n68), .ZN(n69) );
  NAND2_X1 U113 ( .A1(net35056), .A2(net34775), .ZN(net37469) );
  AND2_X1 U114 ( .A1(net35302), .A2(net37430), .ZN(net37480) );
  NAND4_X1 U115 ( .A1(net22458), .A2(net22452), .A3(net22444), .A4(net35187), 
        .ZN(net22634) );
  BUF_X1 U116 ( .A(net22446), .Z(net35187) );
  AOI21_X1 U117 ( .B1(net35187), .B2(n62), .A(n63), .ZN(n59) );
  NAND2_X1 U118 ( .A1(net35187), .A2(net22447), .ZN(net22440) );
  AND2_X1 U119 ( .A1(n60), .A2(n59), .ZN(net35350) );
  CLKBUF_X1 U120 ( .A(net35350), .Z(net37569) );
  INV_X1 U121 ( .A(net22447), .ZN(n63) );
  INV_X1 U122 ( .A(net22443), .ZN(n62) );
  NAND3_X1 U123 ( .A1(n61), .A2(net22452), .A3(n72), .ZN(n60) );
  AND2_X1 U124 ( .A1(net22446), .A2(net22444), .ZN(n72) );
  NAND2_X1 U125 ( .A1(net22451), .A2(net22456), .ZN(n61) );
  CLKBUF_X1 U126 ( .A(A[3]), .Z(net38443) );
  CLKBUF_X1 U127 ( .A(net37442), .Z(net37487) );
  CLKBUF_X1 U128 ( .A(net35056), .Z(net38135) );
  AND4_X1 U129 ( .A1(net22669), .A2(net22670), .A3(n75), .A4(net22439), .ZN(
        net35345) );
  INV_X1 U130 ( .A(net35345), .ZN(net22643) );
  CLKBUF_X1 U131 ( .A(net22434), .Z(n75) );
  NAND2_X1 U132 ( .A1(n75), .A2(net38589), .ZN(net22432) );
  AOI21_X1 U133 ( .B1(net22670), .B2(n73), .A(net35304), .ZN(net22666) );
  CLKBUF_X1 U134 ( .A(net22666), .Z(net35293) );
  OAI21_X1 U135 ( .B1(n74), .B2(net22438), .A(net22435), .ZN(n73) );
  INV_X1 U136 ( .A(net22434), .ZN(n74) );
  NAND2_X1 U137 ( .A1(B[11]), .A2(A[11]), .ZN(net22668) );
  NAND2_X1 U138 ( .A1(net22668), .A2(net22669), .ZN(net22678) );
  OR2_X1 U139 ( .A1(B[11]), .A2(A[11]), .ZN(net22669) );
  INV_X1 U140 ( .A(B[0]), .ZN(n78) );
  CLKBUF_X1 U141 ( .A(net22435), .Z(net38589) );
  OR2_X1 U142 ( .A1(B[5]), .A2(A[5]), .ZN(net22452) );
  CLKBUF_X1 U143 ( .A(net37430), .Z(net38489) );
  CLKBUF_X1 U144 ( .A(A[6]), .Z(n76) );
  XNOR2_X1 U145 ( .A(net34383), .B(net38371), .ZN(SUM[30]) );
  INV_X1 U146 ( .A(net22488), .ZN(net38298) );
  OR2_X1 U147 ( .A1(B[9]), .A2(A[9]), .ZN(net22434) );
  BUF_X1 U148 ( .A(B[13]), .Z(net35051) );
  AND2_X1 U149 ( .A1(B[10]), .A2(A[10]), .ZN(net35304) );
  NAND2_X1 U150 ( .A1(net22488), .A2(net38489), .ZN(net22485) );
  CLKBUF_X1 U151 ( .A(net22438), .Z(net38162) );
  INV_X1 U152 ( .A(B[2]), .ZN(n79) );
  NAND2_X1 U153 ( .A1(n81), .A2(n82), .ZN(net37430) );
  INV_X1 U154 ( .A(A[0]), .ZN(n77) );
  NAND2_X1 U155 ( .A1(A[0]), .A2(B[0]), .ZN(net34775) );
  NAND2_X1 U156 ( .A1(A[2]), .A2(B[2]), .ZN(net37442) );
  OAI21_X1 U157 ( .B1(net22462), .B2(net22463), .A(net37487), .ZN(net22461) );
  NAND2_X1 U158 ( .A1(net35151), .A2(net37487), .ZN(net22484) );
  XNOR2_X1 U159 ( .A(net37898), .B(net38443), .ZN(net22460) );
  INV_X1 U160 ( .A(B[1]), .ZN(n81) );
  NAND2_X1 U161 ( .A1(B[1]), .A2(A[1]), .ZN(net35056) );
  INV_X1 U162 ( .A(A[2]), .ZN(n80) );
  NAND2_X1 U163 ( .A1(net38135), .A2(net38489), .ZN(net22593) );
  NAND2_X1 U164 ( .A1(n79), .A2(n80), .ZN(net35302) );
  INV_X1 U165 ( .A(A[1]), .ZN(n82) );
  OAI21_X1 U166 ( .B1(n74), .B2(net22684), .A(net38589), .ZN(net22682) );
  CLKBUF_X1 U167 ( .A(net22451), .Z(net35340) );
  INV_X1 U168 ( .A(net35304), .ZN(net22673) );
  CLKBUF_X1 U169 ( .A(n120), .Z(n83) );
  INV_X1 U170 ( .A(net22463), .ZN(net35151) );
  CLKBUF_X1 U171 ( .A(A[13]), .Z(net34908) );
  OAI21_X1 U172 ( .B1(net34874), .B2(n119), .A(n83), .ZN(n84) );
  OR2_X1 U173 ( .A1(A[6]), .A2(B[6]), .ZN(net22444) );
  CLKBUF_X1 U174 ( .A(net22577), .Z(net34874) );
  CLKBUF_X1 U175 ( .A(net22456), .Z(net34451) );
  XOR2_X1 U176 ( .A(net22535), .B(net22537), .Z(SUM[24]) );
  INV_X1 U177 ( .A(net34775), .ZN(net22488) );
  INV_X1 U178 ( .A(net34345), .ZN(net22457) );
  INV_X1 U179 ( .A(net34787), .ZN(net22491) );
  XNOR2_X1 U180 ( .A(n141), .B(n140), .ZN(SUM[17]) );
  NAND2_X1 U181 ( .A1(n131), .A2(n132), .ZN(n141) );
  XNOR2_X1 U182 ( .A(net22530), .B(net22529), .ZN(SUM[25]) );
  XNOR2_X1 U183 ( .A(n114), .B(n113), .ZN(SUM[21]) );
  NAND2_X1 U184 ( .A1(n104), .A2(n105), .ZN(n114) );
  XNOR2_X1 U185 ( .A(n6), .B(net22525), .ZN(SUM[26]) );
  XNOR2_X1 U186 ( .A(n138), .B(n137), .ZN(SUM[18]) );
  NAND2_X1 U187 ( .A1(n124), .A2(n127), .ZN(n138) );
  XNOR2_X1 U188 ( .A(n134), .B(n135), .ZN(SUM[19]) );
  NAND2_X1 U189 ( .A1(n133), .A2(n126), .ZN(n135) );
  XOR2_X1 U190 ( .A(n117), .B(n118), .Z(SUM[20]) );
  XNOR2_X1 U191 ( .A(net22646), .B(net22647), .ZN(SUM[15]) );
  OAI21_X1 U192 ( .B1(n91), .B2(net22450), .A(net35340), .ZN(n89) );
  XNOR2_X1 U193 ( .A(net22593), .B(net22488), .ZN(SUM[1]) );
  AOI21_X1 U194 ( .B1(n100), .B2(n109), .A(n110), .ZN(n107) );
  NOR2_X1 U195 ( .A1(n96), .A2(n85), .ZN(net22542) );
  AOI21_X1 U196 ( .B1(n97), .B2(n98), .A(n99), .ZN(n96) );
  OAI21_X1 U197 ( .B1(net22577), .B2(n119), .A(n120), .ZN(n115) );
  NOR2_X1 U198 ( .A1(n122), .A2(n121), .ZN(n120) );
  NAND2_X1 U199 ( .A1(n94), .A2(net34451), .ZN(n92) );
  NAND2_X1 U200 ( .A1(net22457), .A2(net22458), .ZN(n94) );
  NAND2_X1 U201 ( .A1(net34951), .A2(n103), .ZN(n113) );
  NAND2_X1 U202 ( .A1(net34874), .A2(n130), .ZN(n140) );
  NAND2_X1 U203 ( .A1(net22485), .A2(net38135), .ZN(net22465) );
  NAND2_X1 U204 ( .A1(n139), .A2(n131), .ZN(n137) );
  NAND2_X1 U205 ( .A1(n132), .A2(n140), .ZN(n139) );
  NAND2_X1 U206 ( .A1(n112), .A2(n104), .ZN(n109) );
  NAND2_X1 U207 ( .A1(n105), .A2(n113), .ZN(n112) );
  NAND2_X1 U208 ( .A1(n149), .A2(net38162), .ZN(net22433) );
  NAND2_X1 U209 ( .A1(net22437), .A2(net22439), .ZN(n149) );
  NAND2_X1 U210 ( .A1(n143), .A2(net22626), .ZN(net22655) );
  NAND2_X1 U211 ( .A1(n144), .A2(net22636), .ZN(n143) );
  XNOR2_X1 U212 ( .A(net22658), .B(net22655), .ZN(SUM[13]) );
  XNOR2_X1 U213 ( .A(n145), .B(n144), .ZN(SUM[12]) );
  NAND2_X1 U214 ( .A1(net22626), .A2(net22636), .ZN(n145) );
  XNOR2_X1 U215 ( .A(net22653), .B(net22651), .ZN(SUM[14]) );
  XNOR2_X1 U216 ( .A(n1), .B(net31956), .ZN(SUM[28]) );
  XNOR2_X1 U217 ( .A(n95), .B(net22457), .ZN(SUM[4]) );
  NAND2_X1 U218 ( .A1(net34451), .A2(net22458), .ZN(n95) );
  XNOR2_X1 U219 ( .A(n86), .B(n8), .ZN(SUM[8]) );
  NAND2_X1 U220 ( .A1(net38162), .A2(net22439), .ZN(n86) );
  XNOR2_X1 U221 ( .A(net22440), .B(n87), .ZN(SUM[7]) );
  NAND2_X1 U222 ( .A1(n88), .A2(net22443), .ZN(n87) );
  NAND2_X1 U223 ( .A1(net22444), .A2(n89), .ZN(n88) );
  XNOR2_X1 U224 ( .A(net22484), .B(net22465), .ZN(SUM[2]) );
  XNOR2_X1 U225 ( .A(n90), .B(n89), .ZN(SUM[6]) );
  NAND2_X1 U226 ( .A1(net22444), .A2(net22443), .ZN(n90) );
  XNOR2_X1 U227 ( .A(n146), .B(net22678), .ZN(SUM[11]) );
  NAND2_X1 U228 ( .A1(net22673), .A2(n147), .ZN(n146) );
  NAND2_X1 U229 ( .A1(net22682), .A2(net22670), .ZN(n147) );
  XNOR2_X1 U230 ( .A(n148), .B(net22682), .ZN(SUM[10]) );
  NAND2_X1 U231 ( .A1(net22673), .A2(net22670), .ZN(n148) );
  XNOR2_X1 U232 ( .A(net22460), .B(net22461), .ZN(SUM[3]) );
  XNOR2_X1 U233 ( .A(n93), .B(n92), .ZN(SUM[5]) );
  NAND2_X1 U234 ( .A1(net22452), .A2(net35340), .ZN(n93) );
  XNOR2_X1 U235 ( .A(net22490), .B(net22491), .ZN(SUM[29]) );
  XNOR2_X1 U236 ( .A(net22432), .B(net22433), .ZN(SUM[9]) );
  XNOR2_X1 U237 ( .A(n109), .B(n111), .ZN(SUM[22]) );
  NAND2_X1 U238 ( .A1(n98), .A2(n100), .ZN(n111) );
  XNOR2_X1 U239 ( .A(net22518), .B(net22519), .ZN(SUM[27]) );
  XNOR2_X1 U240 ( .A(n107), .B(n108), .ZN(SUM[23]) );
  NOR2_X1 U241 ( .A1(n99), .A2(n85), .ZN(n108) );
  NAND2_X1 U242 ( .A1(n103), .A2(n116), .ZN(n118) );
  AOI21_X1 U243 ( .B1(n123), .B2(n124), .A(n125), .ZN(n122) );
  NAND2_X1 U244 ( .A1(n127), .A2(n128), .ZN(n123) );
  OAI21_X1 U245 ( .B1(n129), .B2(n130), .A(n131), .ZN(n128) );
  NAND2_X1 U246 ( .A1(n130), .A2(net22610), .ZN(n142) );
  NAND2_X1 U247 ( .A1(n124), .A2(n136), .ZN(n134) );
  NAND2_X1 U248 ( .A1(n137), .A2(n127), .ZN(n136) );
  NAND2_X1 U249 ( .A1(n100), .A2(n101), .ZN(n97) );
  OAI21_X1 U250 ( .B1(n102), .B2(n103), .A(n104), .ZN(n101) );
  NAND2_X1 U251 ( .A1(B[25]), .A2(A[25]), .ZN(net22515) );
  NAND2_X1 U252 ( .A1(B[24]), .A2(A[24]), .ZN(net22514) );
  NAND2_X1 U253 ( .A1(B[20]), .A2(A[20]), .ZN(n103) );
  NAND2_X1 U254 ( .A1(B[26]), .A2(A[26]), .ZN(net22509) );
  NAND2_X1 U255 ( .A1(net35051), .A2(net34908), .ZN(net22627) );
  NAND2_X1 U256 ( .A1(B[8]), .A2(A[8]), .ZN(net22438) );
  NAND2_X1 U257 ( .A1(A[5]), .A2(B[5]), .ZN(net22451) );
  NAND2_X1 U258 ( .A1(B[16]), .A2(A[16]), .ZN(n130) );
  NAND2_X1 U259 ( .A1(B[21]), .A2(A[21]), .ZN(n104) );
  NAND2_X1 U260 ( .A1(B[9]), .A2(A[9]), .ZN(net22435) );
  NAND2_X1 U261 ( .A1(B[17]), .A2(A[17]), .ZN(n131) );
  OR2_X1 U262 ( .A1(B[7]), .A2(A[7]), .ZN(net22446) );
  NAND2_X1 U263 ( .A1(B[18]), .A2(A[18]), .ZN(n124) );
  NAND2_X1 U264 ( .A1(B[22]), .A2(A[22]), .ZN(n98) );
  NAND2_X1 U265 ( .A1(B[7]), .A2(A[7]), .ZN(net22447) );
  OR2_X1 U266 ( .A1(B[26]), .A2(A[26]), .ZN(net22511) );
  OR2_X1 U267 ( .A1(B[18]), .A2(A[18]), .ZN(n127) );
  OR2_X1 U268 ( .A1(B[22]), .A2(A[22]), .ZN(n100) );
  NAND2_X1 U269 ( .A1(B[19]), .A2(A[19]), .ZN(n133) );
  OR2_X1 U270 ( .A1(B[8]), .A2(A[8]), .ZN(net22439) );
  OR2_X1 U271 ( .A1(B[25]), .A2(A[25]), .ZN(net22516) );
  AND2_X1 U272 ( .A1(B[27]), .A2(A[27]), .ZN(net31820) );
  AND2_X1 U273 ( .A1(B[23]), .A2(A[23]), .ZN(n85) );
  OR2_X1 U274 ( .A1(A[21]), .A2(B[21]), .ZN(n105) );
  OR2_X1 U275 ( .A1(B[17]), .A2(A[17]), .ZN(n132) );
  OR2_X1 U276 ( .A1(A[4]), .A2(B[4]), .ZN(net22458) );
  OR2_X1 U277 ( .A1(B[19]), .A2(A[19]), .ZN(n126) );
  OR2_X1 U278 ( .A1(B[24]), .A2(A[24]), .ZN(net22532) );
  OR2_X1 U279 ( .A1(B[20]), .A2(A[20]), .ZN(n116) );
  OR2_X1 U280 ( .A1(B[12]), .A2(A[12]), .ZN(net22636) );
  OR2_X1 U281 ( .A1(B[16]), .A2(A[16]), .ZN(net22610) );
  OR2_X1 U282 ( .A1(B[27]), .A2(A[27]), .ZN(net22517) );
  OR2_X1 U283 ( .A1(B[23]), .A2(A[23]), .ZN(n106) );
  NAND2_X1 U284 ( .A1(n76), .A2(B[6]), .ZN(net22443) );
  NAND2_X1 U285 ( .A1(B[4]), .A2(A[4]), .ZN(net22456) );
  INV_X1 U286 ( .A(net22452), .ZN(net22450) );
  INV_X1 U287 ( .A(n92), .ZN(n91) );
  INV_X1 U288 ( .A(net22465), .ZN(net22462) );
  INV_X1 U289 ( .A(net34346), .ZN(net22535) );
  INV_X1 U290 ( .A(n105), .ZN(n102) );
  NAND3_X1 U291 ( .A1(n100), .A2(n106), .A3(n105), .ZN(net22541) );
  INV_X1 U292 ( .A(n106), .ZN(n99) );
  INV_X1 U293 ( .A(n98), .ZN(n110) );
  INV_X1 U294 ( .A(n84), .ZN(n117) );
  INV_X1 U295 ( .A(n126), .ZN(n125) );
  INV_X1 U296 ( .A(n132), .ZN(n129) );
  INV_X1 U297 ( .A(n133), .ZN(n121) );
  NAND3_X1 U298 ( .A1(n127), .A2(n126), .A3(n132), .ZN(n119) );
  XNOR2_X1 U299 ( .A(n142), .B(net34452), .ZN(SUM[16]) );
  INV_X1 U300 ( .A(net22655), .ZN(net22654) );
  INV_X1 U301 ( .A(net34831), .ZN(net22665) );
  INV_X1 U302 ( .A(net22437), .ZN(net22664) );
  INV_X1 U303 ( .A(net22433), .ZN(net22684) );
  INV_X1 U304 ( .A(net35302), .ZN(net22463) );
endmodule


module ALU_DATA_W32 ( .FUNC({\FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), A, 
        B, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   N19, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N794, N795, N796, n121, n123, n127, n131, n136, n146, n148,
         n150, n151, n157, n159, n162, n163, n170, n172, n175, n176, n183,
         n184, n186, n192, n195, n196, n197, n198, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n213, n214, n217, n220, n232,
         n247, n253, n254, n258, n259, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n279, n285, n295, n302, n338, n339, n378,
         n401, n402, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n454, n455, n465, n474, n480, n482, n483, n484,
         n485, n487, n488, n489, n496, n497, n503, n504, n506, n507, n508,
         n509, n512, n513, n518, n519, n520, n521, n522, n523, n524, n527,
         n528, n529, n530, n534, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n547, n549, n550, n551, n552, n553, net18425,
         net18434, net18459, net18461, net19990, net19993, net20016, net20298,
         net24439, net24440, net24456, net24457, net24458, net24463, net24464,
         net24465, net24497, net24555, net24560, net24561, net24562, net24726,
         net24728, net24759, net24772, net24773, net24777, net24891, net24901,
         net24911, net26397, net26387, net26385, net26383, net26407, net26403,
         net26415, net26425, net26423, net26437, net26435, net26433, net26431,
         net26459, net26457, net26455, net26453, net26451, net26449, net26445,
         net26473, net26469, net26467, net26465, net26463, net26461, net26485,
         net26483, net26479, net26495, net26493, net26491, net26501, net26499,
         net26497, net26700, net31345, net31362, net31363, net31364, net31396,
         net31776, net31778, net31788, net32003, net32007, net32250, net32589,
         net34396, net34870, net35295, net35313, net35873, net36181, net36207,
         net36683, net36677, net36652, net36631, net36523, net34274, net34273,
         net31775, net24442, n239, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n19, n20, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n122, n124, n125, n126, n128, n129, n130, n132, n133, n134, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n147, n149,
         n152, n153, n154, n155, n156, n158, n160, n161, n164, n165, n166,
         n167, n168, n169, n171, n173, n174, n177, n178, n179, n180, n181,
         n182, n185, n187, n188, n189, n190, n191, n193, n194, n199, n200,
         n201, n212, n215, n216, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n233, n234, n235, n236, n237,
         n238, n240, n241, n242, n243, n244, n245, n246, n248, n249, n250,
         n251, n252, n255, n256, n257, n260, n261, n262, n273, n274, n275,
         n276, n277, n278, n280, n281, n282, n283, n284, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n296, n297, n298, n299, n300,
         n301, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n403, n404, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n466, n467, n468, n469, n470, n471, n472, n473, n475, n476,
         n477, n478, n479, n481, n486, n490, n491, n492, n493, n494, n495,
         n498, n499, n500, n501, n502, n505, n510, n511, n514, n515, n516,
         n517, n525, n526, n531, n532, n533, n535, n546, n548, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791;
  wire   [3:0] FUNC;

  NOR2_X2 U458 ( .A1(n762), .A2(n274), .ZN(n213) );
  ALU_DATA_W32_DW01_cmp6_0 r80 ( .A({B[31:14], n158, n23, B[11:10], n166, B[8], 
        n190, n225, n231, n96, n168, n143, n83, n142}), .B({A[31:14], n174, 
        A[12:8], n141, n144, n155, n242, n109, n106, n76, A[0]}), .TC(1'b0), 
        .LE(N794), .GE(N795), .NE(N796) );
  ALU_DATA_W32_DW01_sub_2 sub_128 ( .A({A[31], n77, A[29:27], n154, A[25], 
        n169, A[23:9], n234, A[7:4], n236, n261, A[1], n245}), .B({B[31:27], 
        n75, B[25:19], n32, B[17:10], n226, B[8:3], n82, B[1], n171}), .CI(
        1'b0), .DIFF({N122, N121, N120, N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91}) );
  ALU_DATA_W32_DW01_add_2 add_125 ( .A({A[31], n77, A[29:27], n154, A[25], 
        n169, A[23:15], n173, A[13:11], net34396, A[9], n234, A[7:5], n161, 
        n72, n149, A[1], n275}), .B({B[31:27], n31, B[25:19], n32, B[17:15], 
        n156, B[13:12], n108, B[10:9], n228, B[7:6], n107, n178, B[3], n82, 
        n187, n171}), .CI(1'b0), .SUM({N90, N89, N88, N87, N86, N85, N84, N83, 
        N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, N66, N65, N64, N63, N62, N61, N60, N59}) );
  AND3_X1 U3 ( .A1(n1), .A2(n2), .A3(n3), .ZN(n689) );
  NAND2_X1 U4 ( .A1(N86), .A2(net26491), .ZN(n1) );
  NAND2_X1 U6 ( .A1(n255), .A2(net24465), .ZN(n2) );
  NAND2_X1 U7 ( .A1(N118), .A2(net26499), .ZN(n3) );
  NOR2_X1 U8 ( .A1(net18459), .A2(n133), .ZN(n120) );
  INV_X1 U9 ( .A(net24465), .ZN(n124) );
  NOR2_X1 U10 ( .A1(net26700), .A2(net36631), .ZN(n125) );
  NAND2_X1 U12 ( .A1(n61), .A2(n62), .ZN(n59) );
  NAND2_X1 U13 ( .A1(net24456), .A2(n213), .ZN(n61) );
  NAND2_X1 U15 ( .A1(net24457), .A2(n232), .ZN(n62) );
  NOR2_X1 U16 ( .A1(net26700), .A2(n51), .ZN(n52) );
  INV_X1 U17 ( .A(net24458), .ZN(n51) );
  INV_X1 U18 ( .A(net24773), .ZN(n129) );
  NAND2_X1 U19 ( .A1(net35295), .A2(net24772), .ZN(n128) );
  BUF_X1 U20 ( .A(B[2]), .Z(n82) );
  BUF_X1 U21 ( .A(A[8]), .Z(n234) );
  NAND2_X1 U22 ( .A1(net26455), .A2(A[29]), .ZN(n114) );
  AND3_X1 U23 ( .A1(n483), .A2(n548), .A3(n491), .ZN(n47) );
  AND3_X1 U24 ( .A1(n521), .A2(n568), .A3(n505), .ZN(n46) );
  INV_X1 U25 ( .A(A[29]), .ZN(net19993) );
  BUF_X1 U26 ( .A(B[3]), .Z(n168) );
  NAND2_X1 U27 ( .A1(n115), .A2(n214), .ZN(n163) );
  NOR2_X1 U28 ( .A1(n120), .A2(n122), .ZN(n115) );
  INV_X1 U29 ( .A(n84), .ZN(n381) );
  INV_X1 U30 ( .A(n47), .ZN(n472) );
  BUF_X1 U31 ( .A(n174), .Z(n238) );
  INV_X1 U32 ( .A(n46), .ZN(n498) );
  OAI222_X1 U33 ( .A1(n393), .A2(net26700), .B1(net26479), .B2(n715), .C1(n342), .C2(net24561), .ZN(n653) );
  NAND2_X1 U34 ( .A1(n213), .A2(net24464), .ZN(n112) );
  NAND2_X1 U35 ( .A1(net36677), .A2(net24463), .ZN(n111) );
  NAND2_X1 U36 ( .A1(net24562), .A2(net26485), .ZN(net36523) );
  AOI211_X1 U37 ( .C1(n58), .C2(net26483), .A(n59), .B(n52), .ZN(n57) );
  NAND4_X1 U38 ( .A1(net36683), .A2(n4), .A3(n8), .A4(net24439), .ZN(n58) );
  INV_X1 U39 ( .A(net24439), .ZN(n50) );
  NOR2_X1 U40 ( .A1(A[31]), .A2(net26387), .ZN(n53) );
  BUF_X1 U41 ( .A(A[2]), .Z(n149) );
  INV_X1 U42 ( .A(n48), .ZN(n399) );
  NOR2_X1 U43 ( .A1(net24439), .A2(n118), .ZN(n116) );
  NAND2_X1 U44 ( .A1(n128), .A2(n129), .ZN(n117) );
  INV_X1 U45 ( .A(net32250), .ZN(n118) );
  AOI222_X1 U46 ( .A1(n255), .A2(n606), .B1(n256), .B2(n605), .C1(n257), .C2(
        n604), .ZN(n608) );
  AOI221_X1 U47 ( .B1(n250), .B2(net24464), .C1(n251), .C2(net24463), .A(n613), 
        .ZN(n625) );
  AOI221_X1 U48 ( .B1(n246), .B2(n699), .C1(n257), .C2(n636), .A(n635), .ZN(
        n642) );
  AOI221_X1 U49 ( .B1(n678), .B2(n662), .C1(n75), .C2(n661), .A(n660), .ZN(
        n674) );
  INV_X1 U50 ( .A(net26449), .ZN(n134) );
  OR2_X1 U51 ( .A1(net32589), .A2(n119), .ZN(n4) );
  INV_X1 U52 ( .A(net26437), .ZN(n133) );
  AND2_X1 U53 ( .A1(net31362), .A2(net31396), .ZN(n5) );
  AND3_X1 U54 ( .A1(n99), .A2(n100), .A3(n101), .ZN(n6) );
  BUF_X1 U55 ( .A(B[1]), .Z(n83) );
  OR3_X1 U56 ( .A1(B[31]), .A2(B[30]), .A3(n231), .ZN(n7) );
  OR2_X1 U57 ( .A1(net32007), .A2(net19990), .ZN(n8) );
  OR2_X1 U58 ( .A1(B[25]), .A2(B[23]), .ZN(n9) );
  OR2_X1 U59 ( .A1(B[18]), .A2(B[16]), .ZN(n10) );
  BUF_X1 U60 ( .A(A[3]), .Z(n109) );
  AND2_X1 U61 ( .A1(n676), .A2(n675), .ZN(n11) );
  AND2_X1 U62 ( .A1(n759), .A2(FUNC[1]), .ZN(n12) );
  AND2_X1 U63 ( .A1(n758), .A2(FUNC[3]), .ZN(n13) );
  AND2_X1 U64 ( .A1(n54), .A2(n65), .ZN(n14) );
  AND2_X1 U65 ( .A1(n11), .A2(n710), .ZN(n15) );
  OR2_X1 U66 ( .A1(n791), .A2(n273), .ZN(n16) );
  OR2_X1 U67 ( .A1(n791), .A2(n273), .ZN(n19) );
  AND3_X2 U68 ( .A1(n520), .A2(n632), .A3(n600), .ZN(n20) );
  OR2_X1 U69 ( .A1(n791), .A2(n273), .ZN(n104) );
  AND2_X1 U70 ( .A1(n78), .A2(n5), .ZN(n22) );
  CLKBUF_X1 U71 ( .A(A[4]), .Z(n161) );
  CLKBUF_X1 U72 ( .A(A[4]), .Z(n242) );
  CLKBUF_X1 U73 ( .A(B[12]), .Z(n23) );
  NAND2_X1 U74 ( .A1(B[0]), .A2(n240), .ZN(net32007) );
  INV_X1 U75 ( .A(n585), .ZN(n24) );
  NOR2_X1 U76 ( .A1(n116), .A2(n117), .ZN(net24759) );
  AND2_X1 U77 ( .A1(n623), .A2(n625), .ZN(n25) );
  NAND2_X1 U78 ( .A1(N81), .A2(net26491), .ZN(n26) );
  NAND2_X1 U79 ( .A1(n212), .A2(n732), .ZN(n27) );
  NAND2_X1 U80 ( .A1(N113), .A2(net26501), .ZN(n28) );
  AND3_X1 U81 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n607) );
  BUF_X1 U82 ( .A(n68), .Z(net26501) );
  AND2_X1 U83 ( .A1(n22), .A2(n213), .ZN(n29) );
  INV_X1 U84 ( .A(n168), .ZN(n30) );
  INV_X1 U85 ( .A(n168), .ZN(n762) );
  CLKBUF_X1 U86 ( .A(B[26]), .Z(n31) );
  BUF_X1 U87 ( .A(B[18]), .Z(n32) );
  AND3_X1 U88 ( .A1(n88), .A2(n89), .A3(n90), .ZN(n622) );
  BUF_X1 U89 ( .A(B[4]), .Z(n178) );
  INV_X1 U90 ( .A(n649), .ZN(n33) );
  CLKBUF_X1 U91 ( .A(A[2]), .Z(n106) );
  BUF_X1 U92 ( .A(B[1]), .Z(n187) );
  INV_X1 U93 ( .A(n450), .ZN(n34) );
  AND2_X1 U94 ( .A1(N78), .A2(net26493), .ZN(n35) );
  AND2_X1 U95 ( .A1(n687), .A2(net24465), .ZN(n36) );
  AND2_X1 U96 ( .A1(N110), .A2(net26501), .ZN(n37) );
  NOR3_X1 U97 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n558) );
  BUF_X1 U98 ( .A(net31775), .Z(net26493) );
  AOI221_X4 U99 ( .B1(n154), .B2(net26423), .C1(A[27]), .C2(net26435), .A(n285), .ZN(n279) );
  CLKBUF_X3 U100 ( .A(A[26]), .Z(n154) );
  CLKBUF_X1 U101 ( .A(n225), .Z(n38) );
  BUF_X1 U102 ( .A(B[6]), .Z(n225) );
  NOR3_X1 U103 ( .A1(n766), .A2(n91), .A3(n10), .ZN(n771) );
  AOI221_X4 U104 ( .B1(n33), .B2(net36207), .C1(n154), .C2(net26437), .A(n302), 
        .ZN(n295) );
  AND2_X2 U105 ( .A1(n678), .A2(net26483), .ZN(n251) );
  NAND3_X1 U106 ( .A1(n15), .A2(n709), .A3(n708), .ZN(RES[28]) );
  INV_X1 U107 ( .A(net32589), .ZN(n39) );
  INV_X1 U108 ( .A(net32589), .ZN(n40) );
  OR2_X1 U109 ( .A1(n19), .A2(net24891), .ZN(n41) );
  NAND2_X1 U110 ( .A1(n41), .A2(net24901), .ZN(n390) );
  NAND2_X2 U111 ( .A1(n273), .A2(n276), .ZN(net32589) );
  CLKBUF_X1 U112 ( .A(net32589), .Z(net26461) );
  INV_X1 U113 ( .A(n60), .ZN(n64) );
  INV_X1 U114 ( .A(net24562), .ZN(net36631) );
  AOI221_X1 U115 ( .B1(n257), .B2(n408), .C1(n256), .C2(n102), .A(n481), .ZN(
        n494) );
  NAND2_X1 U116 ( .A1(N121), .A2(net26499), .ZN(n42) );
  NAND2_X1 U117 ( .A1(N89), .A2(net26491), .ZN(n43) );
  INV_X1 U118 ( .A(n753), .ZN(n44) );
  AND3_X1 U119 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n754) );
  INV_X1 U120 ( .A(n78), .ZN(n436) );
  CLKBUF_X1 U121 ( .A(n78), .Z(n189) );
  NAND3_X1 U122 ( .A1(n622), .A2(n624), .A3(n25), .ZN(RES[23]) );
  AOI221_X4 U123 ( .B1(n687), .B2(net24457), .C1(n246), .C2(net24456), .A(n619), .ZN(n624) );
  CLKBUF_X1 U124 ( .A(n347), .Z(n45) );
  INV_X1 U125 ( .A(n16), .ZN(net26437) );
  INV_X1 U126 ( .A(net32007), .ZN(net26425) );
  AND3_X2 U127 ( .A1(n484), .A2(n615), .A3(n583), .ZN(n48) );
  AOI22_X1 U128 ( .A1(n445), .A2(net36677), .B1(net26485), .B2(n526), .ZN(n49)
         );
  INV_X1 U129 ( .A(net26700), .ZN(net36677) );
  NAND2_X1 U130 ( .A1(net24464), .A2(n232), .ZN(n132) );
  NAND2_X1 U131 ( .A1(N122), .A2(n68), .ZN(n69) );
  NAND2_X1 U132 ( .A1(net24442), .A2(n14), .ZN(RES[31]) );
  AND2_X1 U133 ( .A1(n56), .A2(n55), .ZN(n65) );
  OAI21_X1 U134 ( .B1(n53), .B2(net31788), .A(B[31]), .ZN(n55) );
  INV_X1 U135 ( .A(net26397), .ZN(net26387) );
  MUX2_X1 U136 ( .A(net26397), .B(net31778), .S(B[29]), .Z(net24497) );
  INV_X1 U137 ( .A(net26397), .ZN(net26385) );
  NAND2_X1 U138 ( .A1(n63), .A2(n50), .ZN(n56) );
  INV_X1 U139 ( .A(net24440), .ZN(n63) );
  NAND2_X1 U140 ( .A1(n64), .A2(net32003), .ZN(n54) );
  MUX2_X1 U141 ( .A(net36652), .B(n57), .S(net35873), .Z(n60) );
  BUF_X1 U142 ( .A(n210), .Z(net35873) );
  AND3_X1 U143 ( .A1(n69), .A2(net34273), .A3(net34274), .ZN(net24442) );
  NAND2_X1 U144 ( .A1(A[31]), .A2(n66), .ZN(net34274) );
  NAND3_X1 U145 ( .A1(n239), .A2(net26403), .A3(n67), .ZN(n66) );
  MUX2_X1 U146 ( .A(net26387), .B(net26415), .S(B[31]), .Z(n67) );
  NAND2_X1 U147 ( .A1(N90), .A2(net26493), .ZN(net34273) );
  NAND2_X1 U148 ( .A1(net31362), .A2(net31345), .ZN(n239) );
  NOR2_X1 U149 ( .A1(n239), .A2(N19), .ZN(n208) );
  AND2_X1 U150 ( .A1(n411), .A2(n239), .ZN(n524) );
  INV_X1 U151 ( .A(n239), .ZN(net24726) );
  AND2_X1 U152 ( .A1(net31776), .A2(net31345), .ZN(net31778) );
  NAND2_X1 U153 ( .A1(net31364), .A2(net31396), .ZN(n123) );
  AND2_X1 U154 ( .A1(net31363), .A2(net31345), .ZN(net31788) );
  AND2_X1 U155 ( .A1(net31776), .A2(net31396), .ZN(net31775) );
  BUF_X1 U156 ( .A(net31775), .Z(net26491) );
  BUF_X1 U157 ( .A(net31775), .Z(net26495) );
  AND2_X1 U158 ( .A1(net31363), .A2(net31396), .ZN(n68) );
  BUF_X1 U159 ( .A(n68), .Z(net26499) );
  BUF_X1 U160 ( .A(n68), .Z(net26497) );
  OR2_X1 U161 ( .A1(net18434), .A2(n752), .ZN(n70) );
  NAND2_X1 U162 ( .A1(n70), .A2(n6), .ZN(n266) );
  CLKBUF_X1 U163 ( .A(n568), .Z(n71) );
  BUF_X1 U164 ( .A(A[0]), .Z(n245) );
  CLKBUF_X1 U165 ( .A(B[12]), .Z(n200) );
  NOR2_X1 U166 ( .A1(net32007), .A2(net18461), .ZN(n122) );
  BUF_X1 U167 ( .A(B[13]), .Z(n158) );
  BUF_X1 U168 ( .A(B[2]), .Z(n143) );
  BUF_X1 U169 ( .A(A[3]), .Z(n72) );
  CLKBUF_X1 U170 ( .A(B[15]), .Z(n73) );
  CLKBUF_X1 U171 ( .A(n205), .Z(n74) );
  AOI221_X1 U172 ( .B1(n241), .B2(net36181), .C1(n177), .C2(net26437), .A(n272), .ZN(n271) );
  AOI221_X1 U173 ( .B1(n244), .B2(net36207), .C1(n241), .C2(net26437), .A(n220), .ZN(n217) );
  CLKBUF_X1 U174 ( .A(n31), .Z(n75) );
  BUF_X1 U175 ( .A(A[3]), .Z(n236) );
  BUF_X1 U176 ( .A(A[1]), .Z(n76) );
  BUF_X1 U177 ( .A(B[11]), .Z(n108) );
  INV_X1 U178 ( .A(n119), .ZN(n77) );
  INV_X1 U179 ( .A(A[30]), .ZN(n119) );
  AND2_X2 U180 ( .A1(n210), .A2(net34870), .ZN(n78) );
  NAND2_X1 U181 ( .A1(N83), .A2(net26491), .ZN(n79) );
  NAND2_X1 U182 ( .A1(n29), .A2(n639), .ZN(n80) );
  NAND2_X1 U183 ( .A1(N115), .A2(net26499), .ZN(n81) );
  AND3_X1 U184 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n640) );
  BUF_X2 U185 ( .A(B[14]), .Z(n156) );
  AND2_X2 U186 ( .A1(net24726), .A2(net20016), .ZN(n84) );
  AOI221_X4 U187 ( .B1(n84), .B2(n652), .C1(n131), .C2(n645), .A(n341), .ZN(
        n346) );
  INV_X1 U188 ( .A(n210), .ZN(net20016) );
  BUF_X1 U189 ( .A(A[0]), .Z(n275) );
  AND2_X1 U190 ( .A1(n444), .A2(n397), .ZN(n85) );
  AND2_X1 U191 ( .A1(n22), .A2(n653), .ZN(n86) );
  AND2_X1 U192 ( .A1(n252), .A2(n472), .ZN(n87) );
  NOR3_X1 U193 ( .A1(n85), .A2(n86), .A3(n87), .ZN(n345) );
  AND2_X2 U194 ( .A1(n299), .A2(n213), .ZN(n252) );
  NAND2_X1 U195 ( .A1(N82), .A2(net26491), .ZN(n88) );
  NAND2_X1 U196 ( .A1(n29), .A2(net24465), .ZN(n89) );
  NAND2_X1 U197 ( .A1(N114), .A2(net26499), .ZN(n90) );
  BUF_X1 U198 ( .A(B[9]), .Z(n226) );
  NAND2_X1 U199 ( .A1(n160), .A2(net34870), .ZN(n210) );
  CLKBUF_X1 U200 ( .A(B[17]), .Z(n91) );
  AND2_X1 U201 ( .A1(n256), .A2(n670), .ZN(n92) );
  AND2_X1 U202 ( .A1(n687), .A2(n739), .ZN(n93) );
  AND2_X1 U203 ( .A1(n29), .A2(n738), .ZN(n94) );
  NOR3_X1 U204 ( .A1(n92), .A2(n93), .A3(n94), .ZN(n672) );
  INV_X1 U205 ( .A(net18461), .ZN(n95) );
  CLKBUF_X1 U206 ( .A(A[10]), .Z(net34396) );
  BUF_X1 U207 ( .A(B[4]), .Z(n96) );
  NAND2_X1 U208 ( .A1(n676), .A2(n675), .ZN(n97) );
  NOR2_X1 U209 ( .A1(n768), .A2(n7), .ZN(n769) );
  BUF_X1 U210 ( .A(B[5]), .Z(n231) );
  CLKBUF_X1 U211 ( .A(B[7]), .Z(n190) );
  OAI221_X1 U212 ( .B1(net26463), .B2(n786), .C1(net26445), .C2(n787), .A(n414), .ZN(n186) );
  OAI22_X1 U213 ( .A1(net26463), .A2(net19993), .B1(net19990), .B2(n133), .ZN(
        n253) );
  OR2_X1 U214 ( .A1(net18434), .A2(n746), .ZN(n98) );
  NAND2_X1 U215 ( .A1(n98), .A2(n6), .ZN(n267) );
  OR2_X1 U216 ( .A1(n499), .A2(net24561), .ZN(n99) );
  OR2_X1 U217 ( .A1(net26479), .A2(n46), .ZN(n100) );
  OR2_X1 U218 ( .A1(n20), .A2(net26700), .ZN(n101) );
  CLKBUF_X1 U219 ( .A(n409), .Z(n102) );
  CLKBUF_X1 U220 ( .A(B[10]), .Z(n103) );
  AOI221_X4 U221 ( .B1(n257), .B2(n645), .C1(B[25]), .C2(n644), .A(n660), .ZN(
        n657) );
  INV_X1 U222 ( .A(net26461), .ZN(net26469) );
  CLKBUF_X1 U223 ( .A(n32), .Z(n105) );
  INV_X2 U224 ( .A(n213), .ZN(net24561) );
  NAND2_X4 U225 ( .A1(n30), .A2(n181), .ZN(net26479) );
  CLKBUF_X1 U226 ( .A(B[5]), .Z(n107) );
  CLKBUF_X3 U227 ( .A(A[2]), .Z(n261) );
  NOR2_X1 U228 ( .A1(n126), .A2(n125), .ZN(net36652) );
  OAI211_X1 U229 ( .C1(net26479), .C2(n124), .A(n130), .B(n132), .ZN(n126) );
  NAND2_X1 U230 ( .A1(n213), .A2(net24463), .ZN(n130) );
  NAND2_X1 U231 ( .A1(net26433), .A2(A[29]), .ZN(net36683) );
  NAND2_X1 U232 ( .A1(A[30]), .A2(net26467), .ZN(n113) );
  NAND2_X1 U233 ( .A1(n113), .A2(n114), .ZN(n480) );
  CLKBUF_X1 U234 ( .A(A[12]), .Z(n110) );
  INV_X2 U235 ( .A(net31788), .ZN(net26407) );
  NAND3_X1 U236 ( .A1(net36523), .A2(n111), .A3(n112), .ZN(net24555) );
  BUF_X2 U237 ( .A(net26425), .Z(net36181) );
  BUF_X2 U238 ( .A(net26425), .Z(net36207) );
  BUF_X2 U239 ( .A(net26431), .Z(n135) );
  BUF_X1 U240 ( .A(A[17]), .Z(n137) );
  CLKBUF_X1 U241 ( .A(B[9]), .Z(n166) );
  OR2_X2 U242 ( .A1(n464), .A2(net26479), .ZN(n441) );
  AND2_X1 U243 ( .A1(B[30]), .A2(n749), .ZN(n138) );
  AND2_X1 U244 ( .A1(net32003), .A2(n748), .ZN(n139) );
  NOR3_X1 U245 ( .A1(n138), .A2(n139), .A3(n747), .ZN(n755) );
  AOI221_X4 U246 ( .B1(B[20]), .B2(n565), .C1(n564), .C2(n563), .A(n660), .ZN(
        n578) );
  NAND2_X1 U247 ( .A1(n299), .A2(n232), .ZN(n442) );
  OR4_X1 U248 ( .A1(n166), .A2(n38), .A3(n190), .A4(n228), .ZN(n768) );
  AOI21_X1 U249 ( .B1(A[31]), .B2(n187), .A(n480), .ZN(n338) );
  OR2_X1 U250 ( .A1(n338), .A2(n745), .ZN(n140) );
  NAND2_X1 U251 ( .A1(n140), .A2(n11), .ZN(n724) );
  AOI221_X4 U252 ( .B1(n256), .B2(n588), .C1(n248), .C2(n718), .A(n587), .ZN(
        n593) );
  BUF_X1 U253 ( .A(B[8]), .Z(n228) );
  CLKBUF_X1 U254 ( .A(A[7]), .Z(n141) );
  OR2_X2 U255 ( .A1(n296), .A2(net26479), .ZN(n466) );
  CLKBUF_X1 U256 ( .A(B[0]), .Z(n142) );
  CLKBUF_X1 U257 ( .A(A[9]), .Z(net35313) );
  CLKBUF_X1 U258 ( .A(A[6]), .Z(n144) );
  AND2_X1 U259 ( .A1(n29), .A2(net24464), .ZN(n145) );
  AND2_X1 U260 ( .A1(n687), .A2(net24463), .ZN(n147) );
  NOR3_X1 U261 ( .A1(n145), .A2(n147), .A3(n360), .ZN(n368) );
  CLKBUF_X1 U262 ( .A(A[15]), .Z(net35295) );
  OR2_X1 U263 ( .A1(n746), .A2(n745), .ZN(n152) );
  NAND2_X1 U264 ( .A1(n152), .A2(n11), .ZN(n747) );
  BUF_X1 U265 ( .A(n173), .Z(n153) );
  CLKBUF_X1 U266 ( .A(A[14]), .Z(n173) );
  INV_X1 U267 ( .A(n763), .ZN(n274) );
  BUF_X1 U268 ( .A(B[1]), .Z(n240) );
  CLKBUF_X1 U269 ( .A(A[5]), .Z(n155) );
  BUF_X1 U270 ( .A(B[0]), .Z(n171) );
  INV_X1 U271 ( .A(n764), .ZN(n273) );
  INV_X1 U272 ( .A(net34870), .ZN(N19) );
  CLKBUF_X1 U273 ( .A(n178), .Z(n160) );
  AOI221_X4 U274 ( .B1(n678), .B2(net24555), .C1(B[27]), .C2(n677), .A(n97), 
        .ZN(n692) );
  OR4_X1 U275 ( .A1(B[21]), .A2(B[19]), .A3(B[22]), .A4(B[20]), .ZN(n766) );
  CLKBUF_X1 U276 ( .A(A[11]), .Z(n164) );
  CLKBUF_X1 U277 ( .A(n275), .Z(n165) );
  CLKBUF_X1 U278 ( .A(n76), .Z(n260) );
  BUF_X1 U279 ( .A(A[22]), .Z(n167) );
  AOI221_X4 U280 ( .B1(n260), .B2(net31778), .C1(net26397), .C2(n790), .A(
        net31788), .ZN(n405) );
  BUF_X2 U281 ( .A(A[24]), .Z(n169) );
  BUF_X1 U282 ( .A(A[13]), .Z(n174) );
  AOI221_X4 U283 ( .B1(n149), .B2(net31778), .C1(net26397), .C2(n789), .A(
        net31788), .ZN(n263) );
  CLKBUF_X1 U284 ( .A(n161), .Z(n177) );
  INV_X1 U285 ( .A(n166), .ZN(n179) );
  INV_X1 U286 ( .A(n179), .ZN(n180) );
  INV_X1 U287 ( .A(n274), .ZN(n181) );
  AND4_X2 U288 ( .A1(n772), .A2(n769), .A3(n771), .A4(n770), .ZN(net34870) );
  INV_X1 U289 ( .A(n466), .ZN(n182) );
  AND2_X1 U290 ( .A1(n299), .A2(n232), .ZN(n185) );
  OR2_X1 U291 ( .A1(n464), .A2(net26700), .ZN(n363) );
  INV_X1 U292 ( .A(net26700), .ZN(net20298) );
  CLKBUF_X1 U293 ( .A(n185), .Z(n188) );
  CLKBUF_X1 U294 ( .A(n144), .Z(n244) );
  AND2_X1 U295 ( .A1(N96), .A2(net26497), .ZN(n191) );
  AND2_X1 U296 ( .A1(n136), .A2(n444), .ZN(n193) );
  AND2_X1 U297 ( .A1(n186), .A2(n370), .ZN(n194) );
  NOR3_X1 U298 ( .A1(n191), .A2(n193), .A3(n194), .ZN(n309) );
  CLKBUF_X1 U299 ( .A(n444), .Z(n199) );
  CLKBUF_X1 U300 ( .A(n108), .Z(n201) );
  OR2_X1 U301 ( .A1(n296), .A2(net26700), .ZN(n467) );
  INV_X1 U302 ( .A(n424), .ZN(n212) );
  NOR3_X1 U303 ( .A1(n767), .A2(B[24]), .A3(n9), .ZN(n770) );
  AND2_X1 U304 ( .A1(n678), .A2(n653), .ZN(n215) );
  AND2_X1 U305 ( .A1(n256), .A2(n652), .ZN(n216) );
  AND2_X1 U306 ( .A1(n29), .A2(n717), .ZN(n218) );
  NOR3_X1 U307 ( .A1(n215), .A2(n216), .A3(n218), .ZN(n655) );
  AND2_X1 U308 ( .A1(n687), .A2(net24562), .ZN(n219) );
  AND2_X1 U309 ( .A1(n255), .A2(net24464), .ZN(n221) );
  AND2_X1 U310 ( .A1(n29), .A2(net24463), .ZN(n222) );
  NOR3_X1 U311 ( .A1(n219), .A2(n221), .A3(n222), .ZN(n448) );
  CLKBUF_X1 U312 ( .A(B[21]), .Z(n223) );
  INV_X1 U313 ( .A(n441), .ZN(n224) );
  CLKBUF_X1 U314 ( .A(A[8]), .Z(n235) );
  AOI221_X1 U315 ( .B1(n238), .B2(n395), .C1(n255), .C2(n712), .A(n394), .ZN(
        n404) );
  CLKBUF_X1 U316 ( .A(n38), .Z(n227) );
  BUF_X2 U317 ( .A(n467), .Z(n249) );
  CLKBUF_X1 U318 ( .A(n141), .Z(n229) );
  INV_X1 U319 ( .A(n569), .ZN(n230) );
  INV_X1 U320 ( .A(n30), .ZN(n233) );
  CLKBUF_X1 U321 ( .A(n228), .Z(n237) );
  CLKBUF_X1 U322 ( .A(n155), .Z(n241) );
  CLKBUF_X1 U323 ( .A(n236), .Z(n243) );
  NAND2_X1 U324 ( .A1(n551), .A2(n13), .ZN(n529) );
  NAND2_X1 U325 ( .A1(N796), .A2(n12), .ZN(n553) );
  INV_X2 U326 ( .A(n467), .ZN(n687) );
  INV_X1 U327 ( .A(n466), .ZN(n246) );
  INV_X1 U328 ( .A(n466), .ZN(n248) );
  INV_X1 U329 ( .A(n466), .ZN(n686) );
  INV_X2 U330 ( .A(net26467), .ZN(net26463) );
  INV_X1 U331 ( .A(net26449), .ZN(net26445) );
  INV_X1 U332 ( .A(n363), .ZN(n444) );
  INV_X1 U333 ( .A(n441), .ZN(n370) );
  INV_X1 U334 ( .A(n19), .ZN(net26435) );
  INV_X1 U335 ( .A(n104), .ZN(net26431) );
  INV_X1 U336 ( .A(n19), .ZN(net26433) );
  AND2_X1 U337 ( .A1(n678), .A2(net20298), .ZN(n250) );
  BUF_X1 U338 ( .A(net26459), .Z(net26451) );
  BUF_X1 U339 ( .A(net26457), .Z(net26453) );
  BUF_X1 U340 ( .A(net26459), .Z(net26449) );
  BUF_X1 U341 ( .A(net26457), .Z(net26455) );
  INV_X1 U342 ( .A(net26397), .ZN(net26383) );
  INV_X1 U343 ( .A(net32007), .ZN(net26423) );
  OAI22_X1 U344 ( .A1(net26465), .A2(n790), .B1(n133), .B2(n789), .ZN(n542) );
  OAI21_X1 U345 ( .B1(n274), .B2(net26383), .A(net26407), .ZN(n264) );
  AND2_X1 U346 ( .A1(n131), .A2(net26485), .ZN(net32250) );
  INV_X1 U347 ( .A(net32589), .ZN(net26467) );
  INV_X1 U348 ( .A(net26461), .ZN(net26473) );
  AND2_X2 U349 ( .A1(n22), .A2(n232), .ZN(n255) );
  AND2_X2 U350 ( .A1(n78), .A2(net24726), .ZN(n256) );
  AOI22_X1 U351 ( .A1(n408), .A2(n206), .B1(n409), .B2(n208), .ZN(n407) );
  AOI22_X1 U352 ( .A1(n205), .A2(n206), .B1(n207), .B2(n208), .ZN(n204) );
  AOI22_X1 U353 ( .A1(n266), .A2(n206), .B1(n267), .B2(n208), .ZN(n265) );
  INV_X1 U354 ( .A(net18425), .ZN(net26457) );
  INV_X1 U355 ( .A(net18425), .ZN(net26459) );
  NOR2_X1 U356 ( .A1(n411), .A2(N19), .ZN(n206) );
  NOR2_X1 U357 ( .A1(n181), .A2(n762), .ZN(n232) );
  NOR2_X1 U358 ( .A1(n411), .A2(n210), .ZN(n131) );
  OAI221_X1 U359 ( .B1(n268), .B2(n781), .C1(n208), .C2(n206), .A(net35873), 
        .ZN(n258) );
  OAI221_X1 U360 ( .B1(n410), .B2(n782), .C1(n208), .C2(n206), .A(net35873), 
        .ZN(n401) );
  AOI22_X1 U361 ( .A1(net20016), .A2(n775), .B1(n260), .B2(n406), .ZN(n402) );
  AOI22_X1 U362 ( .A1(n176), .A2(net20298), .B1(n175), .B2(n213), .ZN(n269) );
  NOR2_X1 U363 ( .A1(N19), .A2(n524), .ZN(n536) );
  OAI22_X1 U364 ( .A1(n455), .A2(net35873), .B1(net20016), .B2(n539), .ZN(n537) );
  AND2_X1 U365 ( .A1(n5), .A2(net34870), .ZN(net32003) );
  INV_X1 U366 ( .A(n260), .ZN(n790) );
  AND2_X2 U367 ( .A1(n189), .A2(net24728), .ZN(n257) );
  AOI22_X1 U368 ( .A1(n186), .A2(net20298), .B1(n136), .B2(n213), .ZN(n412) );
  AOI22_X1 U369 ( .A1(n163), .A2(net20298), .B1(n162), .B2(n213), .ZN(n211) );
  AOI22_X1 U370 ( .A1(n229), .A2(net36181), .B1(n235), .B2(net26433), .ZN(n527) );
  AOI22_X1 U371 ( .A1(n95), .A2(net36207), .B1(n164), .B2(net26435), .ZN(n488)
         );
  OAI221_X1 U372 ( .B1(net18459), .B2(net26463), .C1(net26445), .C2(n784), .A(
        n545), .ZN(n151) );
  AOI22_X1 U373 ( .A1(n164), .A2(net36181), .B1(n95), .B2(net26435), .ZN(n545)
         );
  OAI221_X1 U374 ( .B1(net32589), .B2(n783), .C1(net26445), .C2(net18461), .A(
        n522), .ZN(n175) );
  AOI22_X1 U375 ( .A1(n238), .A2(net36207), .B1(n110), .B2(net26437), .ZN(n522) );
  OAI221_X1 U376 ( .B1(net32589), .B2(n761), .C1(net26445), .C2(n783), .A(n509), .ZN(n162) );
  AOI22_X1 U377 ( .A1(n153), .A2(net36207), .B1(n238), .B2(n135), .ZN(n509) );
  OAI221_X1 U378 ( .B1(net32589), .B2(net18461), .C1(net18459), .C2(net26445), 
        .A(n413), .ZN(n136) );
  AOI22_X1 U379 ( .A1(n110), .A2(net36181), .B1(n164), .B2(n135), .ZN(n413) );
  AOI221_X1 U380 ( .B1(n213), .B2(n151), .C1(net20298), .C2(n196), .A(n540), 
        .ZN(n539) );
  OAI22_X1 U381 ( .A1(n779), .A2(net18434), .B1(n541), .B2(net26479), .ZN(n540) );
  INV_X1 U382 ( .A(n150), .ZN(n779) );
  OAI221_X1 U383 ( .B1(net26463), .B2(n787), .C1(net26445), .C2(n262), .A(n544), .ZN(n196) );
  OAI221_X1 U384 ( .B1(net18459), .B2(net32007), .C1(n133), .C2(n784), .A(n270), .ZN(n176) );
  AOI22_X1 U385 ( .A1(n235), .A2(net26473), .B1(n229), .B2(net26449), .ZN(n214) );
  AOI22_X1 U386 ( .A1(n235), .A2(net36181), .B1(n229), .B2(net26437), .ZN(n414) );
  OAI221_X1 U387 ( .B1(n209), .B2(n780), .C1(n208), .C2(n206), .A(net35873), 
        .ZN(n197) );
  NAND2_X1 U388 ( .A1(n232), .A2(A[31]), .ZN(n378) );
  NAND2_X1 U389 ( .A1(n233), .A2(A[31]), .ZN(n339) );
  OAI221_X1 U390 ( .B1(n164), .B2(net26385), .C1(net26415), .C2(n783), .A(
        net26403), .ZN(n504) );
  OAI221_X1 U391 ( .B1(n229), .B2(net26385), .C1(net26415), .C2(n785), .A(
        net26403), .ZN(n159) );
  OAI22_X1 U392 ( .A1(net26445), .A2(net19993), .B1(net26463), .B2(net19990), 
        .ZN(n285) );
  OAI22_X1 U393 ( .A1(net26445), .A2(net19990), .B1(net26463), .B2(n760), .ZN(
        n302) );
  OAI221_X1 U394 ( .B1(n235), .B2(net26385), .C1(net26415), .C2(n784), .A(
        net26403), .ZN(n148) );
  OAI221_X1 U395 ( .B1(n95), .B2(net26385), .C1(net26415), .C2(net18461), .A(
        net26403), .ZN(n519) );
  OAI221_X1 U396 ( .B1(n241), .B2(net26385), .C1(net26415), .C2(n787), .A(
        net26403), .ZN(n184) );
  OAI221_X1 U397 ( .B1(net35313), .B2(net26385), .C1(net18459), .C2(net26415), 
        .A(net26403), .ZN(n127) );
  AOI22_X1 U398 ( .A1(n110), .A2(net36181), .B1(n238), .B2(net26435), .ZN(n465) );
  AOI22_X1 U399 ( .A1(n164), .A2(net36181), .B1(n110), .B2(net26437), .ZN(n474) );
  AOI22_X1 U400 ( .A1(net35295), .A2(net36181), .B1(n173), .B2(net26437), .ZN(
        n543) );
  AOI211_X1 U401 ( .C1(A[27]), .C2(net36207), .A(n253), .B(n254), .ZN(n247) );
  OAI22_X1 U402 ( .A1(n776), .A2(net18434), .B1(n217), .B2(net26479), .ZN(n209) );
  OAI22_X1 U403 ( .A1(net26445), .A2(n788), .B1(net32589), .B2(n262), .ZN(n220) );
  OAI22_X1 U404 ( .A1(n777), .A2(net18434), .B1(n271), .B2(net26479), .ZN(n268) );
  OAI22_X1 U405 ( .A1(net26445), .A2(n789), .B1(net32589), .B2(n788), .ZN(n272) );
  OAI22_X1 U406 ( .A1(n778), .A2(net18434), .B1(n415), .B2(net26479), .ZN(n410) );
  AOI221_X1 U407 ( .B1(n177), .B2(net36207), .C1(n243), .C2(net26435), .A(n416), .ZN(n415) );
  OAI22_X1 U408 ( .A1(net26445), .A2(n790), .B1(net32589), .B2(n789), .ZN(n416) );
  AOI22_X1 U409 ( .A1(n24), .A2(net26423), .B1(n230), .B2(net26431), .ZN(n521)
         );
  AOI22_X1 U410 ( .A1(n167), .A2(net26423), .B1(n24), .B2(net26433), .ZN(n508)
         );
  AOI22_X1 U411 ( .A1(n230), .A2(net26423), .B1(A[19]), .B2(net26431), .ZN(
        n483) );
  AOI22_X1 U412 ( .A1(A[19]), .A2(net36181), .B1(A[18]), .B2(net26435), .ZN(
        n549) );
  INV_X1 U413 ( .A(n164), .ZN(n783) );
  AOI22_X1 U414 ( .A1(A[23]), .A2(net36181), .B1(n167), .B2(net26433), .ZN(
        n550) );
  AOI22_X1 U415 ( .A1(n34), .A2(net36181), .B1(net35295), .B2(n135), .ZN(n485)
         );
  AOI22_X1 U416 ( .A1(n169), .A2(net26423), .B1(A[23]), .B2(net26431), .ZN(
        n484) );
  AOI22_X1 U417 ( .A1(n238), .A2(net36181), .B1(n153), .B2(net26435), .ZN(n454) );
  OAI21_X1 U418 ( .B1(n233), .B2(net26383), .A(net26403), .ZN(n203) );
  OAI21_X1 U419 ( .B1(n231), .B2(net26383), .A(net26403), .ZN(n183) );
  OAI21_X1 U420 ( .B1(n227), .B2(net26383), .A(net26403), .ZN(n170) );
  OAI21_X1 U421 ( .B1(n190), .B2(net26383), .A(net26403), .ZN(n157) );
  OAI21_X1 U422 ( .B1(n237), .B2(net26383), .A(net26403), .ZN(n146) );
  OAI21_X1 U423 ( .B1(n160), .B2(net26383), .A(net26407), .ZN(n192) );
  OAI21_X1 U424 ( .B1(n180), .B2(net26383), .A(net26407), .ZN(n121) );
  OAI21_X1 U425 ( .B1(n103), .B2(net26383), .A(net26407), .ZN(n518) );
  OAI21_X1 U426 ( .B1(n201), .B2(net26383), .A(net26403), .ZN(n503) );
  AOI22_X1 U427 ( .A1(A[28]), .A2(net26425), .B1(A[27]), .B2(net26431), .ZN(
        n482) );
  AOI22_X1 U428 ( .A1(A[27]), .A2(net36181), .B1(n154), .B2(net26435), .ZN(
        n547) );
  AOI22_X1 U429 ( .A1(n137), .A2(net36207), .B1(n34), .B2(n135), .ZN(n523) );
  AOI22_X1 U430 ( .A1(n33), .A2(net26423), .B1(n169), .B2(net26431), .ZN(n520)
         );
  AOI22_X1 U431 ( .A1(n154), .A2(net26425), .B1(n33), .B2(net26437), .ZN(n506)
         );
  AOI22_X1 U432 ( .A1(A[18]), .A2(net36207), .B1(n137), .B2(n135), .ZN(n507)
         );
  AND2_X1 U433 ( .A1(n758), .A2(n759), .ZN(net31776) );
  AND2_X1 U434 ( .A1(n278), .A2(n277), .ZN(net31396) );
  AND2_X1 U435 ( .A1(FUNC[2]), .A2(n759), .ZN(net31364) );
  AND2_X1 U436 ( .A1(FUNC[0]), .A2(n758), .ZN(net31363) );
  AND2_X1 U437 ( .A1(FUNC[2]), .A2(FUNC[0]), .ZN(net31362) );
  AND2_X1 U438 ( .A1(FUNC[1]), .A2(n278), .ZN(net31345) );
  OAI221_X1 U439 ( .B1(n244), .B2(net26385), .C1(net26415), .C2(n786), .A(
        net26403), .ZN(n172) );
  AOI22_X1 U440 ( .A1(n241), .A2(net36207), .B1(n244), .B2(n135), .ZN(n497) );
  AOI22_X1 U441 ( .A1(n244), .A2(net36181), .B1(n229), .B2(n135), .ZN(n489) );
  AOI22_X1 U442 ( .A1(n229), .A2(net36181), .B1(n244), .B2(n135), .ZN(n544) );
  AOI22_X1 U443 ( .A1(n229), .A2(net26469), .B1(n244), .B2(net26449), .ZN(n270) );
  INV_X1 U444 ( .A(n177), .ZN(n262) );
  AOI221_X1 U445 ( .B1(n243), .B2(net31778), .C1(net26397), .C2(n788), .A(
        net31788), .ZN(n202) );
  AOI22_X1 U446 ( .A1(net20016), .A2(n773), .B1(n243), .B2(n203), .ZN(n198) );
  AOI211_X1 U447 ( .C1(n243), .C2(net36207), .A(n542), .B(n757), .ZN(n541) );
  AOI22_X1 U448 ( .A1(n536), .A2(n537), .B1(n273), .B2(n538), .ZN(n530) );
  AOI22_X1 U449 ( .A1(net26397), .A2(n764), .B1(net31778), .B2(n273), .ZN(n534) );
  OAI21_X1 U450 ( .B1(n83), .B2(net26383), .A(net26407), .ZN(n406) );
  INV_X1 U451 ( .A(n240), .ZN(n791) );
  OAI21_X1 U452 ( .B1(n165), .B2(net26383), .A(net26403), .ZN(n538) );
  AOI22_X1 U453 ( .A1(n165), .A2(net36207), .B1(n260), .B2(n135), .ZN(n512) );
  AOI22_X1 U454 ( .A1(N794), .A2(n759), .B1(N795), .B2(FUNC[0]), .ZN(n552) );
  OAI21_X1 U455 ( .B1(n552), .B2(FUNC[1]), .A(n553), .ZN(n551) );
  AOI22_X1 U456 ( .A1(net20016), .A2(n774), .B1(n261), .B2(n264), .ZN(n259) );
  AOI22_X1 U457 ( .A1(n261), .A2(net36181), .B1(n243), .B2(n135), .ZN(n487) );
  AOI22_X1 U459 ( .A1(n260), .A2(net36181), .B1(n149), .B2(n135), .ZN(n496) );
  OAI221_X1 U460 ( .B1(n177), .B2(net26385), .C1(net26415), .C2(n262), .A(
        net26403), .ZN(n195) );
  AOI22_X1 U461 ( .A1(n243), .A2(net36207), .B1(n177), .B2(net26433), .ZN(n528) );
  AOI22_X1 U462 ( .A1(n177), .A2(net36181), .B1(n241), .B2(n135), .ZN(n513) );
  INV_X1 U463 ( .A(net26479), .ZN(net26483) );
  INV_X1 U464 ( .A(net26479), .ZN(net26485) );
  INV_X1 U465 ( .A(n40), .ZN(net26465) );
  INV_X1 U466 ( .A(net31778), .ZN(net26415) );
  INV_X1 U467 ( .A(net31788), .ZN(net26403) );
  INV_X1 U468 ( .A(n123), .ZN(net26397) );
  INV_X1 U469 ( .A(n240), .ZN(n276) );
  INV_X1 U470 ( .A(B[0]), .ZN(n764) );
  NAND2_X1 U471 ( .A1(n276), .A2(n764), .ZN(net18425) );
  NAND2_X1 U472 ( .A1(n238), .A2(net26469), .ZN(n428) );
  NAND2_X1 U473 ( .A1(net26455), .A2(n110), .ZN(n372) );
  NAND3_X1 U474 ( .A1(n543), .A2(n428), .A3(n372), .ZN(n150) );
  INV_X1 U475 ( .A(FUNC[2]), .ZN(n758) );
  INV_X1 U476 ( .A(FUNC[3]), .ZN(n278) );
  INV_X1 U477 ( .A(B[2]), .ZN(n763) );
  INV_X1 U478 ( .A(FUNC[1]), .ZN(n277) );
  NAND2_X1 U479 ( .A1(n78), .A2(n5), .ZN(n296) );
  NAND2_X1 U480 ( .A1(n165), .A2(net26455), .ZN(n626) );
  INV_X1 U481 ( .A(FUNC[0]), .ZN(n759) );
  INV_X1 U482 ( .A(n165), .ZN(n287) );
  AOI21_X1 U483 ( .B1(n534), .B2(net26403), .A(n287), .ZN(n280) );
  AOI221_X1 U484 ( .B1(N59), .B2(net26493), .C1(N91), .C2(net26497), .A(n280), 
        .ZN(n281) );
  NAND3_X1 U485 ( .A1(A[31]), .A2(N19), .A3(net24726), .ZN(n358) );
  AND3_X1 U486 ( .A1(n281), .A2(n358), .A3(n530), .ZN(n282) );
  OAI211_X1 U487 ( .C1(n466), .C2(n626), .A(n529), .B(n282), .ZN(RES[0]) );
  AOI22_X1 U488 ( .A1(N92), .A2(net26499), .B1(N60), .B2(net26495), .ZN(n286)
         );
  OAI22_X1 U489 ( .A1(net26445), .A2(n790), .B1(net32589), .B2(n287), .ZN(n712) );
  NAND2_X1 U490 ( .A1(n401), .A2(n402), .ZN(n283) );
  INV_X1 U491 ( .A(n358), .ZN(n341) );
  AOI211_X1 U492 ( .C1(n248), .C2(n712), .A(n283), .B(n341), .ZN(n284) );
  OAI211_X1 U493 ( .C1(n405), .C2(n791), .A(n286), .B(n284), .ZN(RES[1]) );
  AOI22_X1 U494 ( .A1(N93), .A2(net26497), .B1(N61), .B2(net26495), .ZN(n290)
         );
  INV_X1 U495 ( .A(n261), .ZN(n789) );
  OAI222_X1 U496 ( .A1(n789), .A2(n134), .B1(n16), .B2(n287), .C1(net26465), 
        .C2(n790), .ZN(n733) );
  NAND2_X1 U497 ( .A1(n259), .A2(n258), .ZN(n288) );
  AOI211_X1 U498 ( .C1(n182), .C2(n733), .A(n288), .B(n341), .ZN(n289) );
  OAI211_X1 U499 ( .C1(n263), .C2(n181), .A(n290), .B(n289), .ZN(RES[2]) );
  AOI22_X1 U500 ( .A1(N94), .A2(net26499), .B1(N62), .B2(net26493), .ZN(n293)
         );
  INV_X1 U501 ( .A(n243), .ZN(n788) );
  OAI221_X1 U502 ( .B1(n789), .B2(net26461), .C1(n788), .C2(n134), .A(n512), 
        .ZN(net24464) );
  NAND2_X1 U503 ( .A1(n197), .A2(n198), .ZN(n291) );
  AOI211_X1 U504 ( .C1(n246), .C2(net24464), .A(n291), .B(n341), .ZN(n292) );
  OAI211_X1 U505 ( .C1(n202), .C2(n30), .A(n293), .B(n292), .ZN(RES[3]) );
  INV_X1 U506 ( .A(A[28]), .ZN(net19990) );
  AOI22_X1 U507 ( .A1(A[30]), .A2(n135), .B1(A[31]), .B2(net26425), .ZN(n294)
         );
  OAI221_X1 U508 ( .B1(net19993), .B2(net32589), .C1(net19990), .C2(n134), .A(
        n294), .ZN(n379) );
  INV_X1 U509 ( .A(n379), .ZN(n462) );
  NAND2_X1 U510 ( .A1(n24), .A2(net26473), .ZN(n599) );
  NAND2_X1 U511 ( .A1(n230), .A2(net26453), .ZN(n567) );
  NAND3_X1 U512 ( .A1(n550), .A2(n599), .A3(n567), .ZN(n459) );
  INV_X1 U513 ( .A(n459), .ZN(n331) );
  NAND2_X1 U514 ( .A1(n33), .A2(net26473), .ZN(n664) );
  NAND2_X1 U515 ( .A1(n169), .A2(net26453), .ZN(n631) );
  NAND3_X1 U516 ( .A1(n547), .A2(n664), .A3(n631), .ZN(n369) );
  INV_X1 U517 ( .A(n369), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n274), .A2(n762), .ZN(net26700) );
  OAI222_X1 U519 ( .A1(n462), .A2(net24561), .B1(net26479), .B2(n331), .C1(
        n461), .C2(net26700), .ZN(n572) );
  NOR2_X1 U520 ( .A1(n233), .A2(n296), .ZN(n297) );
  OAI221_X1 U521 ( .B1(n788), .B2(net32589), .C1(n262), .C2(n134), .A(n496), 
        .ZN(n453) );
  INV_X1 U522 ( .A(n453), .ZN(n627) );
  MUX2_X1 U523 ( .A(n627), .B(n626), .S(n274), .Z(n695) );
  INV_X1 U524 ( .A(n695), .ZN(n563) );
  AOI221_X1 U525 ( .B1(n131), .B2(n572), .C1(n297), .C2(n563), .A(n341), .ZN(
        n304) );
  INV_X1 U526 ( .A(n524), .ZN(net24911) );
  NAND2_X1 U527 ( .A1(n78), .A2(net24911), .ZN(n464) );
  INV_X1 U528 ( .A(n464), .ZN(n299) );
  INV_X1 U529 ( .A(n572), .ZN(n298) );
  NAND2_X1 U530 ( .A1(n298), .A2(n378), .ZN(n574) );
  NAND2_X1 U531 ( .A1(n137), .A2(net26469), .ZN(n502) );
  NAND2_X1 U532 ( .A1(n34), .A2(net26453), .ZN(n456) );
  NAND3_X1 U533 ( .A1(n549), .A2(n502), .A3(n456), .ZN(n458) );
  AOI222_X1 U534 ( .A1(n151), .A2(n444), .B1(n84), .B2(n574), .C1(n185), .C2(
        n458), .ZN(n303) );
  AOI222_X1 U535 ( .A1(N95), .A2(net26497), .B1(n252), .B2(n150), .C1(n196), 
        .C2(n224), .ZN(n301) );
  AOI222_X1 U536 ( .A1(n192), .A2(n177), .B1(N63), .B2(net26495), .C1(n160), 
        .C2(n195), .ZN(n300) );
  NAND4_X1 U537 ( .A1(n301), .A2(n303), .A3(n304), .A4(n300), .ZN(RES[4]) );
  NAND2_X1 U538 ( .A1(n167), .A2(net26467), .ZN(n615) );
  NAND2_X1 U539 ( .A1(n24), .A2(net26453), .ZN(n583) );
  NAND2_X1 U540 ( .A1(n154), .A2(n39), .ZN(n680) );
  NAND2_X1 U541 ( .A1(n33), .A2(net26453), .ZN(n647) );
  NAND3_X1 U542 ( .A1(n482), .A2(n680), .A3(n647), .ZN(n337) );
  INV_X1 U543 ( .A(n337), .ZN(n473) );
  OAI22_X1 U544 ( .A1(net26479), .A2(n48), .B1(n473), .B2(net26700), .ZN(n305)
         );
  INV_X1 U545 ( .A(n305), .ZN(n307) );
  OAI211_X1 U546 ( .C1(n338), .C2(net24561), .A(n307), .B(n378), .ZN(n588) );
  NAND2_X1 U547 ( .A1(A[18]), .A2(net26467), .ZN(n548) );
  NAND2_X1 U548 ( .A1(n137), .A2(net26453), .ZN(n491) );
  INV_X1 U549 ( .A(n712), .ZN(n342) );
  OAI21_X1 U550 ( .B1(n342), .B2(n249), .A(n358), .ZN(n306) );
  AOI221_X1 U551 ( .B1(n84), .B2(n588), .C1(n185), .C2(n472), .A(n306), .ZN(
        n311) );
  INV_X1 U552 ( .A(n241), .ZN(n787) );
  OAI221_X1 U553 ( .B1(n262), .B2(net32589), .C1(n787), .C2(n134), .A(n487), 
        .ZN(n713) );
  NAND2_X1 U554 ( .A1(n153), .A2(net26469), .ZN(n440) );
  NAND2_X1 U555 ( .A1(n238), .A2(net26453), .ZN(n396) );
  NAND3_X1 U556 ( .A1(n485), .A2(n440), .A3(n396), .ZN(n397) );
  INV_X1 U557 ( .A(A[31]), .ZN(net24891) );
  INV_X1 U558 ( .A(n480), .ZN(net24901) );
  INV_X1 U559 ( .A(n390), .ZN(n728) );
  OAI21_X1 U560 ( .B1(n728), .B2(net24561), .A(n307), .ZN(n589) );
  AOI222_X1 U561 ( .A1(n246), .A2(n713), .B1(n252), .B2(n397), .C1(n131), .C2(
        n589), .ZN(n310) );
  AOI222_X1 U562 ( .A1(n183), .A2(n241), .B1(N64), .B2(net26495), .C1(n231), 
        .C2(n184), .ZN(n308) );
  NAND4_X1 U563 ( .A1(n311), .A2(n310), .A3(n309), .A4(n308), .ZN(RES[5]) );
  NAND2_X1 U564 ( .A1(net26455), .A2(A[30]), .ZN(n756) );
  OAI21_X1 U565 ( .B1(net26455), .B2(net24891), .A(n756), .ZN(n312) );
  INV_X1 U566 ( .A(n312), .ZN(n746) );
  NAND2_X1 U567 ( .A1(A[23]), .A2(n39), .ZN(n632) );
  NAND2_X1 U568 ( .A1(n167), .A2(net26451), .ZN(n600) );
  NAND3_X1 U569 ( .A1(n520), .A2(n632), .A3(n600), .ZN(n430) );
  INV_X1 U570 ( .A(A[27]), .ZN(n760) );
  NAND2_X1 U571 ( .A1(n154), .A2(net26451), .ZN(n665) );
  AOI22_X1 U572 ( .A1(A[28]), .A2(net26431), .B1(A[29]), .B2(net26425), .ZN(
        n313) );
  OAI211_X1 U573 ( .C1(n760), .C2(net32589), .A(n665), .B(n313), .ZN(n347) );
  INV_X1 U574 ( .A(n347), .ZN(n499) );
  OAI22_X1 U575 ( .A1(net26479), .A2(n20), .B1(n499), .B2(net26700), .ZN(n314)
         );
  INV_X1 U576 ( .A(n314), .ZN(n316) );
  OAI211_X1 U577 ( .C1(n746), .C2(net24561), .A(n378), .B(n316), .ZN(n605) );
  NAND2_X1 U578 ( .A1(A[19]), .A2(n40), .ZN(n568) );
  NAND2_X1 U579 ( .A1(A[18]), .A2(net26451), .ZN(n505) );
  INV_X1 U580 ( .A(n733), .ZN(n658) );
  OAI21_X1 U581 ( .B1(n658), .B2(n249), .A(n358), .ZN(n315) );
  AOI221_X1 U582 ( .B1(n84), .B2(n605), .C1(n185), .C2(n498), .A(n315), .ZN(
        n320) );
  INV_X1 U583 ( .A(n244), .ZN(n786) );
  OAI221_X1 U584 ( .B1(n787), .B2(net26465), .C1(n786), .C2(n134), .A(n528), 
        .ZN(n734) );
  NAND2_X1 U585 ( .A1(net35295), .A2(net26473), .ZN(n457) );
  NAND2_X1 U586 ( .A1(n153), .A2(net26451), .ZN(n427) );
  NAND3_X1 U587 ( .A1(n523), .A2(n457), .A3(n427), .ZN(n351) );
  OAI21_X1 U588 ( .B1(net26461), .B2(net24891), .A(n756), .ZN(n421) );
  INV_X1 U589 ( .A(n421), .ZN(n752) );
  OAI21_X1 U590 ( .B1(n752), .B2(net24561), .A(n316), .ZN(n604) );
  AOI222_X1 U591 ( .A1(n248), .A2(n734), .B1(n252), .B2(n351), .C1(n131), .C2(
        n604), .ZN(n319) );
  AOI222_X1 U592 ( .A1(N97), .A2(net26497), .B1(n175), .B2(n444), .C1(n176), 
        .C2(n370), .ZN(n318) );
  AOI222_X1 U593 ( .A1(n170), .A2(n244), .B1(N65), .B2(net26495), .C1(n227), 
        .C2(n172), .ZN(n317) );
  NAND4_X1 U594 ( .A1(n320), .A2(n319), .A3(n318), .A4(n317), .ZN(RES[6]) );
  NAND2_X1 U595 ( .A1(n169), .A2(n40), .ZN(n648) );
  NAND2_X1 U596 ( .A1(A[23]), .A2(net26451), .ZN(n616) );
  NAND3_X1 U597 ( .A1(n506), .A2(n648), .A3(n616), .ZN(n445) );
  INV_X1 U598 ( .A(n445), .ZN(n531) );
  NAND2_X1 U599 ( .A1(net26455), .A2(A[27]), .ZN(n681) );
  AOI22_X1 U600 ( .A1(A[29]), .A2(net26435), .B1(A[30]), .B2(net26423), .ZN(
        n321) );
  OAI211_X1 U601 ( .C1(net19990), .C2(net26461), .A(n681), .B(n321), .ZN(n357)
         );
  INV_X1 U602 ( .A(n357), .ZN(n532) );
  OAI22_X1 U603 ( .A1(net26479), .A2(n531), .B1(n532), .B2(net26700), .ZN(n322) );
  INV_X1 U604 ( .A(n322), .ZN(n324) );
  NAND2_X1 U605 ( .A1(n324), .A2(n339), .ZN(n621) );
  NAND2_X1 U606 ( .A1(n230), .A2(n40), .ZN(n584) );
  NAND2_X1 U607 ( .A1(A[19]), .A2(net26451), .ZN(n554) );
  NAND3_X1 U608 ( .A1(n508), .A2(n584), .A3(n554), .ZN(n526) );
  INV_X1 U609 ( .A(net24464), .ZN(net24560) );
  OAI21_X1 U610 ( .B1(net24560), .B2(n249), .A(n358), .ZN(n323) );
  AOI221_X1 U611 ( .B1(n84), .B2(n621), .C1(n188), .C2(n526), .A(n323), .ZN(
        n328) );
  INV_X1 U612 ( .A(n229), .ZN(n785) );
  OAI221_X1 U613 ( .B1(n786), .B2(net32589), .C1(n785), .C2(n134), .A(n513), 
        .ZN(net24463) );
  NAND2_X1 U614 ( .A1(n34), .A2(net26473), .ZN(n490) );
  NAND2_X1 U615 ( .A1(net35295), .A2(net26451), .ZN(n439) );
  NAND3_X1 U616 ( .A1(n507), .A2(n490), .A3(n439), .ZN(n362) );
  NAND2_X1 U617 ( .A1(A[31]), .A2(net26449), .ZN(net24439) );
  OAI21_X1 U618 ( .B1(net24439), .B2(net24561), .A(n324), .ZN(n620) );
  AOI222_X1 U619 ( .A1(n182), .A2(net24463), .B1(n252), .B2(n362), .C1(n131), 
        .C2(n620), .ZN(n327) );
  AOI222_X1 U620 ( .A1(N98), .A2(net26497), .B1(n162), .B2(n444), .C1(n163), 
        .C2(n370), .ZN(n326) );
  AOI222_X1 U621 ( .A1(n157), .A2(n229), .B1(N66), .B2(net26495), .C1(n190), 
        .C2(n159), .ZN(n325) );
  NAND4_X1 U622 ( .A1(n328), .A2(n327), .A3(n326), .A4(n325), .ZN(RES[7]) );
  INV_X1 U623 ( .A(n626), .ZN(n757) );
  NAND2_X1 U624 ( .A1(n22), .A2(n213), .ZN(n424) );
  OAI22_X1 U625 ( .A1(net26479), .A2(n461), .B1(n462), .B2(net26700), .ZN(n636) );
  INV_X1 U626 ( .A(n636), .ZN(n330) );
  INV_X1 U627 ( .A(n131), .ZN(n380) );
  OAI21_X1 U628 ( .B1(n330), .B2(n380), .A(n358), .ZN(n329) );
  AOI221_X1 U629 ( .B1(n757), .B2(n29), .C1(n687), .C2(n453), .A(n329), .ZN(
        n336) );
  NAND2_X1 U630 ( .A1(n330), .A2(n339), .ZN(n637) );
  INV_X1 U631 ( .A(n235), .ZN(n784) );
  OAI221_X1 U632 ( .B1(n785), .B2(net26463), .C1(n784), .C2(n134), .A(n497), 
        .ZN(n573) );
  AOI222_X1 U633 ( .A1(n252), .A2(n458), .B1(n84), .B2(n637), .C1(n686), .C2(
        n573), .ZN(n335) );
  OAI22_X1 U634 ( .A1(n779), .A2(n363), .B1(n331), .B2(n442), .ZN(n332) );
  AOI221_X1 U635 ( .B1(n151), .B2(n224), .C1(N99), .C2(net26497), .A(n332), 
        .ZN(n334) );
  AOI222_X1 U636 ( .A1(n146), .A2(n235), .B1(N67), .B2(net26495), .C1(n237), 
        .C2(n148), .ZN(n333) );
  NAND4_X1 U637 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .ZN(RES[8]) );
  NAND2_X1 U638 ( .A1(n337), .A2(net26483), .ZN(n340) );
  OAI211_X1 U639 ( .C1(n338), .C2(net26700), .A(n339), .B(n340), .ZN(n652) );
  OAI21_X1 U640 ( .B1(n728), .B2(net26700), .A(n340), .ZN(n645) );
  INV_X1 U641 ( .A(n713), .ZN(n393) );
  INV_X1 U642 ( .A(net35313), .ZN(net18459) );
  OAI221_X1 U643 ( .B1(n784), .B2(net26463), .C1(net18459), .C2(n134), .A(n489), .ZN(n590) );
  INV_X1 U644 ( .A(n590), .ZN(n715) );
  AOI222_X1 U645 ( .A1(N100), .A2(net26497), .B1(n185), .B2(n399), .C1(n136), 
        .C2(n370), .ZN(n344) );
  AOI222_X1 U646 ( .A1(n121), .A2(net35313), .B1(N68), .B2(net26495), .C1(n180), .C2(n127), .ZN(n343) );
  NAND4_X1 U647 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(RES[9]) );
  NAND2_X1 U648 ( .A1(n45), .A2(net26485), .ZN(n350) );
  OAI21_X1 U649 ( .B1(n752), .B2(net26700), .A(n350), .ZN(n669) );
  INV_X1 U650 ( .A(n669), .ZN(n348) );
  OAI21_X1 U651 ( .B1(n348), .B2(n380), .A(n358), .ZN(n349) );
  AOI221_X1 U652 ( .B1(n212), .B2(n733), .C1(n687), .C2(n734), .A(n349), .ZN(
        n356) );
  OAI211_X1 U653 ( .C1(n746), .C2(net26700), .A(n339), .B(n350), .ZN(n670) );
  INV_X1 U654 ( .A(net34396), .ZN(net18461) );
  OAI221_X1 U655 ( .B1(net18459), .B2(net32589), .C1(net18461), .C2(n134), .A(
        n527), .ZN(n606) );
  AOI222_X1 U656 ( .A1(n498), .A2(n252), .B1(n84), .B2(n670), .C1(n686), .C2(
        n606), .ZN(n355) );
  INV_X1 U657 ( .A(n351), .ZN(n777) );
  OAI22_X1 U658 ( .A1(n20), .A2(n442), .B1(n777), .B2(n363), .ZN(n352) );
  AOI221_X1 U659 ( .B1(n175), .B2(n224), .C1(N101), .C2(net26497), .A(n352), 
        .ZN(n354) );
  AOI222_X1 U660 ( .A1(n518), .A2(n95), .B1(N69), .B2(net26495), .C1(n103), 
        .C2(n519), .ZN(n353) );
  NAND4_X1 U661 ( .A1(n356), .A2(n355), .A3(n354), .A4(n353), .ZN(RES[10]) );
  NAND2_X1 U662 ( .A1(n357), .A2(net26483), .ZN(n682) );
  NAND3_X1 U663 ( .A1(n84), .A2(A[31]), .A3(net26479), .ZN(n359) );
  NAND2_X1 U664 ( .A1(n359), .A2(n358), .ZN(n382) );
  INV_X1 U665 ( .A(n382), .ZN(n418) );
  OAI21_X1 U666 ( .B1(n682), .B2(n381), .A(n418), .ZN(n360) );
  OAI21_X1 U667 ( .B1(net24439), .B2(net26700), .A(n682), .ZN(n688) );
  AOI22_X1 U668 ( .A1(net36181), .A2(n235), .B1(net26435), .B2(net35313), .ZN(
        n361) );
  OAI221_X1 U669 ( .B1(net18461), .B2(net26461), .C1(n134), .C2(n783), .A(n361), .ZN(net24562) );
  AOI222_X1 U670 ( .A1(n252), .A2(n526), .B1(n131), .B2(n688), .C1(n686), .C2(
        net24562), .ZN(n367) );
  INV_X1 U671 ( .A(n362), .ZN(n776) );
  OAI22_X1 U672 ( .A1(n531), .A2(n442), .B1(n776), .B2(n363), .ZN(n364) );
  AOI221_X1 U673 ( .B1(n162), .B2(n224), .C1(N102), .C2(net26497), .A(n364), 
        .ZN(n366) );
  AOI222_X1 U674 ( .A1(n503), .A2(n164), .B1(N70), .B2(net26495), .C1(n201), 
        .C2(n504), .ZN(n365) );
  NAND4_X1 U675 ( .A1(n368), .A2(n367), .A3(n366), .A4(n365), .ZN(RES[11]) );
  AOI222_X1 U676 ( .A1(n252), .A2(n459), .B1(n444), .B2(n458), .C1(n185), .C2(
        n369), .ZN(n388) );
  AOI222_X1 U677 ( .A1(N71), .A2(net26493), .B1(n224), .B2(n150), .C1(N103), 
        .C2(net26499), .ZN(n387) );
  INV_X1 U678 ( .A(n573), .ZN(n697) );
  AOI22_X1 U679 ( .A1(net36207), .A2(net35313), .B1(n95), .B2(net26433), .ZN(
        n371) );
  OAI211_X1 U680 ( .C1(net26463), .C2(n783), .A(n372), .B(n371), .ZN(n638) );
  INV_X1 U681 ( .A(n638), .ZN(n696) );
  MUX2_X1 U682 ( .A(net26397), .B(net31778), .S(n200), .Z(n373) );
  OAI21_X1 U683 ( .B1(net31788), .B2(n373), .A(n110), .ZN(n374) );
  OAI221_X1 U684 ( .B1(n697), .B2(n249), .C1(n696), .C2(n466), .A(n374), .ZN(
        n385) );
  INV_X1 U685 ( .A(n110), .ZN(n761) );
  AOI21_X1 U686 ( .B1(net26397), .B2(n761), .A(net31788), .ZN(n377) );
  INV_X1 U687 ( .A(n200), .ZN(n376) );
  NAND3_X1 U688 ( .A1(n22), .A2(n233), .A3(n563), .ZN(n375) );
  OAI21_X1 U689 ( .B1(n377), .B2(n376), .A(n375), .ZN(n384) );
  NAND2_X1 U690 ( .A1(n379), .A2(net26485), .ZN(n693) );
  AOI21_X1 U691 ( .B1(n381), .B2(n380), .A(n693), .ZN(n383) );
  NOR4_X1 U692 ( .A1(n385), .A2(n384), .A3(n383), .A4(n382), .ZN(n386) );
  NAND3_X1 U693 ( .A1(n388), .A2(n387), .A3(n386), .ZN(RES[12]) );
  OAI21_X1 U694 ( .B1(n238), .B2(net26385), .A(net26407), .ZN(n391) );
  NAND2_X1 U695 ( .A1(n84), .A2(net26483), .ZN(n419) );
  OAI21_X1 U696 ( .B1(n338), .B2(n419), .A(n418), .ZN(n389) );
  AOI221_X1 U697 ( .B1(n158), .B2(n391), .C1(net32250), .C2(n390), .A(n389), 
        .ZN(n417) );
  MUX2_X1 U698 ( .A(net26387), .B(net26415), .S(n158), .Z(n392) );
  NAND2_X1 U699 ( .A1(n392), .A2(net26407), .ZN(n395) );
  OAI22_X1 U700 ( .A1(n715), .A2(n249), .B1(n393), .B2(n424), .ZN(n394) );
  OAI211_X1 U701 ( .C1(n761), .C2(net26463), .A(n488), .B(n396), .ZN(n711) );
  INV_X1 U702 ( .A(n397), .ZN(n778) );
  OAI22_X1 U703 ( .A1(n473), .A2(n442), .B1(n778), .B2(n441), .ZN(n398) );
  AOI221_X1 U704 ( .B1(n248), .B2(n711), .C1(n199), .C2(n472), .A(n398), .ZN(
        n403) );
  AOI222_X1 U705 ( .A1(N72), .A2(net26493), .B1(n252), .B2(n399), .C1(N104), 
        .C2(net26501), .ZN(n400) );
  NAND4_X1 U706 ( .A1(n403), .A2(n404), .A3(n417), .A4(n400), .ZN(RES[13]) );
  OAI21_X1 U707 ( .B1(n153), .B2(net26385), .A(net26403), .ZN(n422) );
  OAI21_X1 U708 ( .B1(n746), .B2(n419), .A(n418), .ZN(n420) );
  AOI221_X1 U709 ( .B1(n156), .B2(n422), .C1(net32250), .C2(n421), .A(n420), 
        .ZN(n434) );
  MUX2_X1 U710 ( .A(net26385), .B(net26415), .S(n156), .Z(n423) );
  NAND2_X1 U711 ( .A1(n423), .A2(net26407), .ZN(n426) );
  INV_X1 U712 ( .A(n606), .ZN(n736) );
  INV_X1 U713 ( .A(n734), .ZN(n659) );
  OAI22_X1 U714 ( .A1(n736), .A2(n249), .B1(n659), .B2(n424), .ZN(n425) );
  AOI221_X1 U715 ( .B1(n153), .B2(n426), .C1(n255), .C2(n733), .A(n425), .ZN(
        n433) );
  NAND3_X1 U716 ( .A1(n474), .A2(n428), .A3(n427), .ZN(n732) );
  OAI22_X1 U717 ( .A1(n499), .A2(n442), .B1(n777), .B2(n441), .ZN(n429) );
  AOI221_X1 U718 ( .B1(n248), .B2(n732), .C1(n199), .C2(n498), .A(n429), .ZN(
        n432) );
  AOI222_X1 U719 ( .A1(N73), .A2(net26493), .B1(n252), .B2(n430), .C1(N105), 
        .C2(net26501), .ZN(n431) );
  NAND4_X1 U720 ( .A1(n434), .A2(n433), .A3(n432), .A4(n431), .ZN(RES[14]) );
  MUX2_X1 U721 ( .A(net26385), .B(net26415), .S(n73), .Z(n435) );
  NAND2_X1 U722 ( .A1(n435), .A2(net26403), .ZN(net24772) );
  INV_X1 U723 ( .A(net35295), .ZN(net24777) );
  AOI21_X1 U724 ( .B1(net26397), .B2(net24777), .A(net31788), .ZN(n438) );
  INV_X1 U725 ( .A(n73), .ZN(n437) );
  NAND3_X1 U726 ( .A1(A[31]), .A2(net24726), .A3(n436), .ZN(n675) );
  OAI21_X1 U727 ( .B1(n438), .B2(n437), .A(n675), .ZN(net24773) );
  NAND3_X1 U728 ( .A1(n465), .A2(n440), .A3(n439), .ZN(net24465) );
  OAI22_X1 U729 ( .A1(n532), .A2(n442), .B1(n776), .B2(n441), .ZN(n443) );
  AOI221_X1 U730 ( .B1(n248), .B2(net24465), .C1(n199), .C2(n526), .A(n443), 
        .ZN(n447) );
  AOI222_X1 U731 ( .A1(N74), .A2(net26493), .B1(n252), .B2(n445), .C1(N106), 
        .C2(net26501), .ZN(n446) );
  NAND4_X1 U732 ( .A1(n446), .A2(n448), .A3(n447), .A4(net24759), .ZN(RES[15])
         );
  NAND2_X1 U733 ( .A1(n5), .A2(net20016), .ZN(n562) );
  INV_X1 U734 ( .A(n562), .ZN(n678) );
  OAI21_X1 U735 ( .B1(n34), .B2(net26385), .A(net26407), .ZN(n449) );
  INV_X1 U736 ( .A(n675), .ZN(n660) );
  AOI221_X1 U737 ( .B1(n251), .B2(n757), .C1(B[16]), .C2(n449), .A(n660), .ZN(
        n471) );
  MUX2_X1 U738 ( .A(net26385), .B(net26415), .S(B[16]), .Z(n451) );
  INV_X1 U739 ( .A(A[16]), .ZN(n450) );
  AOI21_X1 U740 ( .B1(n451), .B2(net26407), .A(n450), .ZN(n452) );
  AOI221_X1 U741 ( .B1(n29), .B2(n573), .C1(n255), .C2(n453), .A(n452), .ZN(
        n470) );
  NAND3_X1 U742 ( .A1(n454), .A2(n457), .A3(n456), .ZN(n639) );
  INV_X1 U743 ( .A(n639), .ZN(n701) );
  INV_X1 U744 ( .A(n232), .ZN(net18434) );
  AOI22_X1 U745 ( .A1(net20298), .A2(n459), .B1(n458), .B2(net26483), .ZN(n460) );
  OAI221_X1 U746 ( .B1(net18434), .B2(n462), .C1(n461), .C2(net24561), .A(n460), .ZN(n463) );
  INV_X1 U747 ( .A(n463), .ZN(n455) );
  OAI222_X1 U748 ( .A1(n696), .A2(n249), .B1(n701), .B2(n466), .C1(n455), .C2(
        n464), .ZN(n468) );
  AOI221_X1 U749 ( .B1(N107), .B2(net26499), .C1(N75), .C2(net26491), .A(n468), 
        .ZN(n469) );
  NAND3_X1 U750 ( .A1(n471), .A2(n470), .A3(n469), .ZN(RES[16]) );
  OAI222_X1 U751 ( .A1(n473), .A2(net24561), .B1(net26479), .B2(n47), .C1(n48), 
        .C2(net26700), .ZN(n475) );
  INV_X1 U752 ( .A(n475), .ZN(n476) );
  OAI21_X1 U753 ( .B1(n338), .B2(net18434), .A(n476), .ZN(n409) );
  NAND2_X1 U754 ( .A1(net31345), .A2(net31364), .ZN(n411) );
  OAI21_X1 U755 ( .B1(net18434), .B2(n728), .A(n476), .ZN(n408) );
  OAI21_X1 U756 ( .B1(n137), .B2(net26385), .A(net26407), .ZN(n477) );
  AOI221_X1 U757 ( .B1(n251), .B2(n712), .C1(n91), .C2(n477), .A(n660), .ZN(
        n495) );
  INV_X1 U758 ( .A(n411), .ZN(net24728) );
  MUX2_X1 U759 ( .A(net26387), .B(net26415), .S(n91), .Z(n479) );
  INV_X1 U760 ( .A(n137), .ZN(n478) );
  AOI21_X1 U761 ( .B1(n479), .B2(net26407), .A(n478), .ZN(n481) );
  AOI22_X1 U762 ( .A1(n153), .A2(net26423), .B1(net35295), .B2(net26435), .ZN(
        n486) );
  NAND3_X1 U763 ( .A1(n491), .A2(n490), .A3(n486), .ZN(n717) );
  AOI222_X1 U764 ( .A1(n212), .A2(n590), .B1(n686), .B2(n717), .C1(n255), .C2(
        n713), .ZN(n493) );
  AOI222_X1 U765 ( .A1(N76), .A2(net26493), .B1(n687), .B2(n711), .C1(N108), 
        .C2(net26501), .ZN(n492) );
  NAND4_X1 U766 ( .A1(n495), .A2(n494), .A3(n493), .A4(n492), .ZN(RES[17]) );
  OAI21_X1 U767 ( .B1(A[18]), .B2(net26387), .A(net26407), .ZN(n500) );
  AOI221_X1 U768 ( .B1(n251), .B2(n733), .C1(n105), .C2(n500), .A(n660), .ZN(
        n525) );
  AOI22_X1 U769 ( .A1(net35295), .A2(net26423), .B1(n34), .B2(n135), .ZN(n501)
         );
  NAND3_X1 U770 ( .A1(n505), .A2(n502), .A3(n501), .ZN(n738) );
  MUX2_X1 U771 ( .A(net26387), .B(net26415), .S(n105), .Z(n511) );
  INV_X1 U772 ( .A(A[18]), .ZN(n510) );
  AOI21_X1 U773 ( .B1(n511), .B2(net26407), .A(n510), .ZN(n514) );
  AOI221_X1 U774 ( .B1(n256), .B2(n267), .C1(n182), .C2(n738), .A(n514), .ZN(
        n517) );
  AOI222_X1 U775 ( .A1(n29), .A2(n606), .B1(n257), .B2(n266), .C1(n255), .C2(
        n734), .ZN(n516) );
  AOI222_X1 U776 ( .A1(N77), .A2(net26493), .B1(n687), .B2(n732), .C1(N109), 
        .C2(net26501), .ZN(n515) );
  NAND4_X1 U777 ( .A1(n525), .A2(n517), .A3(n516), .A4(n515), .ZN(RES[18]) );
  OAI211_X1 U778 ( .C1(n532), .C2(net24561), .A(n49), .B(n378), .ZN(n207) );
  MUX2_X1 U779 ( .A(n532), .B(net24439), .S(n274), .Z(n533) );
  OAI21_X1 U780 ( .B1(n30), .B2(n533), .A(n49), .ZN(n205) );
  OAI21_X1 U781 ( .B1(A[19]), .B2(net26387), .A(net26407), .ZN(n535) );
  AOI221_X1 U782 ( .B1(n251), .B2(net24464), .C1(B[19]), .C2(n535), .A(n660), 
        .ZN(n561) );
  AOI22_X1 U783 ( .A1(n34), .A2(net26425), .B1(n137), .B2(n135), .ZN(n546) );
  NAND3_X1 U784 ( .A1(n554), .A2(n548), .A3(n546), .ZN(net24457) );
  MUX2_X1 U785 ( .A(net26387), .B(net26415), .S(B[19]), .Z(n556) );
  INV_X1 U786 ( .A(A[19]), .ZN(n555) );
  AOI21_X1 U787 ( .B1(n556), .B2(net26407), .A(n555), .ZN(n557) );
  AOI221_X1 U788 ( .B1(n256), .B2(n207), .C1(n248), .C2(net24457), .A(n557), 
        .ZN(n560) );
  AOI222_X1 U789 ( .A1(n212), .A2(net24562), .B1(n257), .B2(n74), .C1(n255), 
        .C2(net24463), .ZN(n559) );
  NAND4_X1 U790 ( .A1(n558), .A2(n560), .A3(n559), .A4(n561), .ZN(RES[19]) );
  OAI21_X1 U791 ( .B1(n230), .B2(net26387), .A(net26407), .ZN(n565) );
  NOR2_X1 U792 ( .A1(n233), .A2(n562), .ZN(n564) );
  AOI22_X1 U793 ( .A1(n137), .A2(net26423), .B1(A[18]), .B2(net26437), .ZN(
        n566) );
  NAND3_X1 U794 ( .A1(n71), .A2(n567), .A3(n566), .ZN(n698) );
  MUX2_X1 U795 ( .A(net26387), .B(net26415), .S(B[20]), .Z(n570) );
  INV_X1 U796 ( .A(A[20]), .ZN(n569) );
  AOI21_X1 U797 ( .B1(n570), .B2(net26407), .A(n569), .ZN(n571) );
  AOI221_X1 U798 ( .B1(n246), .B2(n698), .C1(n257), .C2(n572), .A(n571), .ZN(
        n577) );
  AOI222_X1 U799 ( .A1(n29), .A2(n638), .B1(n256), .B2(n574), .C1(n255), .C2(
        n573), .ZN(n576) );
  AOI222_X1 U800 ( .A1(N79), .A2(net26491), .B1(n687), .B2(n639), .C1(N111), 
        .C2(net26501), .ZN(n575) );
  NAND4_X1 U801 ( .A1(n578), .A2(n577), .A3(n576), .A4(n575), .ZN(RES[20]) );
  INV_X1 U802 ( .A(A[21]), .ZN(n585) );
  AOI21_X1 U803 ( .B1(net26397), .B2(n585), .A(net31788), .ZN(n580) );
  INV_X1 U804 ( .A(n223), .ZN(n579) );
  OAI21_X1 U805 ( .B1(n580), .B2(n579), .A(n675), .ZN(n581) );
  AOI221_X1 U806 ( .B1(n250), .B2(n712), .C1(n251), .C2(n713), .A(n581), .ZN(
        n594) );
  AOI22_X1 U807 ( .A1(A[18]), .A2(net36181), .B1(A[19]), .B2(net26433), .ZN(
        n582) );
  NAND3_X1 U808 ( .A1(n584), .A2(n583), .A3(n582), .ZN(n718) );
  MUX2_X1 U809 ( .A(net26387), .B(net26415), .S(n223), .Z(n586) );
  AOI21_X1 U810 ( .B1(n586), .B2(net26407), .A(n585), .ZN(n587) );
  AOI222_X1 U811 ( .A1(n255), .A2(n590), .B1(n257), .B2(n589), .C1(n687), .C2(
        n717), .ZN(n592) );
  AOI222_X1 U812 ( .A1(N80), .A2(net26491), .B1(n212), .B2(n711), .C1(N112), 
        .C2(net26501), .ZN(n591) );
  NAND4_X1 U813 ( .A1(n594), .A2(n593), .A3(n592), .A4(n591), .ZN(RES[21]) );
  INV_X1 U814 ( .A(n167), .ZN(n601) );
  AOI21_X1 U815 ( .B1(net26397), .B2(n601), .A(net31788), .ZN(n596) );
  INV_X1 U816 ( .A(B[22]), .ZN(n595) );
  OAI21_X1 U817 ( .B1(n596), .B2(n595), .A(n675), .ZN(n597) );
  AOI221_X1 U818 ( .B1(n250), .B2(n733), .C1(n251), .C2(n734), .A(n597), .ZN(
        n610) );
  AOI22_X1 U819 ( .A1(A[19]), .A2(net36207), .B1(n230), .B2(net26437), .ZN(
        n598) );
  NAND3_X1 U820 ( .A1(n600), .A2(n599), .A3(n598), .ZN(n739) );
  MUX2_X1 U821 ( .A(net26387), .B(net26415), .S(B[22]), .Z(n602) );
  AOI21_X1 U822 ( .B1(n602), .B2(net26407), .A(n601), .ZN(n603) );
  AOI221_X1 U823 ( .B1(n687), .B2(n738), .C1(n246), .C2(n739), .A(n603), .ZN(
        n609) );
  NAND4_X1 U824 ( .A1(n610), .A2(n609), .A3(n608), .A4(n607), .ZN(RES[22]) );
  INV_X1 U825 ( .A(A[23]), .ZN(n617) );
  AOI21_X1 U826 ( .B1(net26397), .B2(n617), .A(net31788), .ZN(n612) );
  INV_X1 U827 ( .A(B[23]), .ZN(n611) );
  OAI21_X1 U828 ( .B1(n612), .B2(n611), .A(n675), .ZN(n613) );
  AOI22_X1 U829 ( .A1(n230), .A2(net26423), .B1(n24), .B2(net26437), .ZN(n614)
         );
  NAND3_X1 U830 ( .A1(n616), .A2(n615), .A3(n614), .ZN(net24456) );
  MUX2_X1 U831 ( .A(net26387), .B(net26415), .S(B[23]), .Z(n618) );
  AOI21_X1 U832 ( .B1(n618), .B2(net26407), .A(n617), .ZN(n619) );
  AOI222_X1 U833 ( .A1(n255), .A2(net24562), .B1(n256), .B2(n621), .C1(n257), 
        .C2(n620), .ZN(n623) );
  OAI222_X1 U834 ( .A1(n627), .A2(net26700), .B1(net26479), .B2(n697), .C1(
        net24561), .C2(n626), .ZN(n629) );
  OAI21_X1 U835 ( .B1(n169), .B2(net26385), .A(net26407), .ZN(n628) );
  AOI221_X1 U836 ( .B1(n678), .B2(n629), .C1(B[24]), .C2(n628), .A(n660), .ZN(
        n643) );
  AOI22_X1 U837 ( .A1(n24), .A2(net36181), .B1(n167), .B2(net26435), .ZN(n630)
         );
  NAND3_X1 U838 ( .A1(n632), .A2(n631), .A3(n630), .ZN(n699) );
  MUX2_X1 U839 ( .A(net26387), .B(net26415), .S(B[24]), .Z(n634) );
  INV_X1 U840 ( .A(n169), .ZN(n633) );
  AOI21_X1 U841 ( .B1(n634), .B2(net26407), .A(n633), .ZN(n635) );
  AOI222_X1 U842 ( .A1(n255), .A2(n638), .B1(n687), .B2(n698), .C1(n256), .C2(
        n637), .ZN(n641) );
  NAND4_X1 U843 ( .A1(n643), .A2(n642), .A3(n641), .A4(n640), .ZN(RES[24]) );
  OAI21_X1 U844 ( .B1(n33), .B2(net26387), .A(net26407), .ZN(n644) );
  AOI22_X1 U845 ( .A1(n167), .A2(net36207), .B1(A[23]), .B2(net26433), .ZN(
        n646) );
  NAND3_X1 U846 ( .A1(n648), .A2(n647), .A3(n646), .ZN(n719) );
  MUX2_X1 U847 ( .A(net26387), .B(net26415), .S(B[25]), .Z(n650) );
  INV_X1 U848 ( .A(A[25]), .ZN(n649) );
  AOI21_X1 U849 ( .B1(n650), .B2(net26407), .A(n649), .ZN(n651) );
  AOI221_X1 U850 ( .B1(n687), .B2(n718), .C1(n182), .C2(n719), .A(n651), .ZN(
        n656) );
  AOI222_X1 U851 ( .A1(N84), .A2(net26491), .B1(n255), .B2(n711), .C1(N116), 
        .C2(net26499), .ZN(n654) );
  NAND4_X1 U852 ( .A1(n657), .A2(n656), .A3(n655), .A4(n654), .ZN(RES[25]) );
  OAI222_X1 U853 ( .A1(n659), .A2(net26700), .B1(net26479), .B2(n736), .C1(
        n658), .C2(net24561), .ZN(n662) );
  OAI21_X1 U854 ( .B1(n154), .B2(net26385), .A(net26407), .ZN(n661) );
  AOI22_X1 U855 ( .A1(A[23]), .A2(net36181), .B1(n169), .B2(n135), .ZN(n663)
         );
  NAND3_X1 U856 ( .A1(n665), .A2(n664), .A3(n663), .ZN(n740) );
  MUX2_X1 U857 ( .A(net26387), .B(net26415), .S(n75), .Z(n667) );
  INV_X1 U858 ( .A(n154), .ZN(n666) );
  AOI21_X1 U859 ( .B1(n667), .B2(net26407), .A(n666), .ZN(n668) );
  AOI221_X1 U860 ( .B1(n182), .B2(n740), .C1(n257), .C2(n669), .A(n668), .ZN(
        n673) );
  AOI222_X1 U861 ( .A1(N85), .A2(net26491), .B1(n255), .B2(n732), .C1(N117), 
        .C2(net26499), .ZN(n671) );
  NAND4_X1 U862 ( .A1(n671), .A2(n673), .A3(n674), .A4(n672), .ZN(RES[26]) );
  OAI21_X1 U863 ( .B1(A[27]), .B2(net26387), .A(net26407), .ZN(n677) );
  NAND3_X1 U864 ( .A1(n256), .A2(A[31]), .A3(net26479), .ZN(n676) );
  AOI22_X1 U865 ( .A1(n169), .A2(net36207), .B1(n33), .B2(n135), .ZN(n679) );
  NAND3_X1 U866 ( .A1(n681), .A2(n680), .A3(n679), .ZN(net24458) );
  INV_X1 U867 ( .A(n682), .ZN(n685) );
  MUX2_X1 U868 ( .A(net26387), .B(net26415), .S(B[27]), .Z(n683) );
  AOI21_X1 U869 ( .B1(n683), .B2(net26403), .A(n760), .ZN(n684) );
  AOI221_X1 U870 ( .B1(n182), .B2(net24458), .C1(n685), .C2(n256), .A(n684), 
        .ZN(n691) );
  AOI222_X1 U871 ( .A1(n257), .A2(n688), .B1(n687), .B2(net24456), .C1(n29), 
        .C2(net24457), .ZN(n690) );
  NAND4_X1 U872 ( .A1(n689), .A2(n691), .A3(n690), .A4(n692), .ZN(RES[27]) );
  INV_X1 U873 ( .A(n693), .ZN(n694) );
  OAI21_X1 U874 ( .B1(n257), .B2(n256), .A(n694), .ZN(n710) );
  OAI21_X1 U875 ( .B1(A[28]), .B2(net26387), .A(net26407), .ZN(n705) );
  OAI222_X1 U876 ( .A1(n697), .A2(net26700), .B1(net26479), .B2(n696), .C1(n30), .C2(n695), .ZN(n703) );
  AOI22_X1 U877 ( .A1(net20298), .A2(n699), .B1(n213), .B2(n698), .ZN(n700) );
  OAI221_X1 U878 ( .B1(net18434), .B2(n701), .C1(n295), .C2(net26479), .A(n700), .ZN(n702) );
  MUX2_X1 U879 ( .A(n703), .B(n702), .S(net35873), .Z(n704) );
  AOI22_X1 U880 ( .A1(B[28]), .A2(n705), .B1(net32003), .B2(n704), .ZN(n709)
         );
  MUX2_X1 U881 ( .A(net26387), .B(net26415), .S(B[28]), .Z(n706) );
  AOI21_X1 U882 ( .B1(n706), .B2(net26407), .A(net19990), .ZN(n707) );
  AOI221_X1 U883 ( .B1(N87), .B2(net26493), .C1(N119), .C2(net26497), .A(n707), 
        .ZN(n708) );
  OAI21_X1 U884 ( .B1(A[29]), .B2(net26387), .A(net26407), .ZN(n726) );
  INV_X1 U885 ( .A(n711), .ZN(n716) );
  AOI22_X1 U886 ( .A1(n213), .A2(n713), .B1(n712), .B2(n232), .ZN(n714) );
  OAI221_X1 U887 ( .B1(net26479), .B2(n716), .C1(n715), .C2(net26700), .A(n714), .ZN(n723) );
  INV_X1 U888 ( .A(n717), .ZN(n721) );
  AOI22_X1 U889 ( .A1(net20298), .A2(n719), .B1(n213), .B2(n718), .ZN(n720) );
  OAI221_X1 U890 ( .B1(net18434), .B2(n721), .C1(n279), .C2(net26479), .A(n720), .ZN(n722) );
  MUX2_X1 U891 ( .A(n723), .B(n722), .S(net35873), .Z(n725) );
  NAND2_X1 U892 ( .A1(n256), .A2(net26485), .ZN(n745) );
  AOI221_X1 U893 ( .B1(B[29]), .B2(n726), .C1(net32003), .C2(n725), .A(n724), 
        .ZN(n731) );
  NAND2_X1 U894 ( .A1(n257), .A2(net26483), .ZN(net24440) );
  OAI21_X1 U895 ( .B1(net31788), .B2(net24497), .A(A[29]), .ZN(n727) );
  OAI21_X1 U896 ( .B1(n728), .B2(net24440), .A(n727), .ZN(n729) );
  AOI221_X1 U897 ( .B1(N120), .B2(net26499), .C1(N88), .C2(net26491), .A(n729), 
        .ZN(n730) );
  NAND2_X1 U898 ( .A1(n731), .A2(n730), .ZN(RES[29]) );
  OAI21_X1 U899 ( .B1(n77), .B2(net26387), .A(net26407), .ZN(n749) );
  INV_X1 U900 ( .A(n732), .ZN(n737) );
  AOI22_X1 U901 ( .A1(n213), .A2(n734), .B1(n733), .B2(n232), .ZN(n735) );
  OAI221_X1 U902 ( .B1(net26479), .B2(n737), .C1(n736), .C2(net26700), .A(n735), .ZN(n744) );
  INV_X1 U903 ( .A(n738), .ZN(n742) );
  AOI22_X1 U904 ( .A1(net20298), .A2(n740), .B1(n213), .B2(n739), .ZN(n741) );
  OAI221_X1 U905 ( .B1(net18434), .B2(n742), .C1(n247), .C2(net26479), .A(n741), .ZN(n743) );
  MUX2_X1 U906 ( .A(n744), .B(n743), .S(net35873), .Z(n748) );
  MUX2_X1 U907 ( .A(net26397), .B(net31778), .S(B[30]), .Z(n750) );
  OAI21_X1 U908 ( .B1(net31788), .B2(n750), .A(n77), .ZN(n751) );
  OAI21_X1 U909 ( .B1(n752), .B2(net24440), .A(n751), .ZN(n753) );
  NAND2_X1 U910 ( .A1(n754), .A2(n755), .ZN(RES[30]) );
  INV_X1 U911 ( .A(n412), .ZN(n782) );
  INV_X1 U912 ( .A(n407), .ZN(n775) );
  INV_X1 U913 ( .A(n269), .ZN(n781) );
  INV_X1 U914 ( .A(n265), .ZN(n774) );
  INV_X1 U915 ( .A(n756), .ZN(n254) );
  INV_X1 U916 ( .A(n211), .ZN(n780) );
  INV_X1 U917 ( .A(n204), .ZN(n773) );
  OR3_X1 U918 ( .A1(n158), .A2(B[15]), .A3(B[14]), .ZN(n765) );
  NOR4_X1 U919 ( .A1(n765), .A2(n103), .A3(n200), .A4(n201), .ZN(n772) );
  OR4_X1 U920 ( .A1(B[28]), .A2(B[26]), .A3(B[29]), .A4(B[27]), .ZN(n767) );
endmodule


module REG_PIPO_6_00_00_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n14), .ZN(n20) );
  INV_X1 U3 ( .A(n21), .ZN(n13) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n20), .B1(n14), .B2(DOUT[0]), .ZN(n21) );
  INV_X1 U5 ( .A(n19), .ZN(n12) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n20), .B1(n14), .B2(DOUT[1]), .ZN(n19) );
  INV_X1 U7 ( .A(n18), .ZN(n11) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n20), .B1(n14), .B2(DOUT[2]), .ZN(n18) );
  INV_X1 U9 ( .A(n17), .ZN(n10) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n20), .B1(n14), .B2(DOUT[3]), .ZN(n17) );
  INV_X1 U11 ( .A(n16), .ZN(n9) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n20), .B1(n14), .B2(DOUT[4]), .ZN(n16) );
  INV_X1 U13 ( .A(n15), .ZN(n3) );
  AOI22_X1 U14 ( .A1(DIN[5]), .A2(n20), .B1(n14), .B2(DOUT[5]), .ZN(n15) );
  INV_X1 U15 ( .A(EN), .ZN(n14) );
endmodule


module REG_PIPO_32_00000000_00000000_6 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_5 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n66, n98, net24417, net34753, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n67, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n98), .CK(CLK), .RN(n11), .Q(DOUT[31]), .QN(
        n66) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n105), .CK(CLK), .RN(n11), .Q(DOUT[30]), .QN(
        n135) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n106), .CK(CLK), .RN(n11), .Q(DOUT[29]), .QN(
        n136) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n107), .CK(CLK), .RN(n11), .Q(DOUT[28]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n108), .CK(CLK), .RN(n11), .Q(DOUT[27]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n109), .CK(CLK), .RN(n11), .Q(DOUT[26]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n110), .CK(CLK), .RN(n11), .Q(DOUT[25]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n111), .CK(CLK), .RN(n11), .Q(DOUT[24]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n112), .CK(CLK), .RN(n11), .Q(DOUT[23]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n113), .CK(CLK), .RN(n11), .Q(DOUT[22]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n114), .CK(CLK), .RN(n10), .Q(DOUT[21]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n115), .CK(CLK), .RN(n10), .Q(DOUT[20]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n116), .CK(CLK), .RN(n10), .Q(DOUT[19]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n117), .CK(CLK), .RN(n10), .Q(DOUT[18]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n118), .CK(CLK), .RN(n10), .Q(DOUT[17]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n119), .CK(CLK), .RN(n10), .Q(DOUT[16]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n120), .CK(CLK), .RN(n10), .Q(DOUT[15]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n121), .CK(CLK), .RN(n10), .Q(DOUT[14]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n122), .CK(CLK), .RN(n10), .Q(DOUT[13]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n123), .CK(CLK), .RN(n10), .Q(DOUT[12]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n124), .CK(CLK), .RN(n10), .Q(DOUT[11]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n125), .CK(CLK), .RN(n9), .Q(DOUT[10]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n126), .CK(CLK), .RN(n9), .Q(DOUT[9]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n127), .CK(CLK), .RN(n9), .Q(DOUT[8]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n128), .CK(CLK), .RN(n9), .Q(DOUT[7]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n129), .CK(CLK), .RN(n9), .Q(DOUT[6]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n130), .CK(CLK), .RN(n9), .Q(DOUT[5]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n131), .CK(CLK), .RN(n9), .Q(DOUT[4]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n132), .CK(CLK), .RN(n9), .Q(DOUT[3]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n133), .CK(CLK), .RN(n9), .Q(DOUT[2]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n134), .CK(CLK), .RN(n9), .Q(DOUT[1]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n5), .CK(CLK), .RN(n9), .Q(DOUT[0]), .QN(n165)
         );
  OR2_X1 U2 ( .A1(INIT), .A2(n7), .ZN(n1) );
  OR2_X1 U3 ( .A1(n142), .A2(EN), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n23), .A2(n2), .ZN(n112) );
  NAND2_X1 U5 ( .A1(DIN[0]), .A2(net24417), .ZN(n3) );
  OR2_X1 U6 ( .A1(n165), .A2(EN), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n3), .A2(n4), .ZN(n5) );
  INV_X2 U8 ( .A(n1), .ZN(net24417) );
  NAND2_X1 U9 ( .A1(n6), .A2(net34753), .ZN(n98) );
  OR2_X1 U10 ( .A1(n66), .A2(EN), .ZN(net34753) );
  NAND2_X1 U11 ( .A1(DIN[31]), .A2(net24417), .ZN(n6) );
  INV_X1 U12 ( .A(EN), .ZN(n7) );
  OR2_X1 U13 ( .A1(n138), .A2(EN), .ZN(n8) );
  NAND2_X1 U14 ( .A1(n27), .A2(n8), .ZN(n108) );
  BUF_X1 U15 ( .A(RST_AN), .Z(n9) );
  BUF_X1 U16 ( .A(RST_AN), .Z(n10) );
  BUF_X1 U17 ( .A(RST_AN), .Z(n11) );
  OAI22_X1 U18 ( .A1(n154), .A2(EN), .B1(n1), .B2(n31), .ZN(n124) );
  INV_X1 U19 ( .A(DIN[11]), .ZN(n31) );
  OAI22_X1 U20 ( .A1(n160), .A2(EN), .B1(n1), .B2(n100), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[5]), .ZN(n100) );
  OAI22_X1 U22 ( .A1(n159), .A2(EN), .B1(n1), .B2(n99), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[6]), .ZN(n99) );
  OAI22_X1 U24 ( .A1(n162), .A2(EN), .B1(n1), .B2(n102), .ZN(n132) );
  INV_X1 U25 ( .A(DIN[3]), .ZN(n102) );
  OAI22_X1 U26 ( .A1(n164), .A2(EN), .B1(n1), .B2(n104), .ZN(n134) );
  INV_X1 U27 ( .A(DIN[1]), .ZN(n104) );
  OAI22_X1 U28 ( .A1(n163), .A2(EN), .B1(n103), .B2(n1), .ZN(n133) );
  INV_X1 U29 ( .A(DIN[2]), .ZN(n103) );
  OAI22_X1 U30 ( .A1(n155), .A2(EN), .B1(n1), .B2(n32), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[10]), .ZN(n32) );
  OAI22_X1 U32 ( .A1(n161), .A2(EN), .B1(n1), .B2(n101), .ZN(n131) );
  INV_X1 U33 ( .A(DIN[4]), .ZN(n101) );
  OAI22_X1 U34 ( .A1(n156), .A2(EN), .B1(n1), .B2(n33), .ZN(n126) );
  INV_X1 U35 ( .A(DIN[9]), .ZN(n33) );
  OAI22_X1 U36 ( .A1(n157), .A2(EN), .B1(n1), .B2(n34), .ZN(n127) );
  INV_X1 U37 ( .A(DIN[8]), .ZN(n34) );
  OAI22_X1 U38 ( .A1(n158), .A2(EN), .B1(n1), .B2(n67), .ZN(n128) );
  INV_X1 U39 ( .A(DIN[7]), .ZN(n67) );
  NAND2_X1 U40 ( .A1(DIN[12]), .A2(net24417), .ZN(n12) );
  OAI21_X1 U41 ( .B1(n153), .B2(EN), .A(n12), .ZN(n123) );
  NAND2_X1 U42 ( .A1(DIN[13]), .A2(net24417), .ZN(n13) );
  OAI21_X1 U43 ( .B1(n152), .B2(EN), .A(n13), .ZN(n122) );
  NAND2_X1 U44 ( .A1(DIN[14]), .A2(net24417), .ZN(n14) );
  OAI21_X1 U45 ( .B1(n151), .B2(EN), .A(n14), .ZN(n121) );
  NAND2_X1 U46 ( .A1(DIN[15]), .A2(net24417), .ZN(n15) );
  OAI21_X1 U47 ( .B1(n150), .B2(EN), .A(n15), .ZN(n120) );
  NAND2_X1 U48 ( .A1(DIN[16]), .A2(net24417), .ZN(n16) );
  OAI21_X1 U49 ( .B1(n149), .B2(EN), .A(n16), .ZN(n119) );
  NAND2_X1 U50 ( .A1(DIN[17]), .A2(net24417), .ZN(n17) );
  OAI21_X1 U51 ( .B1(n148), .B2(EN), .A(n17), .ZN(n118) );
  NAND2_X1 U52 ( .A1(DIN[18]), .A2(net24417), .ZN(n18) );
  OAI21_X1 U53 ( .B1(n147), .B2(EN), .A(n18), .ZN(n117) );
  NAND2_X1 U54 ( .A1(DIN[19]), .A2(net24417), .ZN(n19) );
  OAI21_X1 U55 ( .B1(n146), .B2(EN), .A(n19), .ZN(n116) );
  NAND2_X1 U56 ( .A1(DIN[20]), .A2(net24417), .ZN(n20) );
  OAI21_X1 U57 ( .B1(n145), .B2(EN), .A(n20), .ZN(n115) );
  NAND2_X1 U58 ( .A1(DIN[21]), .A2(net24417), .ZN(n21) );
  OAI21_X1 U59 ( .B1(n144), .B2(EN), .A(n21), .ZN(n114) );
  NAND2_X1 U60 ( .A1(DIN[22]), .A2(net24417), .ZN(n22) );
  OAI21_X1 U61 ( .B1(n143), .B2(EN), .A(n22), .ZN(n113) );
  NAND2_X1 U62 ( .A1(DIN[23]), .A2(net24417), .ZN(n23) );
  NAND2_X1 U63 ( .A1(DIN[24]), .A2(net24417), .ZN(n24) );
  OAI21_X1 U64 ( .B1(n141), .B2(EN), .A(n24), .ZN(n111) );
  NAND2_X1 U65 ( .A1(DIN[25]), .A2(net24417), .ZN(n25) );
  OAI21_X1 U66 ( .B1(n140), .B2(EN), .A(n25), .ZN(n110) );
  NAND2_X1 U67 ( .A1(DIN[26]), .A2(net24417), .ZN(n26) );
  OAI21_X1 U68 ( .B1(n139), .B2(EN), .A(n26), .ZN(n109) );
  NAND2_X1 U69 ( .A1(DIN[27]), .A2(net24417), .ZN(n27) );
  NAND2_X1 U70 ( .A1(DIN[28]), .A2(net24417), .ZN(n28) );
  OAI21_X1 U71 ( .B1(n137), .B2(EN), .A(n28), .ZN(n107) );
  NAND2_X1 U72 ( .A1(DIN[29]), .A2(net24417), .ZN(n29) );
  OAI21_X1 U73 ( .B1(n136), .B2(EN), .A(n29), .ZN(n106) );
  NAND2_X1 U74 ( .A1(DIN[30]), .A2(net24417), .ZN(n30) );
  OAI21_X1 U75 ( .B1(n135), .B2(EN), .A(n30), .ZN(n105) );
endmodule


module REG_PIPO_32_00000000_00000000_4 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_5_00_00_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(n11) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  INV_X1 U5 ( .A(n16), .ZN(n10) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  INV_X1 U9 ( .A(n14), .ZN(n8) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  INV_X1 U11 ( .A(n13), .ZN(n3) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  INV_X1 U13 ( .A(EN), .ZN(n12) );
endmodule


module REG_PIPO_1_0_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [0:0] DIN;
  output [0:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n3, n4, n2;

  DFFR_X1 \reg_mem_reg[0]  ( .D(n4), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]), .QN(
        n3) );
  NAND3_X1 U3 ( .A1(DIN[0]), .A2(n2), .A3(EN), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n4) );
  INV_X1 U4 ( .A(INIT), .ZN(n2) );
endmodule


module REG_PIPO_32_00000000_00000000_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n168), .A2(EN), .B1(n2), .B2(n103), .ZN(n136) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n103) );
  OAI22_X1 U10 ( .A1(n167), .A2(EN), .B1(n2), .B2(n102), .ZN(n135) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n102) );
  OAI22_X1 U12 ( .A1(n166), .A2(EN), .B1(n2), .B2(n101), .ZN(n134) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n101) );
  OAI22_X1 U14 ( .A1(n165), .A2(EN), .B1(n2), .B2(n100), .ZN(n133) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n100) );
  OAI22_X1 U16 ( .A1(n164), .A2(EN), .B1(n2), .B2(n99), .ZN(n132) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n99) );
  OAI22_X1 U18 ( .A1(n163), .A2(EN), .B1(n2), .B2(n34), .ZN(n131) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n34) );
  OAI22_X1 U20 ( .A1(n162), .A2(EN), .B1(n2), .B2(n33), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n33) );
  OAI22_X1 U22 ( .A1(n161), .A2(EN), .B1(n2), .B2(n32), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n160), .A2(EN), .B1(n2), .B2(n31), .ZN(n128) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n159), .A2(EN), .B1(n2), .B2(n30), .ZN(n127) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n158), .A2(EN), .B1(n2), .B2(n29), .ZN(n126) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n29) );
  OAI22_X1 U30 ( .A1(n157), .A2(EN), .B1(n3), .B2(n28), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n28) );
  OAI22_X1 U32 ( .A1(n156), .A2(EN), .B1(n3), .B2(n27), .ZN(n124) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n27) );
  OAI22_X1 U34 ( .A1(n155), .A2(EN), .B1(n3), .B2(n26), .ZN(n123) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n154), .A2(EN), .B1(n3), .B2(n25), .ZN(n122) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n25) );
  OAI22_X1 U38 ( .A1(n153), .A2(EN), .B1(n3), .B2(n24), .ZN(n121) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n24) );
  OAI22_X1 U40 ( .A1(n152), .A2(EN), .B1(n3), .B2(n23), .ZN(n120) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n151), .A2(EN), .B1(n3), .B2(n22), .ZN(n119) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n22) );
  OAI22_X1 U44 ( .A1(n150), .A2(EN), .B1(n3), .B2(n21), .ZN(n118) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n21) );
  OAI22_X1 U46 ( .A1(n149), .A2(EN), .B1(n3), .B2(n20), .ZN(n117) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n20) );
  OAI22_X1 U48 ( .A1(n148), .A2(EN), .B1(n3), .B2(n19), .ZN(n116) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n19) );
  OAI22_X1 U50 ( .A1(n147), .A2(EN), .B1(n3), .B2(n18), .ZN(n115) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n18) );
  OAI22_X1 U52 ( .A1(n146), .A2(EN), .B1(n4), .B2(n17), .ZN(n114) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n17) );
  OAI22_X1 U54 ( .A1(n145), .A2(EN), .B1(n4), .B2(n16), .ZN(n113) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n16) );
  OAI22_X1 U56 ( .A1(n144), .A2(EN), .B1(n4), .B2(n15), .ZN(n112) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n15) );
  OAI22_X1 U58 ( .A1(n143), .A2(EN), .B1(n4), .B2(n14), .ZN(n111) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n14) );
  OAI22_X1 U60 ( .A1(n142), .A2(EN), .B1(n4), .B2(n13), .ZN(n110) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n13) );
  OAI22_X1 U62 ( .A1(n141), .A2(EN), .B1(n4), .B2(n12), .ZN(n109) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n12) );
  OAI22_X1 U64 ( .A1(n140), .A2(EN), .B1(n4), .B2(n11), .ZN(n108) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n11) );
  OAI22_X1 U66 ( .A1(n139), .A2(EN), .B1(n4), .B2(n10), .ZN(n107) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n10) );
  OAI22_X1 U68 ( .A1(n138), .A2(EN), .B1(n4), .B2(n9), .ZN(n106) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n9) );
  OAI22_X1 U70 ( .A1(n137), .A2(EN), .B1(n4), .B2(n8), .ZN(n105) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n8) );
  NAND2_X1 U72 ( .A1(n104), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n168), .A2(EN), .B1(n2), .B2(n103), .ZN(n136) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n103) );
  OAI22_X1 U10 ( .A1(n167), .A2(EN), .B1(n2), .B2(n102), .ZN(n135) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n102) );
  OAI22_X1 U12 ( .A1(n166), .A2(EN), .B1(n2), .B2(n101), .ZN(n134) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n101) );
  OAI22_X1 U14 ( .A1(n165), .A2(EN), .B1(n2), .B2(n100), .ZN(n133) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n100) );
  OAI22_X1 U16 ( .A1(n164), .A2(EN), .B1(n2), .B2(n99), .ZN(n132) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n99) );
  OAI22_X1 U18 ( .A1(n163), .A2(EN), .B1(n2), .B2(n34), .ZN(n131) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n34) );
  OAI22_X1 U20 ( .A1(n162), .A2(EN), .B1(n2), .B2(n33), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n33) );
  OAI22_X1 U22 ( .A1(n161), .A2(EN), .B1(n2), .B2(n32), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n160), .A2(EN), .B1(n2), .B2(n31), .ZN(n128) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n159), .A2(EN), .B1(n2), .B2(n30), .ZN(n127) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n158), .A2(EN), .B1(n2), .B2(n29), .ZN(n126) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n29) );
  OAI22_X1 U30 ( .A1(n157), .A2(EN), .B1(n3), .B2(n28), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n28) );
  OAI22_X1 U32 ( .A1(n156), .A2(EN), .B1(n3), .B2(n27), .ZN(n124) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n27) );
  OAI22_X1 U34 ( .A1(n155), .A2(EN), .B1(n3), .B2(n26), .ZN(n123) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n154), .A2(EN), .B1(n3), .B2(n25), .ZN(n122) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n25) );
  OAI22_X1 U38 ( .A1(n153), .A2(EN), .B1(n3), .B2(n24), .ZN(n121) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n24) );
  OAI22_X1 U40 ( .A1(n152), .A2(EN), .B1(n3), .B2(n23), .ZN(n120) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n151), .A2(EN), .B1(n3), .B2(n22), .ZN(n119) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n22) );
  OAI22_X1 U44 ( .A1(n150), .A2(EN), .B1(n3), .B2(n21), .ZN(n118) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n21) );
  OAI22_X1 U46 ( .A1(n149), .A2(EN), .B1(n3), .B2(n20), .ZN(n117) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n20) );
  OAI22_X1 U48 ( .A1(n148), .A2(EN), .B1(n3), .B2(n19), .ZN(n116) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n19) );
  OAI22_X1 U50 ( .A1(n147), .A2(EN), .B1(n3), .B2(n18), .ZN(n115) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n18) );
  OAI22_X1 U52 ( .A1(n146), .A2(EN), .B1(n4), .B2(n17), .ZN(n114) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n17) );
  OAI22_X1 U54 ( .A1(n145), .A2(EN), .B1(n4), .B2(n16), .ZN(n113) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n16) );
  OAI22_X1 U56 ( .A1(n144), .A2(EN), .B1(n4), .B2(n15), .ZN(n112) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n15) );
  OAI22_X1 U58 ( .A1(n143), .A2(EN), .B1(n4), .B2(n14), .ZN(n111) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n14) );
  OAI22_X1 U60 ( .A1(n142), .A2(EN), .B1(n4), .B2(n13), .ZN(n110) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n13) );
  OAI22_X1 U62 ( .A1(n141), .A2(EN), .B1(n4), .B2(n12), .ZN(n109) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n12) );
  OAI22_X1 U64 ( .A1(n140), .A2(EN), .B1(n4), .B2(n11), .ZN(n108) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n11) );
  OAI22_X1 U66 ( .A1(n139), .A2(EN), .B1(n4), .B2(n10), .ZN(n107) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n10) );
  OAI22_X1 U68 ( .A1(n138), .A2(EN), .B1(n4), .B2(n9), .ZN(n106) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n9) );
  OAI22_X1 U70 ( .A1(n137), .A2(EN), .B1(n4), .B2(n8), .ZN(n105) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n8) );
  NAND2_X1 U72 ( .A1(n104), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U10 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U12 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U14 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U16 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U18 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U20 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U22 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U24 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U28 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U30 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U32 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U34 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U36 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U38 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U42 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U44 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U46 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U48 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U50 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n19) );
  OAI22_X1 U52 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U54 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U56 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U58 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U60 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U62 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U64 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U66 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U68 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U70 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n9) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_5_00_00_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  INV_X1 U2 ( .A(n18), .ZN(n11) );
  AOI22_X1 U3 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  INV_X1 U4 ( .A(n16), .ZN(n10) );
  AOI22_X1 U5 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  INV_X1 U6 ( .A(n15), .ZN(n9) );
  AOI22_X1 U7 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  INV_X1 U8 ( .A(n14), .ZN(n8) );
  AOI22_X1 U9 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  INV_X1 U10 ( .A(n13), .ZN(n3) );
  AOI22_X1 U11 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  INV_X1 U12 ( .A(EN), .ZN(n12) );
  NOR2_X1 U13 ( .A1(INIT), .A2(n12), .ZN(n17) );
endmodule


module DATAPATH_DW01_add_2 ( A, B, CI, SUM, CO );
  input [30:0] A;
  input [30:0] B;
  output [30:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X1 U2 ( .A1(n1), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n35), .A2(n36), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n33), .A2(n34), .ZN(n2) );
  XOR2_X1 U5 ( .A(A[11]), .B(n3), .Z(SUM[11]) );
  NOR2_X1 U6 ( .A1(n7), .A2(n45), .ZN(n3) );
  XNOR2_X1 U7 ( .A(n4), .B(A[23]), .ZN(SUM[23]) );
  NAND2_X1 U8 ( .A1(A[22]), .A2(n10), .ZN(n4) );
  XOR2_X1 U9 ( .A(n24), .B(A[24]), .Z(SUM[24]) );
  XOR2_X1 U10 ( .A(n19), .B(A[28]), .Z(SUM[28]) );
  XNOR2_X1 U11 ( .A(n5), .B(A[27]), .ZN(SUM[27]) );
  NAND2_X1 U12 ( .A1(A[26]), .A2(n12), .ZN(n5) );
  XNOR2_X1 U13 ( .A(n6), .B(A[30]), .ZN(SUM[30]) );
  NAND2_X1 U14 ( .A1(n11), .A2(A[29]), .ZN(n6) );
  XOR2_X1 U15 ( .A(n13), .B(n49), .Z(SUM[9]) );
  XOR2_X1 U16 ( .A(n7), .B(n45), .Z(SUM[10]) );
  NOR2_X1 U17 ( .A1(n47), .A2(n39), .ZN(n14) );
  NOR2_X1 U18 ( .A1(n44), .A2(n36), .ZN(n43) );
  OR2_X1 U19 ( .A1(n49), .A2(n13), .ZN(n7) );
  INV_X1 U20 ( .A(n25), .ZN(n27) );
  INV_X1 U21 ( .A(n29), .ZN(n32) );
  INV_X1 U22 ( .A(n20), .ZN(n23) );
  NAND2_X1 U23 ( .A1(n37), .A2(n38), .ZN(n35) );
  XOR2_X1 U24 ( .A(A[5]), .B(n17), .Z(SUM[5]) );
  XOR2_X1 U25 ( .A(A[13]), .B(n42), .Z(SUM[13]) );
  XOR2_X1 U26 ( .A(A[8]), .B(n14), .Z(SUM[8]) );
  AND2_X1 U27 ( .A1(n42), .A2(A[13]), .ZN(n41) );
  AND2_X1 U28 ( .A1(n17), .A2(A[5]), .ZN(n16) );
  XOR2_X1 U29 ( .A(A[20]), .B(n28), .Z(SUM[20]) );
  NAND4_X1 U30 ( .A1(A[11]), .A2(A[10]), .A3(A[9]), .A4(A[8]), .ZN(n36) );
  NOR2_X1 U31 ( .A1(n29), .A2(n30), .ZN(n28) );
  XNOR2_X1 U32 ( .A(n40), .B(A[15]), .ZN(SUM[15]) );
  NAND2_X1 U33 ( .A1(n41), .A2(A[14]), .ZN(n40) );
  XNOR2_X1 U34 ( .A(A[3]), .B(SUM[2]), .ZN(SUM[3]) );
  XNOR2_X1 U35 ( .A(n15), .B(A[7]), .ZN(SUM[7]) );
  NAND2_X1 U36 ( .A1(n16), .A2(A[6]), .ZN(n15) );
  XOR2_X1 U37 ( .A(A[14]), .B(n41), .Z(SUM[14]) );
  XOR2_X1 U38 ( .A(A[6]), .B(n16), .Z(SUM[6]) );
  XOR2_X1 U39 ( .A(A[12]), .B(n43), .Z(SUM[12]) );
  XOR2_X1 U40 ( .A(A[17]), .B(n32), .Z(SUM[17]) );
  XOR2_X1 U41 ( .A(A[4]), .B(n38), .Z(SUM[4]) );
  XOR2_X1 U42 ( .A(n8), .B(A[16]), .Z(SUM[16]) );
  NOR2_X1 U43 ( .A1(SUM[2]), .A2(n48), .ZN(n38) );
  NAND4_X1 U44 ( .A1(A[4]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n39) );
  NOR2_X1 U45 ( .A1(n25), .A2(n26), .ZN(n24) );
  AND2_X1 U46 ( .A1(A[12]), .A2(n43), .ZN(n42) );
  NOR2_X1 U47 ( .A1(n46), .A2(n47), .ZN(n17) );
  XOR2_X1 U48 ( .A(A[21]), .B(n27), .Z(SUM[21]) );
  XOR2_X1 U49 ( .A(A[18]), .B(n9), .Z(SUM[18]) );
  XOR2_X1 U50 ( .A(n10), .B(A[22]), .Z(SUM[22]) );
  XOR2_X1 U51 ( .A(n23), .B(A[25]), .Z(SUM[25]) );
  XNOR2_X1 U52 ( .A(n31), .B(A[19]), .ZN(SUM[19]) );
  NAND2_X1 U53 ( .A1(n9), .A2(A[18]), .ZN(n31) );
  XOR2_X1 U54 ( .A(n11), .B(A[29]), .Z(SUM[29]) );
  XNOR2_X1 U55 ( .A(n12), .B(n22), .ZN(SUM[26]) );
  NOR2_X1 U56 ( .A1(n20), .A2(n21), .ZN(n19) );
  NAND2_X1 U57 ( .A1(n8), .A2(A[16]), .ZN(n29) );
  NAND2_X1 U58 ( .A1(n28), .A2(A[20]), .ZN(n25) );
  NAND2_X1 U59 ( .A1(n24), .A2(A[24]), .ZN(n20) );
  NAND2_X1 U60 ( .A1(n14), .A2(A[8]), .ZN(n13) );
  AND2_X1 U61 ( .A1(A[17]), .A2(n32), .ZN(n9) );
  AND2_X1 U62 ( .A1(A[21]), .A2(n27), .ZN(n10) );
  AND2_X1 U63 ( .A1(n19), .A2(A[28]), .ZN(n11) );
  NAND2_X1 U64 ( .A1(A[12]), .A2(A[13]), .ZN(n34) );
  AND2_X1 U65 ( .A1(A[25]), .A2(n23), .ZN(n12) );
  NAND2_X1 U66 ( .A1(A[14]), .A2(A[15]), .ZN(n33) );
  INV_X1 U67 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U68 ( .A(A[4]), .ZN(n46) );
  INV_X1 U69 ( .A(A[9]), .ZN(n49) );
  INV_X1 U70 ( .A(A[3]), .ZN(n48) );
  INV_X1 U71 ( .A(A[26]), .ZN(n22) );
  NAND3_X1 U72 ( .A1(A[26]), .A2(A[27]), .A3(A[25]), .ZN(n21) );
  NAND3_X1 U73 ( .A1(A[22]), .A2(A[23]), .A3(A[21]), .ZN(n26) );
  NAND3_X1 U74 ( .A1(A[18]), .A2(A[19]), .A3(A[17]), .ZN(n30) );
  INV_X1 U75 ( .A(n39), .ZN(n37) );
  INV_X1 U76 ( .A(n14), .ZN(n44) );
  INV_X1 U77 ( .A(A[10]), .ZN(n45) );
  INV_X1 U78 ( .A(n38), .ZN(n47) );
endmodule


module DATAPATH ( CLK, RST_AN, .CTRL_WORD({\CTRL_WORD[J_TYPE_IMM_SEL] , 
        \CTRL_WORD[R_TYPE_SEL] , \CTRL_WORD[IMM_SEL] , 
        \CTRL_WORD[PC_PLS_4_SEL] , \CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] , \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }), INSTR_CU, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .DP_SIG({
        \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] , 
        \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] , 
        \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] , 
        \DP_SIG[INSTR_OPCODE_M][0] }), IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] INSTR_CU;
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN, \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] , \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  wire   \npc_f[31] , n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n162, n163, n164, n165,
         n166, n167, n169, n170, n172, n184, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n277, n278, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n291, n302, net17718, net17723,
         net25305, net32890, net32889, net34337, net34366, net35180, net35179,
         net35178, net35228, net34800, net37560, n1, n2, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n160, n161, n168, n171, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n238, n239;
  wire   [30:0] pc_pls_4_f;
  wire   [31:0] pc_pls_4_d;
  wire   [31:0] instr_d;
  wire   [4:0] rf_waddr_d;
  wire   [31:0] rf_dout1_d;
  wire   [31:0] rf_dout2_d;
  wire   [4:0] rf_waddr_wb;
  wire   [31:16] imm_d;
  wire   [5:0] instr_opcode_e;
  wire   [31:0] pc_pls_4_e;
  wire   [31:0] rf_dout1_e;
  wire   [31:0] rf_dout2_e;
  wire   [31:0] imm_e;
  wire   [4:0] rs2_e;
  wire   [4:0] rs3_e;
  wire   [31:0] alu_a_e;
  wire   [31:0] alu_out_e;
  wire   [31:0] pc_pls_4_m;
  wire   [4:0] rf_waddr_m;
  wire   [31:0] pc_pls_4_wb;
  wire   [31:0] alu_out_wb;
  wire   [31:0] dmem_dout_wb;
  assign INSTR_CU[31] = IMEM_DOUT[31];
  assign INSTR_CU[30] = IMEM_DOUT[30];
  assign INSTR_CU[29] = IMEM_DOUT[29];
  assign INSTR_CU[28] = IMEM_DOUT[28];
  assign INSTR_CU[27] = IMEM_DOUT[27];
  assign INSTR_CU[26] = IMEM_DOUT[26];
  assign INSTR_CU[25] = IMEM_DOUT[25];
  assign INSTR_CU[24] = IMEM_DOUT[24];
  assign INSTR_CU[23] = IMEM_DOUT[23];
  assign INSTR_CU[22] = IMEM_DOUT[22];
  assign INSTR_CU[21] = IMEM_DOUT[21];
  assign INSTR_CU[20] = IMEM_DOUT[20];
  assign INSTR_CU[19] = IMEM_DOUT[19];
  assign INSTR_CU[18] = IMEM_DOUT[18];
  assign INSTR_CU[17] = IMEM_DOUT[17];
  assign INSTR_CU[16] = IMEM_DOUT[16];
  assign INSTR_CU[15] = IMEM_DOUT[15];
  assign INSTR_CU[14] = IMEM_DOUT[14];
  assign INSTR_CU[13] = IMEM_DOUT[13];
  assign INSTR_CU[12] = IMEM_DOUT[12];
  assign INSTR_CU[11] = IMEM_DOUT[11];
  assign INSTR_CU[10] = IMEM_DOUT[10];
  assign INSTR_CU[9] = IMEM_DOUT[9];
  assign INSTR_CU[8] = IMEM_DOUT[8];
  assign INSTR_CU[7] = IMEM_DOUT[7];
  assign INSTR_CU[6] = IMEM_DOUT[6];
  assign INSTR_CU[5] = IMEM_DOUT[5];
  assign INSTR_CU[4] = IMEM_DOUT[4];
  assign INSTR_CU[3] = IMEM_DOUT[3];
  assign INSTR_CU[2] = IMEM_DOUT[2];
  assign INSTR_CU[1] = IMEM_DOUT[1];
  assign INSTR_CU[0] = IMEM_DOUT[0];

  OR2_X2 U14 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[2]), .ZN(
        rf_waddr_d[2]) );
  OR2_X2 U15 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[1]), .ZN(
        rf_waddr_d[1]) );
  OR2_X2 U16 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[0]), .ZN(
        rf_waddr_d[0]) );
  OAI21_X2 U174 ( .B1(n86), .B2(n132), .A(n282), .ZN(alu_a_e[27]) );
  OAI21_X2 U182 ( .B1(n86), .B2(n136), .A(n286), .ZN(alu_a_e[23]) );
  REG_PIPO_32_fffffffc_fffffffc U_PC_REG ( .CLK(CLK), .RST_AN(n90), .EN(1'b1), 
        .INIT(1'b0), .DIN({\npc_f[31] , n93, n94, n95, n96, n97, n98, n99, 
        n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
        n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n197}), .DOUT(IMEM_ADDR) );
  REG_PIPO_32_00000000_00000000_0 U_PC_PLS_4_REG_FD ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN({1'b0, pc_pls_4_f}), 
        .DOUT(pc_pls_4_d) );
  REG_PIPO_32_00000000_00000000_11 U_INSTR_REG_FD ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN(IMEM_DOUT), .DOUT(instr_d) );
  RF_ADDR_W5_DATA_W32 U_RF ( .CLK(CLK), .RST_AN(n89), .ENABLE(1'b1), .RD1(1'b1), .RD2(1'b1), .WR(\CTRL_WORD[RF_WEN] ), .ADD_WR(rf_waddr_d), .ADD_RD1(
        instr_d[25:21]), .ADD_RD2(instr_d[20:16]), .DATAIN({n198, n199, n7, 
        n200, n201, n202, n203, n204, n205, n8, n206, n207, n208, n10, n26, 
        n12, n23, n24, n13, n25, n35, n36, n209, n210, n211, n212, n213, n214, 
        n215, n6, n9, n38}), .OUT1(rf_dout1_d), .OUT2(rf_dout2_d) );
  REG_PIPO_6_00_00_0 U_INSTR_OPCODE_REG_DE ( .CLK(CLK), .RST_AN(n89), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[31:26]), .DOUT(instr_opcode_e) );
  REG_PIPO_32_00000000_00000000_10 U_PC_PLS_4_REG_DE ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(pc_pls_4_d), .DOUT(
        pc_pls_4_e) );
  REG_PIPO_32_00000000_00000000_9 U_RF_DOUT1_REG_DE ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout1_d), .DOUT(
        rf_dout1_e) );
  REG_PIPO_32_00000000_00000000_8 U_RF_DOUT2_REG_DE ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout2_d), .DOUT(
        rf_dout2_e) );
  REG_PIPO_32_00000000_00000000_7 U_IMM_REG_DE ( .CLK(CLK), .RST_AN(n90), .EN(
        1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN({imm_d[31], imm_d[31], 
        imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[24:16], 
        instr_d[15:0]}), .DOUT(imm_e) );
  REG_PIPO_5_00_00_0 U_RS2_REG_DE ( .CLK(CLK), .RST_AN(n89), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[20:16]), .DOUT(rs2_e) );
  REG_PIPO_5_00_00_3 U_RS3_REG_DE ( .CLK(CLK), .RST_AN(n89), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[15:11]), .DOUT(rs3_e) );
  ALU_DATA_W32 U_ALU ( .FUNC({\CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] }), .A(alu_a_e), .B({n141, n142, n143, n160, 
        n161, n168, n171, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
        n182, n183, n185, n186, n187, n188, n189, n190, n191, net17723, n192, 
        n193, n194, n195, net17718, n196}), .RES(alu_out_e) );
  REG_PIPO_6_00_00_1 U_INSTR_OPCODE_REG_EM ( .CLK(CLK), .RST_AN(n89), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(instr_opcode_e), .DOUT({
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }) );
  REG_PIPO_32_00000000_00000000_6 U_PC_PLS_4_REG_EM ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(pc_pls_4_e), .DOUT(
        pc_pls_4_m) );
  REG_PIPO_32_00000000_00000000_5 U_ALU_OUT_REG_EM ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(alu_out_e), .DOUT(
        DMEM_RWADDR) );
  REG_PIPO_32_00000000_00000000_4 U_DMEM_DOUT_REG_EM ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(rf_dout2_e), .DOUT(
        DMEM_DIN) );
  REG_PIPO_5_00_00_2 U_RF_WADDR_REG_EM ( .CLK(CLK), .RST_AN(n89), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN({n123, n124, n125, n126, n127}), 
        .DOUT(rf_waddr_m) );
  REG_PIPO_1_0_0 U_IS_0_REG_EM ( .CLK(CLK), .RST_AN(n90), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_EM] ), .DIN(n302), .DOUT(\DP_SIG[CMPR_0_IS_0_M] ) );
  REG_PIPO_32_00000000_00000000_3 U_PC_PLS_4_REG_MWB ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(pc_pls_4_m), .DOUT(
        pc_pls_4_wb) );
  REG_PIPO_32_00000000_00000000_2 U_ALU_OUT_REG_MWB ( .CLK(CLK), .RST_AN(n90), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_RWADDR), .DOUT(
        alu_out_wb) );
  REG_PIPO_32_00000000_00000000_1 U_DMEM_DOUT_REG_MWB ( .CLK(CLK), .RST_AN(n90), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_DOUT), .DOUT(dmem_dout_wb) );
  REG_PIPO_5_00_00_1 U_RF_WADDR_REG_MWB ( .CLK(CLK), .RST_AN(n89), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(rf_waddr_m), .DOUT(rf_waddr_wb) );
  DATAPATH_DW01_add_2 add_242 ( .A(IMEM_ADDR[30:0]), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_pls_4_f) );
  BUF_X2 U5 ( .A(n2), .Z(n29) );
  BUF_X2 U7 ( .A(n2), .Z(n76) );
  BUF_X1 U8 ( .A(n151), .Z(n1) );
  BUF_X2 U9 ( .A(n150), .Z(n81) );
  NOR2_X1 U10 ( .A1(n239), .A2(n82), .ZN(n2) );
  BUF_X1 U11 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n72) );
  OAI21_X2 U12 ( .B1(n11), .B2(n128), .A(n277), .ZN(alu_a_e[31]) );
  NAND2_X1 U13 ( .A1(n37), .A2(n288), .ZN(alu_a_e[21]) );
  OAI21_X1 U17 ( .B1(n86), .B2(n134), .A(n284), .ZN(alu_a_e[25]) );
  NAND3_X1 U18 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n6) );
  NAND3_X1 U19 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n7) );
  NAND3_X1 U20 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n8) );
  CLKBUF_X1 U21 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n33) );
  CLKBUF_X1 U22 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n84) );
  OR3_X2 U23 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n9) );
  OR3_X2 U24 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n10) );
  BUF_X2 U25 ( .A(n72), .Z(n86) );
  MUX2_X1 U26 ( .A(rf_dout1_e[16]), .B(pc_pls_4_e[16]), .S(n39), .Z(
        alu_a_e[16]) );
  BUF_X1 U27 ( .A(n72), .Z(n39) );
  CLKBUF_X3 U28 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net25305) );
  CLKBUF_X1 U29 ( .A(net25305), .Z(net35228) );
  BUF_X1 U30 ( .A(net32890), .Z(net34366) );
  BUF_X1 U31 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n82) );
  CLKBUF_X1 U32 ( .A(n86), .Z(n11) );
  BUF_X2 U33 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net32889) );
  OR3_X2 U34 ( .A1(n48), .A2(n47), .A3(n46), .ZN(n12) );
  OR3_X2 U35 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n13) );
  NAND2_X1 U36 ( .A1(dmem_dout_wb[22]), .A2(n84), .ZN(n14) );
  NAND2_X1 U37 ( .A1(alu_out_wb[22]), .A2(n81), .ZN(n15) );
  NAND2_X1 U38 ( .A1(pc_pls_4_wb[22]), .A2(n76), .ZN(n16) );
  NAND2_X1 U39 ( .A1(dmem_dout_wb[2]), .A2(n84), .ZN(n17) );
  NAND2_X1 U40 ( .A1(alu_out_wb[2]), .A2(n79), .ZN(n18) );
  NAND2_X1 U41 ( .A1(n76), .A2(pc_pls_4_wb[2]), .ZN(n19) );
  NAND2_X1 U42 ( .A1(dmem_dout_wb[29]), .A2(n33), .ZN(n20) );
  NAND2_X1 U43 ( .A1(alu_out_wb[29]), .A2(n80), .ZN(n21) );
  NAND2_X1 U44 ( .A1(n76), .A2(pc_pls_4_wb[29]), .ZN(n22) );
  CLKBUF_X1 U45 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n34) );
  BUF_X2 U46 ( .A(n150), .Z(n80) );
  OR3_X2 U47 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n23) );
  OR3_X2 U48 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n24) );
  OR3_X2 U49 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n25) );
  OAI21_X2 U50 ( .B1(n39), .B2(n140), .A(n291), .ZN(alu_a_e[19]) );
  OR3_X2 U51 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n26) );
  MUX2_X1 U52 ( .A(rf_dout2_e[6]), .B(imm_e[6]), .S(net32889), .Z(net17723) );
  CLKBUF_X1 U53 ( .A(net32890), .Z(net35180) );
  BUF_X1 U54 ( .A(n151), .Z(n27) );
  BUF_X1 U55 ( .A(n151), .Z(n77) );
  BUF_X1 U56 ( .A(n2), .Z(n28) );
  BUF_X1 U57 ( .A(n151), .Z(n78) );
  OAI21_X2 U58 ( .B1(n86), .B2(n130), .A(n280), .ZN(alu_a_e[29]) );
  BUF_X1 U59 ( .A(n72), .Z(n71) );
  BUF_X1 U60 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n87) );
  AND2_X1 U61 ( .A1(dmem_dout_wb[1]), .A2(n34), .ZN(n30) );
  AND2_X1 U62 ( .A1(alu_out_wb[1]), .A2(n79), .ZN(n31) );
  AND2_X1 U63 ( .A1(n28), .A2(pc_pls_4_wb[1]), .ZN(n32) );
  MUX2_X1 U64 ( .A(rf_dout1_e[1]), .B(pc_pls_4_e[1]), .S(n87), .Z(alu_a_e[1])
         );
  CLKBUF_X3 U65 ( .A(n72), .Z(n85) );
  OR3_X4 U66 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n35) );
  BUF_X1 U67 ( .A(net35180), .Z(net37560) );
  MUX2_X1 U68 ( .A(rf_dout2_e[1]), .B(imm_e[1]), .S(net34800), .Z(net17718) );
  BUF_X1 U69 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net34800) );
  MUX2_X1 U70 ( .A(rf_dout1_e[12]), .B(pc_pls_4_e[12]), .S(n71), .Z(
        alu_a_e[12]) );
  MUX2_X1 U71 ( .A(rf_dout1_e[17]), .B(pc_pls_4_e[17]), .S(n85), .Z(
        alu_a_e[17]) );
  BUF_X1 U72 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net34337) );
  MUX2_X1 U73 ( .A(rf_dout1_e[15]), .B(pc_pls_4_e[15]), .S(n70), .Z(
        alu_a_e[15]) );
  OR3_X4 U74 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n36) );
  OR2_X1 U75 ( .A1(n86), .A2(n138), .ZN(n37) );
  OR3_X4 U76 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n38) );
  OAI21_X1 U77 ( .B1(n86), .B2(n133), .A(n283), .ZN(alu_a_e[26]) );
  BUF_X1 U78 ( .A(net34800), .Z(net35178) );
  BUF_X1 U79 ( .A(net32890), .Z(net35179) );
  BUF_X1 U80 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net32890) );
  BUF_X1 U81 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n88) );
  INV_X1 U82 ( .A(n172), .ZN(n208) );
  AND2_X1 U83 ( .A1(dmem_dout_wb[18]), .A2(n34), .ZN(n40) );
  AND2_X1 U84 ( .A1(alu_out_wb[18]), .A2(n81), .ZN(n41) );
  AND2_X1 U85 ( .A1(n27), .A2(pc_pls_4_wb[18]), .ZN(n42) );
  AND2_X1 U86 ( .A1(dmem_dout_wb[17]), .A2(n33), .ZN(n43) );
  AND2_X1 U87 ( .A1(alu_out_wb[17]), .A2(n80), .ZN(n44) );
  AND2_X1 U88 ( .A1(n1), .A2(pc_pls_4_wb[17]), .ZN(n45) );
  AND2_X1 U89 ( .A1(dmem_dout_wb[16]), .A2(n34), .ZN(n46) );
  AND2_X1 U90 ( .A1(alu_out_wb[16]), .A2(n79), .ZN(n47) );
  AND2_X1 U91 ( .A1(n27), .A2(pc_pls_4_wb[16]), .ZN(n48) );
  AND2_X1 U92 ( .A1(dmem_dout_wb[15]), .A2(n33), .ZN(n49) );
  AND2_X1 U93 ( .A1(alu_out_wb[15]), .A2(n79), .ZN(n50) );
  AND2_X1 U94 ( .A1(n27), .A2(pc_pls_4_wb[15]), .ZN(n51) );
  INV_X1 U95 ( .A(n152), .ZN(n210) );
  INV_X1 U96 ( .A(n153), .ZN(n211) );
  INV_X1 U97 ( .A(n155), .ZN(n213) );
  INV_X1 U98 ( .A(n157), .ZN(n215) );
  INV_X1 U99 ( .A(n159), .ZN(n199) );
  INV_X1 U100 ( .A(n162), .ZN(n200) );
  INV_X1 U101 ( .A(n164), .ZN(n202) );
  INV_X1 U102 ( .A(n166), .ZN(n204) );
  INV_X1 U103 ( .A(n170), .ZN(n207) );
  AND2_X1 U104 ( .A1(dmem_dout_wb[14]), .A2(n34), .ZN(n52) );
  AND2_X1 U105 ( .A1(alu_out_wb[14]), .A2(n80), .ZN(n53) );
  AND2_X1 U106 ( .A1(n27), .A2(pc_pls_4_wb[14]), .ZN(n54) );
  OAI21_X1 U107 ( .B1(n11), .B2(n137), .A(n287), .ZN(alu_a_e[22]) );
  AND2_X1 U108 ( .A1(dmem_dout_wb[13]), .A2(n33), .ZN(n55) );
  AND2_X1 U109 ( .A1(alu_out_wb[13]), .A2(n80), .ZN(n56) );
  AND2_X1 U110 ( .A1(n27), .A2(pc_pls_4_wb[13]), .ZN(n57) );
  AND2_X1 U111 ( .A1(dmem_dout_wb[12]), .A2(n84), .ZN(n58) );
  AND2_X1 U112 ( .A1(alu_out_wb[12]), .A2(n81), .ZN(n59) );
  AND2_X1 U113 ( .A1(n78), .A2(pc_pls_4_wb[12]), .ZN(n60) );
  INV_X1 U114 ( .A(n158), .ZN(n198) );
  INV_X1 U115 ( .A(n149), .ZN(n209) );
  INV_X1 U116 ( .A(n154), .ZN(n212) );
  INV_X1 U117 ( .A(n156), .ZN(n214) );
  AND2_X1 U118 ( .A1(dmem_dout_wb[11]), .A2(n83), .ZN(n61) );
  AND2_X1 U119 ( .A1(alu_out_wb[11]), .A2(n79), .ZN(n62) );
  AND2_X1 U120 ( .A1(n29), .A2(pc_pls_4_wb[11]), .ZN(n63) );
  INV_X1 U121 ( .A(n163), .ZN(n201) );
  INV_X1 U122 ( .A(n165), .ZN(n203) );
  INV_X1 U123 ( .A(n167), .ZN(n205) );
  INV_X1 U124 ( .A(n169), .ZN(n206) );
  OAI21_X1 U125 ( .B1(n86), .B2(n135), .A(n285), .ZN(alu_a_e[24]) );
  AND2_X1 U126 ( .A1(dmem_dout_wb[10]), .A2(n84), .ZN(n64) );
  AND2_X1 U127 ( .A1(alu_out_wb[10]), .A2(n79), .ZN(n65) );
  AND2_X1 U128 ( .A1(n28), .A2(pc_pls_4_wb[10]), .ZN(n66) );
  AND2_X1 U129 ( .A1(dmem_dout_wb[0]), .A2(n83), .ZN(n67) );
  AND2_X1 U130 ( .A1(alu_out_wb[0]), .A2(n80), .ZN(n68) );
  AND2_X1 U131 ( .A1(n77), .A2(pc_pls_4_wb[0]), .ZN(n69) );
  OAI21_X1 U132 ( .B1(n86), .B2(n129), .A(n278), .ZN(alu_a_e[30]) );
  OAI21_X1 U133 ( .B1(n86), .B2(n131), .A(n281), .ZN(alu_a_e[28]) );
  OAI21_X1 U134 ( .B1(n86), .B2(n139), .A(n289), .ZN(alu_a_e[20]) );
  BUF_X2 U135 ( .A(n150), .Z(n79) );
  CLKBUF_X1 U136 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n83) );
  MUX2_X1 U137 ( .A(rf_dout2_e[3]), .B(imm_e[3]), .S(net34337), .Z(n194) );
  MUX2_X1 U138 ( .A(rf_dout1_e[9]), .B(pc_pls_4_e[9]), .S(n70), .Z(alu_a_e[9])
         );
  MUX2_X1 U139 ( .A(rf_dout1_e[7]), .B(pc_pls_4_e[7]), .S(n88), .Z(alu_a_e[7])
         );
  MUX2_X1 U140 ( .A(rf_dout1_e[8]), .B(pc_pls_4_e[8]), .S(n87), .Z(alu_a_e[8])
         );
  BUF_X1 U141 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n70) );
  BUF_X1 U142 ( .A(n92), .Z(n73) );
  BUF_X1 U143 ( .A(n92), .Z(n74) );
  BUF_X1 U144 ( .A(n92), .Z(n75) );
  INV_X1 U145 ( .A(rf_dout1_e[31]), .ZN(n128) );
  NAND2_X1 U146 ( .A1(pc_pls_4_e[31]), .A2(n85), .ZN(n277) );
  INV_X1 U147 ( .A(rf_dout1_e[26]), .ZN(n133) );
  NAND2_X1 U148 ( .A1(pc_pls_4_e[26]), .A2(n85), .ZN(n283) );
  INV_X1 U149 ( .A(rf_dout1_e[25]), .ZN(n134) );
  NAND2_X1 U150 ( .A1(pc_pls_4_e[25]), .A2(n85), .ZN(n284) );
  INV_X1 U151 ( .A(rf_dout1_e[27]), .ZN(n132) );
  NAND2_X1 U152 ( .A1(pc_pls_4_e[27]), .A2(n85), .ZN(n282) );
  INV_X1 U153 ( .A(rf_dout1_e[19]), .ZN(n140) );
  NAND2_X1 U154 ( .A1(pc_pls_4_e[19]), .A2(n85), .ZN(n291) );
  INV_X1 U155 ( .A(rf_dout1_e[24]), .ZN(n135) );
  NAND2_X1 U156 ( .A1(pc_pls_4_e[24]), .A2(n85), .ZN(n285) );
  INV_X1 U157 ( .A(rf_dout1_e[20]), .ZN(n139) );
  NAND2_X1 U158 ( .A1(pc_pls_4_e[20]), .A2(n85), .ZN(n289) );
  INV_X1 U159 ( .A(rf_dout1_e[22]), .ZN(n137) );
  NAND2_X1 U160 ( .A1(pc_pls_4_e[22]), .A2(n85), .ZN(n287) );
  INV_X1 U161 ( .A(rf_dout1_e[21]), .ZN(n138) );
  NAND2_X1 U162 ( .A1(pc_pls_4_e[21]), .A2(n86), .ZN(n288) );
  INV_X1 U163 ( .A(rf_dout1_e[23]), .ZN(n136) );
  NAND2_X1 U164 ( .A1(pc_pls_4_e[23]), .A2(n85), .ZN(n286) );
  INV_X1 U165 ( .A(rf_dout1_e[30]), .ZN(n129) );
  NAND2_X1 U166 ( .A1(pc_pls_4_e[30]), .A2(n85), .ZN(n278) );
  INV_X1 U167 ( .A(rf_dout1_e[29]), .ZN(n130) );
  NAND2_X1 U168 ( .A1(pc_pls_4_e[29]), .A2(n85), .ZN(n280) );
  AOI222_X1 U169 ( .A1(dmem_dout_wb[8]), .A2(n34), .B1(alu_out_wb[8]), .B2(n80), .C1(n77), .C2(pc_pls_4_wb[8]), .ZN(n152) );
  AOI222_X1 U170 ( .A1(dmem_dout_wb[9]), .A2(n33), .B1(alu_out_wb[9]), .B2(n81), .C1(n1), .C2(pc_pls_4_wb[9]), .ZN(n149) );
  AOI222_X1 U171 ( .A1(dmem_dout_wb[19]), .A2(n33), .B1(alu_out_wb[19]), .B2(
        n81), .C1(n29), .C2(pc_pls_4_wb[19]), .ZN(n172) );
  AOI222_X1 U172 ( .A1(dmem_dout_wb[20]), .A2(n83), .B1(alu_out_wb[20]), .B2(
        n81), .C1(n1), .C2(pc_pls_4_wb[20]), .ZN(n170) );
  AOI222_X1 U173 ( .A1(dmem_dout_wb[21]), .A2(n33), .B1(alu_out_wb[21]), .B2(
        n79), .C1(n29), .C2(pc_pls_4_wb[21]), .ZN(n169) );
  AOI222_X1 U175 ( .A1(dmem_dout_wb[23]), .A2(n83), .B1(alu_out_wb[23]), .B2(
        n80), .C1(n77), .C2(pc_pls_4_wb[23]), .ZN(n167) );
  AOI222_X1 U176 ( .A1(dmem_dout_wb[24]), .A2(n83), .B1(alu_out_wb[24]), .B2(
        n80), .C1(n29), .C2(pc_pls_4_wb[24]), .ZN(n166) );
  AOI222_X1 U177 ( .A1(dmem_dout_wb[25]), .A2(n34), .B1(alu_out_wb[25]), .B2(
        n81), .C1(n1), .C2(pc_pls_4_wb[25]), .ZN(n165) );
  AOI222_X1 U178 ( .A1(dmem_dout_wb[26]), .A2(n33), .B1(alu_out_wb[26]), .B2(
        n79), .C1(n78), .C2(pc_pls_4_wb[26]), .ZN(n164) );
  AOI222_X1 U179 ( .A1(dmem_dout_wb[27]), .A2(n84), .B1(alu_out_wb[27]), .B2(
        n79), .C1(n78), .C2(pc_pls_4_wb[27]), .ZN(n163) );
  AOI222_X1 U180 ( .A1(dmem_dout_wb[28]), .A2(n34), .B1(alu_out_wb[28]), .B2(
        n81), .C1(n78), .C2(pc_pls_4_wb[28]), .ZN(n162) );
  AOI222_X1 U181 ( .A1(dmem_dout_wb[30]), .A2(n34), .B1(alu_out_wb[30]), .B2(
        n80), .C1(n28), .C2(pc_pls_4_wb[30]), .ZN(n159) );
  AOI222_X1 U183 ( .A1(dmem_dout_wb[3]), .A2(n84), .B1(alu_out_wb[3]), .B2(n80), .C1(n28), .C2(pc_pls_4_wb[3]), .ZN(n157) );
  AOI222_X1 U184 ( .A1(dmem_dout_wb[4]), .A2(n34), .B1(alu_out_wb[4]), .B2(n79), .C1(n76), .C2(pc_pls_4_wb[4]), .ZN(n156) );
  AOI222_X1 U185 ( .A1(dmem_dout_wb[5]), .A2(n33), .B1(alu_out_wb[5]), .B2(n79), .C1(n29), .C2(pc_pls_4_wb[5]), .ZN(n155) );
  AOI222_X1 U186 ( .A1(dmem_dout_wb[6]), .A2(n83), .B1(alu_out_wb[6]), .B2(n81), .C1(n76), .C2(pc_pls_4_wb[6]), .ZN(n154) );
  AOI222_X1 U187 ( .A1(dmem_dout_wb[7]), .A2(n34), .B1(alu_out_wb[7]), .B2(n81), .C1(n28), .C2(pc_pls_4_wb[7]), .ZN(n153) );
  AOI222_X1 U188 ( .A1(dmem_dout_wb[31]), .A2(n33), .B1(alu_out_wb[31]), .B2(
        n80), .C1(n77), .C2(pc_pls_4_wb[31]), .ZN(n158) );
  NOR4_X1 U189 ( .A1(rf_dout1_e[23]), .A2(rf_dout1_e[22]), .A3(rf_dout1_e[21]), 
        .A4(rf_dout1_e[20]), .ZN(n222) );
  NOR4_X1 U190 ( .A1(rf_dout1_e[5]), .A2(rf_dout1_e[4]), .A3(rf_dout1_e[3]), 
        .A4(rf_dout1_e[31]), .ZN(n225) );
  NAND2_X1 U191 ( .A1(n227), .A2(n228), .ZN(imm_d[31]) );
  NAND2_X1 U192 ( .A1(instr_d[25]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n228) );
  INV_X1 U193 ( .A(\CTRL_WORD[R_TYPE_SEL] ), .ZN(n238) );
  NAND2_X1 U194 ( .A1(n227), .A2(n231), .ZN(imm_d[22]) );
  NAND2_X1 U195 ( .A1(instr_d[22]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n231) );
  NAND2_X1 U196 ( .A1(n227), .A2(n230), .ZN(imm_d[23]) );
  NAND2_X1 U197 ( .A1(instr_d[23]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n230) );
  NAND2_X1 U198 ( .A1(n227), .A2(n229), .ZN(imm_d[24]) );
  NAND2_X1 U199 ( .A1(instr_d[24]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n229) );
  NAND2_X1 U200 ( .A1(n227), .A2(n237), .ZN(imm_d[16]) );
  NAND2_X1 U201 ( .A1(instr_d[16]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n237) );
  NAND2_X1 U202 ( .A1(n227), .A2(n236), .ZN(imm_d[17]) );
  NAND2_X1 U203 ( .A1(instr_d[17]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n236) );
  NAND2_X1 U204 ( .A1(n227), .A2(n235), .ZN(imm_d[18]) );
  NAND2_X1 U205 ( .A1(instr_d[18]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n235) );
  NAND2_X1 U206 ( .A1(n227), .A2(n234), .ZN(imm_d[19]) );
  NAND2_X1 U207 ( .A1(instr_d[19]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n234) );
  NAND2_X1 U208 ( .A1(n227), .A2(n233), .ZN(imm_d[20]) );
  NAND2_X1 U209 ( .A1(instr_d[20]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n233) );
  NAND2_X1 U210 ( .A1(n227), .A2(n232), .ZN(imm_d[21]) );
  NAND2_X1 U211 ( .A1(instr_d[21]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n232) );
  NOR2_X1 U212 ( .A1(n82), .A2(\CTRL_WORD[JAL_EN] ), .ZN(n150) );
  NAND4_X1 U213 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(n218) );
  NOR4_X1 U214 ( .A1(rf_dout1_e[12]), .A2(rf_dout1_e[11]), .A3(rf_dout1_e[10]), 
        .A4(rf_dout1_e[0]), .ZN(n219) );
  NOR4_X1 U215 ( .A1(rf_dout1_e[16]), .A2(rf_dout1_e[15]), .A3(rf_dout1_e[14]), 
        .A4(rf_dout1_e[13]), .ZN(n220) );
  NOR4_X1 U216 ( .A1(rf_dout1_e[1]), .A2(rf_dout1_e[19]), .A3(rf_dout1_e[18]), 
        .A4(rf_dout1_e[17]), .ZN(n221) );
  NAND4_X1 U217 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(n217) );
  NOR4_X1 U218 ( .A1(rf_dout1_e[27]), .A2(rf_dout1_e[26]), .A3(rf_dout1_e[25]), 
        .A4(rf_dout1_e[24]), .ZN(n223) );
  NOR4_X1 U219 ( .A1(rf_dout1_e[30]), .A2(rf_dout1_e[2]), .A3(rf_dout1_e[29]), 
        .A4(rf_dout1_e[28]), .ZN(n224) );
  NOR4_X1 U220 ( .A1(rf_dout1_e[9]), .A2(rf_dout1_e[8]), .A3(rf_dout1_e[7]), 
        .A4(rf_dout1_e[6]), .ZN(n226) );
  NAND2_X1 U221 ( .A1(instr_d[15]), .A2(n216), .ZN(n227) );
  INV_X1 U222 ( .A(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n216) );
  NOR2_X1 U223 ( .A1(n239), .A2(n82), .ZN(n151) );
  INV_X1 U224 ( .A(\CTRL_WORD[JAL_EN] ), .ZN(n239) );
  OR2_X1 U225 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[4]), .ZN(
        rf_waddr_d[4]) );
  OR2_X1 U226 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[3]), .ZN(
        rf_waddr_d[3]) );
  NOR2_X1 U227 ( .A1(n217), .A2(n218), .ZN(n302) );
  INV_X1 U228 ( .A(rf_dout1_e[28]), .ZN(n131) );
  NAND2_X1 U229 ( .A1(pc_pls_4_e[28]), .A2(n85), .ZN(n281) );
  AND2_X1 U230 ( .A1(DMEM_RWADDR[31]), .A2(n184), .ZN(\npc_f[31] ) );
  INV_X1 U231 ( .A(n148), .ZN(n127) );
  AOI22_X1 U232 ( .A1(rs2_e[0]), .A2(n238), .B1(rs3_e[0]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n148) );
  INV_X1 U233 ( .A(n147), .ZN(n126) );
  AOI22_X1 U234 ( .A1(rs2_e[1]), .A2(n238), .B1(rs3_e[1]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n147) );
  INV_X1 U235 ( .A(n146), .ZN(n125) );
  AOI22_X1 U236 ( .A1(rs2_e[2]), .A2(n238), .B1(rs3_e[2]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n146) );
  INV_X1 U237 ( .A(n145), .ZN(n124) );
  AOI22_X1 U238 ( .A1(rs2_e[3]), .A2(n238), .B1(rs3_e[3]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n145) );
  INV_X1 U239 ( .A(n144), .ZN(n123) );
  AOI22_X1 U240 ( .A1(rs2_e[4]), .A2(n238), .B1(rs3_e[4]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n144) );
  BUF_X2 U241 ( .A(RST_AN), .Z(n89) );
  BUF_X2 U242 ( .A(RST_AN), .Z(n90) );
  MUX2_X1 U243 ( .A(rf_dout1_e[2]), .B(pc_pls_4_e[2]), .S(n88), .Z(alu_a_e[2])
         );
  MUX2_X1 U244 ( .A(rf_dout1_e[4]), .B(pc_pls_4_e[4]), .S(n87), .Z(alu_a_e[4])
         );
  MUX2_X1 U245 ( .A(rf_dout2_e[0]), .B(imm_e[0]), .S(\CTRL_WORD[IMM_SEL] ), 
        .Z(n196) );
  MUX2_X1 U246 ( .A(rf_dout2_e[2]), .B(imm_e[2]), .S(net34337), .Z(n195) );
  MUX2_X1 U247 ( .A(rf_dout2_e[4]), .B(imm_e[4]), .S(net32889), .Z(n193) );
  MUX2_X1 U248 ( .A(rf_dout2_e[5]), .B(imm_e[5]), .S(net32889), .Z(n192) );
  MUX2_X1 U249 ( .A(rf_dout2_e[7]), .B(imm_e[7]), .S(net32889), .Z(n191) );
  MUX2_X1 U250 ( .A(rf_dout2_e[8]), .B(imm_e[8]), .S(net32889), .Z(n190) );
  MUX2_X1 U251 ( .A(rf_dout2_e[9]), .B(imm_e[9]), .S(net35178), .Z(n189) );
  MUX2_X1 U252 ( .A(rf_dout2_e[10]), .B(imm_e[10]), .S(net35178), .Z(n188) );
  MUX2_X1 U253 ( .A(rf_dout2_e[11]), .B(imm_e[11]), .S(net25305), .Z(n187) );
  MUX2_X1 U254 ( .A(rf_dout2_e[12]), .B(imm_e[12]), .S(net35179), .Z(n186) );
  MUX2_X1 U255 ( .A(rf_dout2_e[13]), .B(imm_e[13]), .S(net34366), .Z(n185) );
  MUX2_X1 U256 ( .A(rf_dout2_e[14]), .B(imm_e[14]), .S(net35180), .Z(n183) );
  MUX2_X1 U257 ( .A(rf_dout2_e[15]), .B(imm_e[15]), .S(net35179), .Z(n182) );
  MUX2_X1 U258 ( .A(rf_dout2_e[16]), .B(imm_e[16]), .S(net25305), .Z(n181) );
  MUX2_X1 U259 ( .A(rf_dout2_e[17]), .B(imm_e[17]), .S(net37560), .Z(n180) );
  MUX2_X1 U260 ( .A(rf_dout2_e[18]), .B(imm_e[18]), .S(net35228), .Z(n179) );
  MUX2_X1 U261 ( .A(rf_dout2_e[19]), .B(imm_e[19]), .S(net25305), .Z(n178) );
  MUX2_X1 U262 ( .A(rf_dout2_e[20]), .B(imm_e[20]), .S(net25305), .Z(n177) );
  MUX2_X1 U263 ( .A(rf_dout2_e[21]), .B(imm_e[21]), .S(net25305), .Z(n176) );
  MUX2_X1 U264 ( .A(rf_dout2_e[22]), .B(imm_e[22]), .S(net34366), .Z(n175) );
  MUX2_X1 U265 ( .A(rf_dout2_e[23]), .B(imm_e[23]), .S(net25305), .Z(n174) );
  MUX2_X1 U266 ( .A(rf_dout2_e[24]), .B(imm_e[24]), .S(net25305), .Z(n173) );
  MUX2_X1 U267 ( .A(rf_dout2_e[25]), .B(imm_e[25]), .S(net25305), .Z(n171) );
  MUX2_X1 U268 ( .A(rf_dout2_e[26]), .B(imm_e[26]), .S(net37560), .Z(n168) );
  MUX2_X1 U269 ( .A(rf_dout2_e[27]), .B(imm_e[27]), .S(net25305), .Z(n161) );
  MUX2_X1 U270 ( .A(rf_dout2_e[28]), .B(imm_e[28]), .S(net35180), .Z(n160) );
  MUX2_X1 U271 ( .A(rf_dout2_e[29]), .B(imm_e[29]), .S(net25305), .Z(n143) );
  MUX2_X1 U272 ( .A(rf_dout2_e[30]), .B(imm_e[30]), .S(net34366), .Z(n142) );
  MUX2_X1 U273 ( .A(rf_dout2_e[31]), .B(imm_e[31]), .S(net35228), .Z(n141) );
  MUX2_X1 U274 ( .A(rf_dout1_e[0]), .B(pc_pls_4_e[0]), .S(n87), .Z(alu_a_e[0])
         );
  MUX2_X1 U275 ( .A(rf_dout1_e[3]), .B(pc_pls_4_e[3]), .S(n88), .Z(alu_a_e[3])
         );
  MUX2_X1 U276 ( .A(rf_dout1_e[5]), .B(pc_pls_4_e[5]), .S(n71), .Z(alu_a_e[5])
         );
  MUX2_X1 U277 ( .A(rf_dout1_e[6]), .B(pc_pls_4_e[6]), .S(n87), .Z(alu_a_e[6])
         );
  MUX2_X1 U278 ( .A(rf_dout1_e[10]), .B(pc_pls_4_e[10]), .S(n70), .Z(
        alu_a_e[10]) );
  MUX2_X1 U279 ( .A(rf_dout1_e[11]), .B(pc_pls_4_e[11]), .S(n70), .Z(
        alu_a_e[11]) );
  MUX2_X1 U280 ( .A(rf_dout1_e[13]), .B(pc_pls_4_e[13]), .S(n70), .Z(
        alu_a_e[13]) );
  MUX2_X1 U281 ( .A(rf_dout1_e[14]), .B(pc_pls_4_e[14]), .S(n39), .Z(
        alu_a_e[14]) );
  MUX2_X1 U282 ( .A(rf_dout1_e[18]), .B(pc_pls_4_e[18]), .S(n70), .Z(
        alu_a_e[18]) );
  XOR2_X1 U283 ( .A(\DP_SIG[CMPR_0_IS_0_M] ), .B(\CTRL_WORD[COMP_0_INVERT] ), 
        .Z(n91) );
  MUX2_X1 U284 ( .A(\CTRL_WORD[JUMP_EN] ), .B(n91), .S(\CTRL_WORD[BRANCH_EN] ), 
        .Z(n184) );
  INV_X1 U285 ( .A(n184), .ZN(n92) );
  MUX2_X1 U286 ( .A(DMEM_RWADDR[0]), .B(pc_pls_4_f[0]), .S(n73), .Z(n197) );
  MUX2_X1 U287 ( .A(DMEM_RWADDR[1]), .B(pc_pls_4_f[1]), .S(n73), .Z(n122) );
  MUX2_X1 U288 ( .A(DMEM_RWADDR[2]), .B(pc_pls_4_f[2]), .S(n73), .Z(n121) );
  MUX2_X1 U289 ( .A(DMEM_RWADDR[3]), .B(pc_pls_4_f[3]), .S(n73), .Z(n120) );
  MUX2_X1 U290 ( .A(DMEM_RWADDR[4]), .B(pc_pls_4_f[4]), .S(n73), .Z(n119) );
  MUX2_X1 U291 ( .A(DMEM_RWADDR[5]), .B(pc_pls_4_f[5]), .S(n73), .Z(n118) );
  MUX2_X1 U292 ( .A(DMEM_RWADDR[6]), .B(pc_pls_4_f[6]), .S(n73), .Z(n117) );
  MUX2_X1 U293 ( .A(DMEM_RWADDR[7]), .B(pc_pls_4_f[7]), .S(n73), .Z(n116) );
  MUX2_X1 U294 ( .A(DMEM_RWADDR[8]), .B(pc_pls_4_f[8]), .S(n73), .Z(n115) );
  MUX2_X1 U295 ( .A(DMEM_RWADDR[9]), .B(pc_pls_4_f[9]), .S(n73), .Z(n114) );
  MUX2_X1 U296 ( .A(DMEM_RWADDR[10]), .B(pc_pls_4_f[10]), .S(n73), .Z(n113) );
  MUX2_X1 U297 ( .A(DMEM_RWADDR[11]), .B(pc_pls_4_f[11]), .S(n74), .Z(n112) );
  MUX2_X1 U298 ( .A(DMEM_RWADDR[12]), .B(pc_pls_4_f[12]), .S(n74), .Z(n111) );
  MUX2_X1 U299 ( .A(DMEM_RWADDR[13]), .B(pc_pls_4_f[13]), .S(n74), .Z(n110) );
  MUX2_X1 U300 ( .A(DMEM_RWADDR[14]), .B(pc_pls_4_f[14]), .S(n74), .Z(n109) );
  MUX2_X1 U301 ( .A(DMEM_RWADDR[15]), .B(pc_pls_4_f[15]), .S(n74), .Z(n108) );
  MUX2_X1 U302 ( .A(DMEM_RWADDR[16]), .B(pc_pls_4_f[16]), .S(n74), .Z(n107) );
  MUX2_X1 U303 ( .A(DMEM_RWADDR[17]), .B(pc_pls_4_f[17]), .S(n74), .Z(n106) );
  MUX2_X1 U304 ( .A(DMEM_RWADDR[18]), .B(pc_pls_4_f[18]), .S(n74), .Z(n105) );
  MUX2_X1 U305 ( .A(DMEM_RWADDR[19]), .B(pc_pls_4_f[19]), .S(n74), .Z(n104) );
  MUX2_X1 U306 ( .A(DMEM_RWADDR[20]), .B(pc_pls_4_f[20]), .S(n74), .Z(n103) );
  MUX2_X1 U307 ( .A(DMEM_RWADDR[21]), .B(pc_pls_4_f[21]), .S(n74), .Z(n102) );
  MUX2_X1 U308 ( .A(DMEM_RWADDR[22]), .B(pc_pls_4_f[22]), .S(n75), .Z(n101) );
  MUX2_X1 U309 ( .A(DMEM_RWADDR[23]), .B(pc_pls_4_f[23]), .S(n75), .Z(n100) );
  MUX2_X1 U310 ( .A(DMEM_RWADDR[24]), .B(pc_pls_4_f[24]), .S(n75), .Z(n99) );
  MUX2_X1 U311 ( .A(DMEM_RWADDR[25]), .B(pc_pls_4_f[25]), .S(n75), .Z(n98) );
  MUX2_X1 U312 ( .A(DMEM_RWADDR[26]), .B(pc_pls_4_f[26]), .S(n75), .Z(n97) );
  MUX2_X1 U313 ( .A(DMEM_RWADDR[27]), .B(pc_pls_4_f[27]), .S(n75), .Z(n96) );
  MUX2_X1 U314 ( .A(DMEM_RWADDR[28]), .B(pc_pls_4_f[28]), .S(n75), .Z(n95) );
  MUX2_X1 U315 ( .A(DMEM_RWADDR[29]), .B(pc_pls_4_f[29]), .S(n75), .Z(n94) );
  MUX2_X1 U316 ( .A(DMEM_RWADDR[30]), .B(pc_pls_4_f[30]), .S(n75), .Z(n93) );
endmodule


module HU ( CLK, RST_AN, .DP_SIG({\DP_SIG[CMPR_0_IS_0_M] , 
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }), 
    .HZRD_SIG({\HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , 
        \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , 
        \HZRD_SIG[FLUSH_MWB] }) );
  input CLK, RST_AN, \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  output \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] ,
         \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] ;
  wire   n2, n3, n4, n1, \HZRD_SIG[FLUSH_FD] , n6;
  assign \HZRD_SIG[FLUSH_MWB]  = 1'b0;
  assign \HZRD_SIG[STALL_DE]  = 1'b0;
  assign \HZRD_SIG[STALL_FD]  = 1'b0;
  assign \HZRD_SIG[FLUSH_DE]  = \HZRD_SIG[FLUSH_FD] ;
  assign \HZRD_SIG[FLUSH_EM]  = \HZRD_SIG[FLUSH_FD] ;

  OR4_X1 U3 ( .A1(\DP_SIG[INSTR_OPCODE_M][3] ), .A2(n2), .A3(
        \DP_SIG[INSTR_OPCODE_M][5] ), .A4(\DP_SIG[INSTR_OPCODE_M][4] ), .ZN(n1) );
  INV_X2 U4 ( .A(n1), .ZN(\HZRD_SIG[FLUSH_FD] ) );
  AOI22_X1 U5 ( .A1(n3), .A2(\DP_SIG[INSTR_OPCODE_M][2] ), .B1(
        \DP_SIG[INSTR_OPCODE_M][1] ), .B2(n6), .ZN(n2) );
  INV_X1 U6 ( .A(\DP_SIG[INSTR_OPCODE_M][2] ), .ZN(n6) );
  NOR2_X1 U7 ( .A1(\DP_SIG[INSTR_OPCODE_M][1] ), .A2(n4), .ZN(n3) );
  XNOR2_X1 U8 ( .A(\DP_SIG[INSTR_OPCODE_M][0] ), .B(\DP_SIG[CMPR_0_IS_0_M] ), 
        .ZN(n4) );
endmodule


module CPU ( CLK, RST_AN, IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, DMEM_WEN, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN;
  output DMEM_WEN;
  wire   \hzrd_sig[FLUSH_FD] , \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] ,
         \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] ,
         \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] ,
         \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] ,
         \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] ,
         \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] ,
         \ctrl_word[COMP_0_INVERT] , \ctrl_word[RF_WB_DMEM_DOUT_SEL] ,
         \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] , \dp_sig[CMPR_0_IS_0_M] ,
         \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] ,
         \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] ,
         \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] ;
  wire   [31:0] instr_cu;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  CU U_CU ( .CLK(CLK), .RST_AN(RST_AN), .INSTR(instr_cu), .HZRD_SIG({1'b0, 
        \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        1'b0}), .CTRL_WORD({\ctrl_word[J_TYPE_IMM_SEL] , 
        \ctrl_word[R_TYPE_SEL] , \ctrl_word[IMM_SEL] , 
        \ctrl_word[PC_PLS_4_SEL] , \ctrl_word[ALU_FUNC][3] , 
        \ctrl_word[ALU_FUNC][2] , \ctrl_word[ALU_FUNC][1] , 
        \ctrl_word[ALU_FUNC][0] , \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }) );
  DATAPATH U_DATAPATH ( .CLK(CLK), .RST_AN(RST_AN), .CTRL_WORD({
        \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] , 
        \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] , 
        \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] , 
        \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] , 
        \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }), .INSTR_CU(instr_cu), 
        .HZRD_SIG({1'b0, \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , 
        \hzrd_sig[FLUSH_EM] , 1'b0}), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), 
        .IMEM_ADDR(IMEM_ADDR), .IMEM_DOUT(IMEM_DOUT), .DMEM_RWADDR(DMEM_RWADDR), .DMEM_DIN(DMEM_DIN), .DMEM_DOUT(DMEM_DOUT) );
  HU U_HU ( .CLK(CLK), .RST_AN(RST_AN), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), .HZRD_SIG(
        {SYNOPSYS_UNCONNECTED__0, \hzrd_sig[FLUSH_FD] , 
        SYNOPSYS_UNCONNECTED__1, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        SYNOPSYS_UNCONNECTED__2}) );
endmodule

