
module CU ( CLK, RST_AN, INSTR, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .CTRL_WORD({
        \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] , 
        \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] , 
        \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] , 
        \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] , 
        \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }) );
  input [31:0] INSTR;
  input CLK, RST_AN, \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] ;
  wire   INSTR_31, INSTR_30, INSTR_29, INSTR_28, INSTR_27, INSTR_26,
         \execute_sig_d1[R_TYPE_SEL] , \execute_sig_d1[IMM_SEL] ,
         \execute_sig_d1[ALU_FUNC][2] , \memory_sig_d1[DMEM_WEN] ,
         \memory_sig_d1[BRANCH_EN] , \memory_sig_d1[JUMP_EN] ,
         \memory_sig_d1[COMP_0_INVERT] ,
         \writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d1[JAL_EN] ,
         \writeback_sig_d1[RF_WEN] , \memory_sig_d2[DMEM_WEN] ,
         \memory_sig_d2[BRANCH_EN] , \memory_sig_d2[JUMP_EN] ,
         \memory_sig_d2[COMP_0_INVERT] ,
         \writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d2[JAL_EN] ,
         \writeback_sig_d2[RF_WEN] , \writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ,
         \writeback_sig_d3[JAL_EN] , N213, N215, N216, N217, N218, N224, N228,
         N229, N231, n1, n26, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178;
  assign INSTR_31 = INSTR[31];
  assign INSTR_30 = INSTR[30];
  assign INSTR_29 = INSTR[29];
  assign INSTR_28 = INSTR[28];
  assign INSTR_27 = INSTR[27];
  assign INSTR_26 = INSTR[26];

  DFFR_X1 \decode_sig_d1_reg[J_TYPE_IMM_SEL]  ( .D(n157), .CK(CLK), .RN(n150), 
        .Q(\CTRL_WORD[J_TYPE_IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[IMM_SEL]  ( .D(N218), .CK(CLK), .RN(n150), .Q(
        \execute_sig_d1[IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[PC_PLS_4_SEL]  ( .D(N217), .CK(CLK), .RN(n150), 
        .QN(n110) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][3]  ( .D(N216), .CK(CLK), .SN(n152), 
        .QN(n113) );
  DFFR_X1 \execute_sig_d1_reg[ALU_FUNC][2]  ( .D(N215), .CK(CLK), .RN(n150), 
        .Q(\execute_sig_d1[ALU_FUNC][2] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][1]  ( .D(n158), .CK(CLK), .SN(n152), 
        .QN(n112) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][0]  ( .D(N213), .CK(CLK), .SN(n152), 
        .QN(n111) );
  DFFR_X1 \memory_sig_d1_reg[BRANCH_EN]  ( .D(n114), .CK(CLK), .RN(n150), .Q(
        \memory_sig_d1[BRANCH_EN] ) );
  DFFR_X1 \memory_sig_d1_reg[JUMP_EN]  ( .D(n157), .CK(CLK), .RN(n150), .Q(
        \memory_sig_d1[JUMP_EN] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n156), .CK(CLK), 
        .RN(n150), .Q(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WEN]  ( .D(N224), .CK(CLK), .RN(n150), .Q(
        \writeback_sig_d1[RF_WEN] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][3]  ( .D(N231), .CK(CLK), .SN(n153), 
        .Q(\CTRL_WORD[ALU_FUNC][3] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][1]  ( .D(N229), .CK(CLK), .SN(n152), 
        .Q(\CTRL_WORD[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][0]  ( .D(N228), .CK(CLK), .SN(n153), 
        .Q(\CTRL_WORD[ALU_FUNC][0] ) );
  DFFRS_X2 \execute_sig_d2_reg[PC_PLS_4_SEL]  ( .D(n26), .CK(CLK), .RN(n150), 
        .SN(1'b1), .Q(\CTRL_WORD[PC_PLS_4_SEL] ) );
  DFFR_X1 \writeback_sig_d4_reg[RF_WEN]  ( .D(n1), .CK(CLK), .RN(n150), .Q(
        \CTRL_WORD[RF_WEN] ) );
  NAND3_X1 U110 ( .A1(n159), .A2(n169), .A3(n56), .ZN(n55) );
  NAND3_X1 U111 ( .A1(n56), .A2(n159), .A3(INSTR_31), .ZN(n52) );
  NAND3_X1 U112 ( .A1(n168), .A2(INSTR_27), .A3(INSTR_30), .ZN(n65) );
  NAND3_X1 U113 ( .A1(n68), .A2(n159), .A3(INSTR_27), .ZN(n62) );
  NAND3_X1 U114 ( .A1(INSTR_26), .A2(n75), .A3(INSTR_29), .ZN(n74) );
  OAI33_X1 U115 ( .A1(n89), .A2(INSTR_31), .A3(n163), .B1(n81), .B2(INSTR[2]), 
        .B3(n90), .ZN(n87) );
  NAND3_X1 U116 ( .A1(n60), .A2(n76), .A3(n63), .ZN(n91) );
  OAI33_X1 U117 ( .A1(n97), .A2(INSTR[0]), .A3(n98), .B1(n164), .B2(INSTR[5]), 
        .B3(INSTR[1]), .ZN(n96) );
  NAND3_X1 U118 ( .A1(n101), .A2(n102), .A3(INSTR[3]), .ZN(n90) );
  NAND3_X1 U119 ( .A1(n101), .A2(n177), .A3(INSTR[2]), .ZN(n82) );
  NAND3_X1 U120 ( .A1(n173), .A2(n172), .A3(n68), .ZN(n97) );
  DFFRS_X2 \execute_sig_d2_reg[IMM_SEL]  ( .D(n146), .CK(CLK), .RN(n151), .SN(
        1'b1), .Q(\CTRL_WORD[IMM_SEL] ) );
  DFFR_X1 \writeback_sig_d3_reg[RF_WEN]  ( .D(n144), .CK(CLK), .RN(RST_AN), 
        .QN(n109) );
  DFFR_X1 \writeback_sig_d4_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n143), .CK(CLK), 
        .RN(RST_AN), .Q(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d4_reg[JAL_EN]  ( .D(n142), .CK(CLK), .RN(n152), .Q(
        \CTRL_WORD[JAL_EN] ) );
  DFFR_X1 \writeback_sig_d3_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n141), .CK(CLK), 
        .RN(n152), .Q(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d3_reg[JAL_EN]  ( .D(n140), .CK(CLK), .RN(n152), .Q(
        \writeback_sig_d3[JAL_EN] ) );
  DFFR_X1 \memory_sig_d3_reg[JUMP_EN]  ( .D(n139), .CK(CLK), .RN(n152), .Q(
        \CTRL_WORD[JUMP_EN] ) );
  DFFR_X1 \memory_sig_d3_reg[DMEM_WEN]  ( .D(n138), .CK(CLK), .RN(n152), .Q(
        \CTRL_WORD[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d3_reg[COMP_0_INVERT]  ( .D(n137), .CK(CLK), .RN(n152), 
        .Q(\CTRL_WORD[COMP_0_INVERT] ) );
  DFFR_X1 \memory_sig_d3_reg[BRANCH_EN]  ( .D(n136), .CK(CLK), .RN(n151), .Q(
        \CTRL_WORD[BRANCH_EN] ) );
  DFFR_X1 \execute_sig_d1_reg[R_TYPE_SEL]  ( .D(n135), .CK(CLK), .RN(n151), 
        .Q(\execute_sig_d1[R_TYPE_SEL] ) );
  DFFR_X1 \writeback_sig_d2_reg[RF_WEN]  ( .D(n134), .CK(CLK), .RN(n151), .Q(
        \writeback_sig_d2[RF_WEN] ) );
  DFFR_X1 \writeback_sig_d2_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n133), .CK(CLK), 
        .RN(n151), .Q(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d2_reg[JAL_EN]  ( .D(n132), .CK(CLK), .RN(n151), .Q(
        \writeback_sig_d2[JAL_EN] ) );
  DFFR_X1 \memory_sig_d2_reg[JUMP_EN]  ( .D(n131), .CK(CLK), .RN(n151), .Q(
        \memory_sig_d2[JUMP_EN] ) );
  DFFR_X1 \memory_sig_d2_reg[DMEM_WEN]  ( .D(n130), .CK(CLK), .RN(n151), .Q(
        \memory_sig_d2[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d2_reg[COMP_0_INVERT]  ( .D(n129), .CK(CLK), .RN(n151), 
        .Q(\memory_sig_d2[COMP_0_INVERT] ) );
  DFFR_X1 \memory_sig_d2_reg[BRANCH_EN]  ( .D(n128), .CK(CLK), .RN(n151), .Q(
        \memory_sig_d2[BRANCH_EN] ) );
  DFFR_X1 \execute_sig_d2_reg[R_TYPE_SEL]  ( .D(n127), .CK(CLK), .RN(n151), 
        .Q(\CTRL_WORD[R_TYPE_SEL] ) );
  DFFR_X1 \memory_sig_d1_reg[DMEM_WEN]  ( .D(n126), .CK(CLK), .RN(n152), .Q(
        \memory_sig_d1[DMEM_WEN] ) );
  DFFR_X1 \writeback_sig_d1_reg[JAL_EN]  ( .D(n125), .CK(CLK), .RN(n150), .Q(
        \writeback_sig_d1[JAL_EN] ) );
  DFFR_X1 \memory_sig_d1_reg[COMP_0_INVERT]  ( .D(n124), .CK(CLK), .RN(n151), 
        .Q(\memory_sig_d1[COMP_0_INVERT] ) );
  DFFR_X1 \execute_sig_d2_reg[ALU_FUNC][2]  ( .D(n147), .CK(CLK), .RN(RST_AN), 
        .Q(\CTRL_WORD[ALU_FUNC][2] ) );
  AND2_X1 U3 ( .A1(INSTR_26), .A2(n114), .ZN(n124) );
  AND2_X1 U4 ( .A1(INSTR_26), .A2(n157), .ZN(n125) );
  AND2_X1 U5 ( .A1(INSTR_29), .A2(n156), .ZN(n126) );
  AND2_X1 U6 ( .A1(\execute_sig_d1[R_TYPE_SEL] ), .A2(n155), .ZN(n127) );
  AND2_X1 U7 ( .A1(\memory_sig_d1[BRANCH_EN] ), .A2(n155), .ZN(n128) );
  AND2_X1 U8 ( .A1(\memory_sig_d1[COMP_0_INVERT] ), .A2(n155), .ZN(n129) );
  AND2_X1 U9 ( .A1(\memory_sig_d1[DMEM_WEN] ), .A2(n155), .ZN(n130) );
  AND2_X1 U10 ( .A1(\memory_sig_d1[JUMP_EN] ), .A2(n155), .ZN(n131) );
  AND2_X1 U11 ( .A1(\writeback_sig_d1[JAL_EN] ), .A2(n155), .ZN(n132) );
  AND2_X1 U12 ( .A1(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ), .A2(n155), .ZN(
        n133) );
  AND2_X1 U13 ( .A1(\writeback_sig_d1[RF_WEN] ), .A2(n155), .ZN(n134) );
  AND2_X1 U14 ( .A1(n163), .A2(n159), .ZN(n135) );
  AND2_X1 U15 ( .A1(\memory_sig_d2[BRANCH_EN] ), .A2(n154), .ZN(n136) );
  AND2_X1 U16 ( .A1(\memory_sig_d2[COMP_0_INVERT] ), .A2(n154), .ZN(n137) );
  AND2_X1 U17 ( .A1(\memory_sig_d2[DMEM_WEN] ), .A2(n154), .ZN(n138) );
  AND2_X1 U18 ( .A1(\memory_sig_d2[JUMP_EN] ), .A2(n154), .ZN(n139) );
  AND2_X1 U19 ( .A1(\writeback_sig_d2[JAL_EN] ), .A2(n154), .ZN(n140) );
  AND2_X1 U20 ( .A1(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ), .A2(n154), .ZN(
        n141) );
  AND2_X1 U22 ( .A1(\writeback_sig_d3[JAL_EN] ), .A2(n160), .ZN(n142) );
  AND2_X1 U23 ( .A1(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ), .A2(n160), .ZN(
        n143) );
  AND2_X1 U24 ( .A1(\writeback_sig_d2[RF_WEN] ), .A2(n154), .ZN(n144) );
  INV_X1 U25 ( .A(n97), .ZN(n163) );
  INV_X1 U26 ( .A(\HZRD_SIG[FLUSH_DE] ), .ZN(n155) );
  INV_X1 U27 ( .A(\HZRD_SIG[FLUSH_FD] ), .ZN(n159) );
  INV_X1 U28 ( .A(\HZRD_SIG[FLUSH_EM] ), .ZN(n154) );
  OAI221_X1 U29 ( .B1(n82), .B2(n103), .C1(n56), .C2(n161), .A(n159), .ZN(n88)
         );
  NAND2_X1 U30 ( .A1(n162), .A2(n86), .ZN(n103) );
  INV_X1 U31 ( .A(n81), .ZN(n162) );
  NAND2_X1 U32 ( .A1(n159), .A2(n161), .ZN(n54) );
  OAI211_X1 U33 ( .C1(n61), .C2(n54), .A(n62), .B(n52), .ZN(N218) );
  AOI21_X1 U34 ( .B1(n171), .B2(n63), .A(n58), .ZN(n61) );
  INV_X1 U35 ( .A(n62), .ZN(n157) );
  INV_X1 U36 ( .A(n52), .ZN(n156) );
  OR2_X1 U37 ( .A1(n114), .A2(n157), .ZN(N217) );
  BUF_X1 U38 ( .A(n149), .Z(n152) );
  BUF_X1 U39 ( .A(n148), .Z(n150) );
  BUF_X1 U40 ( .A(n148), .Z(n151) );
  OAI21_X1 U41 ( .B1(n67), .B2(n93), .A(n94), .ZN(n92) );
  NAND2_X1 U42 ( .A1(n172), .A2(n170), .ZN(n60) );
  INV_X1 U43 ( .A(n90), .ZN(n174) );
  INV_X1 U44 ( .A(n59), .ZN(n168) );
  AND2_X1 U45 ( .A1(n73), .A2(n166), .ZN(n56) );
  INV_X1 U46 ( .A(n67), .ZN(n171) );
  NAND2_X1 U47 ( .A1(n165), .A2(n173), .ZN(n66) );
  INV_X1 U48 ( .A(n63), .ZN(n167) );
  INV_X1 U49 ( .A(n78), .ZN(n164) );
  INV_X1 U50 ( .A(n93), .ZN(n165) );
  INV_X1 U51 ( .A(n102), .ZN(n175) );
  OR2_X1 U52 ( .A1(n66), .A2(n172), .ZN(n83) );
  BUF_X1 U53 ( .A(n149), .Z(n153) );
  NOR2_X1 U54 ( .A1(\HZRD_SIG[FLUSH_FD] ), .A2(n77), .ZN(N215) );
  AOI221_X1 U55 ( .B1(n78), .B2(n175), .C1(n79), .C2(INSTR_28), .A(n80), .ZN(
        n77) );
  AOI21_X1 U56 ( .B1(n83), .B2(n84), .A(INSTR_31), .ZN(n79) );
  NOR4_X1 U57 ( .A1(INSTR[5]), .A2(n81), .A3(n82), .A4(n178), .ZN(n80) );
  NOR4_X1 U58 ( .A1(n54), .A2(n67), .A3(INSTR_29), .A4(INSTR_30), .ZN(n114) );
  OAI211_X1 U59 ( .C1(n163), .C2(n69), .A(n70), .B(n159), .ZN(N216) );
  OAI211_X1 U60 ( .C1(INSTR[0]), .C2(INSTR[2]), .A(n174), .B(n163), .ZN(n70)
         );
  AOI221_X1 U61 ( .B1(n71), .B2(n169), .C1(n167), .C2(n172), .A(n72), .ZN(n69)
         );
  OAI221_X1 U62 ( .B1(n73), .B2(n161), .C1(n168), .C2(n166), .A(n74), .ZN(n72)
         );
  NAND2_X1 U63 ( .A1(n112), .A2(n155), .ZN(N229) );
  NAND2_X1 U64 ( .A1(n111), .A2(n155), .ZN(N228) );
  NAND2_X1 U65 ( .A1(n113), .A2(n155), .ZN(N231) );
  OAI211_X1 U66 ( .C1(n53), .C2(n54), .A(n55), .B(n52), .ZN(N224) );
  AOI221_X1 U67 ( .B1(n57), .B2(n173), .C1(INSTR_29), .C2(n171), .A(n58), .ZN(
        n53) );
  OAI22_X1 U68 ( .A1(n59), .A2(n166), .B1(INSTR_30), .B2(n60), .ZN(n57) );
  OR3_X1 U69 ( .A1(n95), .A2(n88), .A3(n96), .ZN(N213) );
  NOR3_X1 U70 ( .A1(n105), .A2(INSTR_31), .A3(n163), .ZN(n95) );
  AOI221_X1 U71 ( .B1(INSTR_30), .B2(n106), .C1(n71), .C2(n169), .A(n107), 
        .ZN(n105) );
  INV_X1 U72 ( .A(n85), .ZN(n158) );
  AOI211_X1 U73 ( .C1(n78), .C2(n86), .A(n87), .B(n88), .ZN(n85) );
  AOI221_X1 U74 ( .B1(n91), .B2(n169), .C1(INSTR_30), .C2(n67), .A(n92), .ZN(
        n89) );
  NOR2_X1 U75 ( .A1(\HZRD_SIG[FLUSH_MWB] ), .A2(n109), .ZN(n1) );
  NOR4_X1 U76 ( .A1(INSTR[6]), .A2(INSTR[4]), .A3(INSTR[10]), .A4(n104), .ZN(
        n101) );
  OR3_X1 U77 ( .A1(INSTR[9]), .A2(INSTR[8]), .A3(INSTR[7]), .ZN(n104) );
  NOR3_X1 U78 ( .A1(n97), .A2(INSTR[0]), .A3(n82), .ZN(n78) );
  NOR4_X1 U79 ( .A1(INSTR_28), .A2(INSTR_29), .A3(INSTR_30), .A4(INSTR_31), 
        .ZN(n68) );
  INV_X1 U80 ( .A(INSTR[3]), .ZN(n177) );
  NOR3_X1 U81 ( .A1(n172), .A2(INSTR_28), .A3(n173), .ZN(n73) );
  INV_X1 U82 ( .A(INSTR_27), .ZN(n172) );
  OAI211_X1 U83 ( .C1(n63), .C2(n64), .A(n65), .B(n66), .ZN(n58) );
  NAND2_X1 U84 ( .A1(INSTR_29), .A2(n172), .ZN(n64) );
  OAI22_X1 U85 ( .A1(INSTR_29), .A2(INSTR_27), .B1(INSTR_26), .B2(n168), .ZN(
        n106) );
  OAI21_X1 U86 ( .B1(INSTR[5]), .B2(n178), .A(n175), .ZN(n86) );
  OAI21_X1 U87 ( .B1(INSTR_30), .B2(n76), .A(n60), .ZN(n71) );
  INV_X1 U88 ( .A(INSTR_29), .ZN(n169) );
  NAND2_X1 U89 ( .A1(INSTR_28), .A2(n172), .ZN(n67) );
  INV_X1 U90 ( .A(INSTR_26), .ZN(n173) );
  OAI211_X1 U91 ( .C1(INSTR_27), .C2(n173), .A(n169), .B(INSTR_30), .ZN(n84)
         );
  NOR2_X1 U92 ( .A1(n176), .A2(INSTR[1]), .ZN(n102) );
  NAND2_X1 U93 ( .A1(INSTR_30), .A2(INSTR_26), .ZN(n63) );
  OAI21_X1 U94 ( .B1(n108), .B2(n172), .A(n94), .ZN(n107) );
  AOI21_X1 U95 ( .B1(INSTR_29), .B2(n170), .A(n167), .ZN(n108) );
  INV_X1 U96 ( .A(INSTR_30), .ZN(n166) );
  AOI21_X1 U97 ( .B1(INSTR[2]), .B2(n174), .A(n99), .ZN(n98) );
  NOR4_X1 U98 ( .A1(n100), .A2(n176), .A3(INSTR[3]), .A4(INSTR[2]), .ZN(n99)
         );
  NAND2_X1 U99 ( .A1(INSTR[1]), .A2(n101), .ZN(n100) );
  OAI21_X1 U100 ( .B1(INSTR_31), .B2(INSTR_28), .A(n76), .ZN(n75) );
  NAND2_X1 U101 ( .A1(INSTR[0]), .A2(n163), .ZN(n81) );
  NAND2_X1 U102 ( .A1(INSTR_27), .A2(INSTR_28), .ZN(n76) );
  INV_X1 U103 ( .A(INSTR_31), .ZN(n161) );
  NAND2_X1 U104 ( .A1(INSTR_29), .A2(n166), .ZN(n93) );
  NAND2_X1 U105 ( .A1(INSTR_28), .A2(n169), .ZN(n59) );
  NAND2_X1 U106 ( .A1(n165), .A2(INSTR_26), .ZN(n94) );
  INV_X1 U107 ( .A(INSTR[1]), .ZN(n178) );
  INV_X1 U108 ( .A(INSTR_28), .ZN(n170) );
  INV_X1 U109 ( .A(INSTR[5]), .ZN(n176) );
  BUF_X1 U121 ( .A(RST_AN), .Z(n149) );
  BUF_X1 U122 ( .A(RST_AN), .Z(n148) );
  INV_X1 U123 ( .A(\HZRD_SIG[FLUSH_MWB] ), .ZN(n160) );
  AND2_X1 U125 ( .A1(\execute_sig_d1[IMM_SEL] ), .A2(n155), .ZN(n146) );
  AND2_X1 U126 ( .A1(\execute_sig_d1[ALU_FUNC][2] ), .A2(n155), .ZN(n147) );
  NOR2_X1 U127 ( .A1(n110), .A2(\HZRD_SIG[FLUSH_DE] ), .ZN(n26) );
endmodule


module REG_PIPO_32_fffffffc_fffffffc_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n21, n22, n23;

  DFFS_X1 \reg_mem_reg[31]  ( .D(n96), .CK(CLK), .SN(n23), .Q(DOUT[31]), .QN(
        n64) );
  DFFS_X1 \reg_mem_reg[30]  ( .D(n95), .CK(CLK), .SN(n23), .Q(DOUT[30]) );
  DFFS_X1 \reg_mem_reg[29]  ( .D(n94), .CK(CLK), .SN(n23), .Q(DOUT[29]) );
  DFFS_X1 \reg_mem_reg[28]  ( .D(n93), .CK(CLK), .SN(n23), .Q(DOUT[28]) );
  DFFS_X1 \reg_mem_reg[27]  ( .D(n92), .CK(CLK), .SN(n23), .Q(DOUT[27]) );
  DFFS_X1 \reg_mem_reg[26]  ( .D(n91), .CK(CLK), .SN(n23), .Q(DOUT[26]) );
  DFFS_X1 \reg_mem_reg[25]  ( .D(n90), .CK(CLK), .SN(n22), .Q(DOUT[25]) );
  DFFS_X1 \reg_mem_reg[24]  ( .D(n89), .CK(CLK), .SN(n22), .Q(DOUT[24]) );
  DFFS_X1 \reg_mem_reg[23]  ( .D(n88), .CK(CLK), .SN(n22), .Q(DOUT[23]) );
  DFFS_X1 \reg_mem_reg[22]  ( .D(n87), .CK(CLK), .SN(n22), .Q(DOUT[22]) );
  DFFS_X1 \reg_mem_reg[21]  ( .D(n86), .CK(CLK), .SN(n22), .Q(DOUT[21]) );
  DFFS_X1 \reg_mem_reg[20]  ( .D(n85), .CK(CLK), .SN(n22), .Q(DOUT[20]) );
  DFFS_X1 \reg_mem_reg[19]  ( .D(n84), .CK(CLK), .SN(n22), .Q(DOUT[19]), .QN(
        n52) );
  DFFS_X1 \reg_mem_reg[18]  ( .D(n83), .CK(CLK), .SN(n22), .Q(DOUT[18]), .QN(
        n51) );
  DFFS_X1 \reg_mem_reg[17]  ( .D(n82), .CK(CLK), .SN(n22), .Q(DOUT[17]), .QN(
        n50) );
  DFFS_X1 \reg_mem_reg[16]  ( .D(n81), .CK(CLK), .SN(n22), .Q(DOUT[16]), .QN(
        n49) );
  DFFS_X1 \reg_mem_reg[15]  ( .D(n80), .CK(CLK), .SN(n22), .Q(DOUT[15]), .QN(
        n48) );
  DFFS_X1 \reg_mem_reg[14]  ( .D(n79), .CK(CLK), .SN(n22), .Q(DOUT[14]), .QN(
        n47) );
  DFFS_X1 \reg_mem_reg[13]  ( .D(n78), .CK(CLK), .SN(n22), .Q(DOUT[13]), .QN(
        n46) );
  DFFS_X1 \reg_mem_reg[12]  ( .D(n77), .CK(CLK), .SN(n21), .Q(DOUT[12]), .QN(
        n45) );
  DFFS_X1 \reg_mem_reg[11]  ( .D(n76), .CK(CLK), .SN(n21), .Q(DOUT[11]), .QN(
        n44) );
  DFFS_X1 \reg_mem_reg[10]  ( .D(n75), .CK(CLK), .SN(n21), .Q(DOUT[10]), .QN(
        n43) );
  DFFS_X1 \reg_mem_reg[9]  ( .D(n74), .CK(CLK), .SN(n21), .Q(DOUT[9]), .QN(n42) );
  DFFS_X1 \reg_mem_reg[8]  ( .D(n73), .CK(CLK), .SN(n21), .Q(DOUT[8]), .QN(n41) );
  DFFS_X1 \reg_mem_reg[7]  ( .D(n72), .CK(CLK), .SN(n21), .Q(DOUT[7]), .QN(n40) );
  DFFS_X1 \reg_mem_reg[6]  ( .D(n71), .CK(CLK), .SN(n21), .Q(DOUT[6]), .QN(n39) );
  DFFS_X1 \reg_mem_reg[5]  ( .D(n70), .CK(CLK), .SN(n21), .Q(DOUT[5]), .QN(n38) );
  DFFS_X1 \reg_mem_reg[4]  ( .D(n69), .CK(CLK), .SN(n21), .Q(DOUT[4]), .QN(n37) );
  DFFS_X1 \reg_mem_reg[3]  ( .D(n68), .CK(CLK), .SN(n21), .Q(DOUT[3]), .QN(n36) );
  DFFS_X1 \reg_mem_reg[2]  ( .D(n67), .CK(CLK), .SN(n21), .Q(DOUT[2]), .QN(n35) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n66), .CK(CLK), .RN(n21), .Q(DOUT[1]), .QN(n34) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n65), .CK(CLK), .RN(n21), .Q(DOUT[0]), .QN(n33) );
  BUF_X1 U2 ( .A(RST_AN), .Z(n21) );
  BUF_X1 U3 ( .A(RST_AN), .Z(n22) );
  BUF_X1 U4 ( .A(RST_AN), .Z(n23) );
  OAI21_X1 U5 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X1 U6 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U7 ( .B1(n48), .B2(EN), .A(n16), .ZN(n80) );
  NAND2_X1 U8 ( .A1(DIN[15]), .A2(EN), .ZN(n16) );
  OAI21_X1 U9 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X1 U10 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U11 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X1 U12 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X1 U13 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  NAND2_X1 U14 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U15 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  NAND2_X1 U16 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X1 U17 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X1 U18 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  OAI21_X1 U19 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  NAND2_X1 U20 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  OAI21_X1 U21 ( .B1(n41), .B2(EN), .A(n9), .ZN(n73) );
  NAND2_X1 U22 ( .A1(DIN[8]), .A2(EN), .ZN(n9) );
  OAI21_X1 U23 ( .B1(n42), .B2(EN), .A(n10), .ZN(n74) );
  NAND2_X1 U24 ( .A1(DIN[9]), .A2(EN), .ZN(n10) );
  OAI21_X1 U25 ( .B1(n43), .B2(EN), .A(n11), .ZN(n75) );
  NAND2_X1 U26 ( .A1(DIN[10]), .A2(EN), .ZN(n11) );
  OAI21_X1 U27 ( .B1(n44), .B2(EN), .A(n12), .ZN(n76) );
  NAND2_X1 U28 ( .A1(DIN[11]), .A2(EN), .ZN(n12) );
  OAI21_X1 U29 ( .B1(n45), .B2(EN), .A(n13), .ZN(n77) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n13) );
  OAI21_X1 U31 ( .B1(n46), .B2(EN), .A(n14), .ZN(n78) );
  NAND2_X1 U32 ( .A1(DIN[13]), .A2(EN), .ZN(n14) );
  OAI21_X1 U33 ( .B1(n47), .B2(EN), .A(n15), .ZN(n79) );
  NAND2_X1 U34 ( .A1(DIN[14]), .A2(EN), .ZN(n15) );
  OAI21_X1 U35 ( .B1(n49), .B2(EN), .A(n17), .ZN(n81) );
  NAND2_X1 U36 ( .A1(DIN[16]), .A2(EN), .ZN(n17) );
  OAI21_X1 U37 ( .B1(n50), .B2(EN), .A(n18), .ZN(n82) );
  NAND2_X1 U38 ( .A1(DIN[17]), .A2(EN), .ZN(n18) );
  OAI21_X1 U39 ( .B1(n51), .B2(EN), .A(n19), .ZN(n83) );
  NAND2_X1 U40 ( .A1(DIN[18]), .A2(EN), .ZN(n19) );
  OAI21_X1 U41 ( .B1(n52), .B2(EN), .A(n20), .ZN(n84) );
  NAND2_X1 U42 ( .A1(DIN[19]), .A2(EN), .ZN(n20) );
  OAI21_X1 U43 ( .B1(n64), .B2(EN), .A(n32), .ZN(n96) );
  NAND2_X1 U44 ( .A1(DIN[31]), .A2(EN), .ZN(n32) );
  OAI21_X1 U45 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X1 U46 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  MUX2_X1 U47 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n85) );
  MUX2_X1 U48 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n86) );
  MUX2_X1 U49 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n87) );
  MUX2_X1 U50 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n88) );
  MUX2_X1 U51 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n89) );
  MUX2_X1 U52 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n90) );
  MUX2_X1 U53 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n91) );
  MUX2_X1 U54 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n92) );
  MUX2_X1 U55 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n93) );
  MUX2_X1 U56 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n94) );
  MUX2_X1 U57 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n95) );
endmodule


module REG_PIPO_32_00000000_00000000_23 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n174), .Q(DOUT[31]), 
        .QN(n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n174), .Q(DOUT[30]), 
        .QN(n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n174), .Q(DOUT[29]), 
        .QN(n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n174), .Q(DOUT[28]), 
        .QN(n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n174), .Q(DOUT[27]), 
        .QN(n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n174), .Q(DOUT[26]), 
        .QN(n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n174), .Q(DOUT[25]), 
        .QN(n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n174), .Q(DOUT[24]), 
        .QN(n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n174), .Q(DOUT[23]), 
        .QN(n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n174), .Q(DOUT[22]), 
        .QN(n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n173), .Q(DOUT[21]), 
        .QN(n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n173), .Q(DOUT[20]), 
        .QN(n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n173), .Q(DOUT[19]), 
        .QN(n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n173), .Q(DOUT[18]), 
        .QN(n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n173), .Q(DOUT[17]), 
        .QN(n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n173), .Q(DOUT[16]), 
        .QN(n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n173), .Q(DOUT[15]), 
        .QN(n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n173), .Q(DOUT[14]), 
        .QN(n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n173), .Q(DOUT[13]), 
        .QN(n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n173), .Q(DOUT[12]), 
        .QN(n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n173), .Q(DOUT[11]), 
        .QN(n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n172), .Q(DOUT[10]), 
        .QN(n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n172), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n172), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n172), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n172), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n172), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n172), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n172), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n172), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n172), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n172), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n170) );
  BUF_X1 U3 ( .A(n169), .Z(n171) );
  BUF_X1 U4 ( .A(RST_AN), .Z(n172) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  OAI22_X1 U7 ( .A1(n168), .A2(EN), .B1(n171), .B2(n207), .ZN(n136) );
  INV_X1 U8 ( .A(DIN[0]), .ZN(n207) );
  OAI22_X1 U9 ( .A1(n167), .A2(EN), .B1(n171), .B2(n206), .ZN(n135) );
  INV_X1 U10 ( .A(DIN[1]), .ZN(n206) );
  OAI22_X1 U11 ( .A1(n166), .A2(EN), .B1(n170), .B2(n205), .ZN(n134) );
  INV_X1 U12 ( .A(DIN[2]), .ZN(n205) );
  OAI22_X1 U13 ( .A1(n165), .A2(EN), .B1(n170), .B2(n204), .ZN(n133) );
  INV_X1 U14 ( .A(DIN[3]), .ZN(n204) );
  OAI22_X1 U15 ( .A1(n164), .A2(EN), .B1(n171), .B2(n203), .ZN(n132) );
  INV_X1 U16 ( .A(DIN[4]), .ZN(n203) );
  OAI22_X1 U17 ( .A1(n163), .A2(EN), .B1(n171), .B2(n202), .ZN(n131) );
  INV_X1 U18 ( .A(DIN[5]), .ZN(n202) );
  OAI22_X1 U19 ( .A1(n162), .A2(EN), .B1(n170), .B2(n201), .ZN(n130) );
  INV_X1 U20 ( .A(DIN[6]), .ZN(n201) );
  OAI22_X1 U21 ( .A1(n161), .A2(EN), .B1(n170), .B2(n200), .ZN(n129) );
  INV_X1 U22 ( .A(DIN[7]), .ZN(n200) );
  OAI22_X1 U23 ( .A1(n160), .A2(EN), .B1(n171), .B2(n199), .ZN(n128) );
  INV_X1 U24 ( .A(DIN[8]), .ZN(n199) );
  OAI22_X1 U25 ( .A1(n159), .A2(EN), .B1(n171), .B2(n198), .ZN(n127) );
  INV_X1 U26 ( .A(DIN[9]), .ZN(n198) );
  OAI22_X1 U27 ( .A1(n158), .A2(EN), .B1(n170), .B2(n197), .ZN(n126) );
  INV_X1 U28 ( .A(DIN[10]), .ZN(n197) );
  OAI22_X1 U29 ( .A1(n157), .A2(EN), .B1(n170), .B2(n196), .ZN(n125) );
  INV_X1 U30 ( .A(DIN[11]), .ZN(n196) );
  OAI22_X1 U31 ( .A1(n156), .A2(EN), .B1(n171), .B2(n195), .ZN(n124) );
  INV_X1 U32 ( .A(DIN[12]), .ZN(n195) );
  OAI22_X1 U33 ( .A1(n155), .A2(EN), .B1(n171), .B2(n194), .ZN(n123) );
  INV_X1 U34 ( .A(DIN[13]), .ZN(n194) );
  OAI22_X1 U35 ( .A1(n154), .A2(EN), .B1(n170), .B2(n193), .ZN(n122) );
  INV_X1 U36 ( .A(DIN[14]), .ZN(n193) );
  OAI22_X1 U37 ( .A1(n153), .A2(EN), .B1(n170), .B2(n192), .ZN(n121) );
  INV_X1 U38 ( .A(DIN[15]), .ZN(n192) );
  OAI22_X1 U39 ( .A1(n152), .A2(EN), .B1(n171), .B2(n191), .ZN(n120) );
  INV_X1 U40 ( .A(DIN[16]), .ZN(n191) );
  OAI22_X1 U41 ( .A1(n151), .A2(EN), .B1(n171), .B2(n190), .ZN(n119) );
  INV_X1 U42 ( .A(DIN[17]), .ZN(n190) );
  OAI22_X1 U43 ( .A1(n150), .A2(EN), .B1(n170), .B2(n189), .ZN(n118) );
  INV_X1 U44 ( .A(DIN[18]), .ZN(n189) );
  OAI22_X1 U45 ( .A1(n149), .A2(EN), .B1(n170), .B2(n188), .ZN(n117) );
  INV_X1 U46 ( .A(DIN[19]), .ZN(n188) );
  OAI22_X1 U47 ( .A1(n137), .A2(EN), .B1(n170), .B2(n208), .ZN(n105) );
  INV_X1 U48 ( .A(DIN[31]), .ZN(n208) );
  INV_X1 U49 ( .A(EN), .ZN(n175) );
  OR2_X1 U50 ( .A1(INIT), .A2(n175), .ZN(n169) );
  INV_X1 U51 ( .A(n169), .ZN(n186) );
  NAND2_X1 U52 ( .A1(DIN[20]), .A2(n186), .ZN(n176) );
  OAI21_X1 U53 ( .B1(n148), .B2(EN), .A(n176), .ZN(n116) );
  NAND2_X1 U54 ( .A1(DIN[21]), .A2(n186), .ZN(n177) );
  OAI21_X1 U55 ( .B1(n147), .B2(EN), .A(n177), .ZN(n115) );
  NAND2_X1 U56 ( .A1(DIN[22]), .A2(n186), .ZN(n178) );
  OAI21_X1 U57 ( .B1(n146), .B2(EN), .A(n178), .ZN(n114) );
  NAND2_X1 U58 ( .A1(DIN[23]), .A2(n186), .ZN(n179) );
  OAI21_X1 U59 ( .B1(n145), .B2(EN), .A(n179), .ZN(n113) );
  NAND2_X1 U60 ( .A1(DIN[24]), .A2(n186), .ZN(n180) );
  OAI21_X1 U61 ( .B1(n144), .B2(EN), .A(n180), .ZN(n112) );
  NAND2_X1 U62 ( .A1(DIN[25]), .A2(n186), .ZN(n181) );
  OAI21_X1 U63 ( .B1(n143), .B2(EN), .A(n181), .ZN(n111) );
  NAND2_X1 U64 ( .A1(DIN[26]), .A2(n186), .ZN(n182) );
  OAI21_X1 U65 ( .B1(n142), .B2(EN), .A(n182), .ZN(n110) );
  NAND2_X1 U66 ( .A1(DIN[27]), .A2(n186), .ZN(n183) );
  OAI21_X1 U67 ( .B1(n141), .B2(EN), .A(n183), .ZN(n109) );
  NAND2_X1 U68 ( .A1(DIN[28]), .A2(n186), .ZN(n184) );
  OAI21_X1 U69 ( .B1(n140), .B2(EN), .A(n184), .ZN(n108) );
  NAND2_X1 U70 ( .A1(DIN[29]), .A2(n186), .ZN(n185) );
  OAI21_X1 U71 ( .B1(n139), .B2(EN), .A(n185), .ZN(n107) );
  NAND2_X1 U72 ( .A1(DIN[30]), .A2(n186), .ZN(n187) );
  OAI21_X1 U73 ( .B1(n138), .B2(EN), .A(n187), .ZN(n106) );
endmodule


module REG_PIPO_32_00000000_00000000_22 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module RF_ADDR_W5_DATA_W32_1 ( CLK, RST_AN, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST_AN, ENABLE, RD1, RD2, WR;
  wire   \registers[1][31] , \registers[1][30] , \registers[1][29] ,
         \registers[1][28] , \registers[1][27] , \registers[1][26] ,
         \registers[1][25] , \registers[1][24] , \registers[1][23] ,
         \registers[1][22] , \registers[1][21] , \registers[1][20] ,
         \registers[1][19] , \registers[1][18] , \registers[1][17] ,
         \registers[1][16] , \registers[1][15] , \registers[1][14] ,
         \registers[1][13] , \registers[1][12] , \registers[1][11] ,
         \registers[1][10] , \registers[1][9] , \registers[1][8] ,
         \registers[1][7] , \registers[1][6] , \registers[1][5] ,
         \registers[1][4] , \registers[1][3] , \registers[1][2] ,
         \registers[1][1] , \registers[1][0] , \registers[6][31] ,
         \registers[6][30] , \registers[6][29] , \registers[6][28] ,
         \registers[6][27] , \registers[6][26] , \registers[6][25] ,
         \registers[6][24] , \registers[6][23] , \registers[6][22] ,
         \registers[6][21] , \registers[6][20] , \registers[6][19] ,
         \registers[6][18] , \registers[6][17] , \registers[6][16] ,
         \registers[6][15] , \registers[6][14] , \registers[6][13] ,
         \registers[6][12] , \registers[6][11] , \registers[6][10] ,
         \registers[6][9] , \registers[6][8] , \registers[6][7] ,
         \registers[6][6] , \registers[6][5] , \registers[6][4] ,
         \registers[6][3] , \registers[6][2] , \registers[6][1] ,
         \registers[6][0] , \registers[7][31] , \registers[7][30] ,
         \registers[7][29] , \registers[7][28] , \registers[7][27] ,
         \registers[7][26] , \registers[7][25] , \registers[7][24] ,
         \registers[7][23] , \registers[7][22] , \registers[7][21] ,
         \registers[7][20] , \registers[7][19] , \registers[7][18] ,
         \registers[7][17] , \registers[7][16] , \registers[7][15] ,
         \registers[7][14] , \registers[7][13] , \registers[7][12] ,
         \registers[7][11] , \registers[7][10] , \registers[7][9] ,
         \registers[7][8] , \registers[7][7] , \registers[7][6] ,
         \registers[7][5] , \registers[7][4] , \registers[7][3] ,
         \registers[7][2] , \registers[7][1] , \registers[7][0] ,
         \registers[8][31] , \registers[8][30] , \registers[8][29] ,
         \registers[8][28] , \registers[8][27] , \registers[8][26] ,
         \registers[8][25] , \registers[8][24] , \registers[8][23] ,
         \registers[8][22] , \registers[8][21] , \registers[8][20] ,
         \registers[8][19] , \registers[8][18] , \registers[8][17] ,
         \registers[8][16] , \registers[8][15] , \registers[8][14] ,
         \registers[8][13] , \registers[8][12] , \registers[8][11] ,
         \registers[8][10] , \registers[8][9] , \registers[8][8] ,
         \registers[8][7] , \registers[8][6] , \registers[8][5] ,
         \registers[8][4] , \registers[8][3] , \registers[8][2] ,
         \registers[8][1] , \registers[8][0] , \registers[9][31] ,
         \registers[9][30] , \registers[9][29] , \registers[9][28] ,
         \registers[9][27] , \registers[9][26] , \registers[9][25] ,
         \registers[9][24] , \registers[9][23] , \registers[9][22] ,
         \registers[9][21] , \registers[9][20] , \registers[9][19] ,
         \registers[9][18] , \registers[9][17] , \registers[9][16] ,
         \registers[9][15] , \registers[9][14] , \registers[9][13] ,
         \registers[9][12] , \registers[9][11] , \registers[9][10] ,
         \registers[9][9] , \registers[9][8] , \registers[9][7] ,
         \registers[9][6] , \registers[9][5] , \registers[9][4] ,
         \registers[9][3] , \registers[9][2] , \registers[9][1] ,
         \registers[9][0] , \registers[12][31] , \registers[12][30] ,
         \registers[12][29] , \registers[12][28] , \registers[12][27] ,
         \registers[12][26] , \registers[12][25] , \registers[12][24] ,
         \registers[12][23] , \registers[12][22] , \registers[12][21] ,
         \registers[12][20] , \registers[12][19] , \registers[12][18] ,
         \registers[12][17] , \registers[12][16] , \registers[12][15] ,
         \registers[12][14] , \registers[12][13] , \registers[12][12] ,
         \registers[12][11] , \registers[12][10] , \registers[12][9] ,
         \registers[12][8] , \registers[12][7] , \registers[12][6] ,
         \registers[12][5] , \registers[12][4] , \registers[12][3] ,
         \registers[12][2] , \registers[12][1] , \registers[12][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[18][31] ,
         \registers[18][30] , \registers[18][29] , \registers[18][28] ,
         \registers[18][27] , \registers[18][26] , \registers[18][25] ,
         \registers[18][24] , \registers[18][23] , \registers[18][22] ,
         \registers[18][21] , \registers[18][20] , \registers[18][19] ,
         \registers[18][18] , \registers[18][17] , \registers[18][16] ,
         \registers[18][15] , \registers[18][14] , \registers[18][13] ,
         \registers[18][12] , \registers[18][11] , \registers[18][10] ,
         \registers[18][9] , \registers[18][8] , \registers[18][7] ,
         \registers[18][6] , \registers[18][5] , \registers[18][4] ,
         \registers[18][3] , \registers[18][2] , \registers[18][1] ,
         \registers[18][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[22][31] , \registers[22][30] , \registers[22][29] ,
         \registers[22][28] , \registers[22][27] , \registers[22][26] ,
         \registers[22][25] , \registers[22][24] , \registers[22][23] ,
         \registers[22][22] , \registers[22][21] , \registers[22][20] ,
         \registers[22][19] , \registers[22][18] , \registers[22][17] ,
         \registers[22][16] , \registers[22][15] , \registers[22][14] ,
         \registers[22][13] , \registers[22][12] , \registers[22][11] ,
         \registers[22][10] , \registers[22][9] , \registers[22][8] ,
         \registers[22][7] , \registers[22][6] , \registers[22][5] ,
         \registers[22][4] , \registers[22][3] , \registers[22][2] ,
         \registers[22][1] , \registers[22][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[24][31] , \registers[24][30] ,
         \registers[24][29] , \registers[24][28] , \registers[24][27] ,
         \registers[24][26] , \registers[24][25] , \registers[24][24] ,
         \registers[24][23] , \registers[24][22] , \registers[24][21] ,
         \registers[24][20] , \registers[24][19] , \registers[24][18] ,
         \registers[24][17] , \registers[24][16] , \registers[24][15] ,
         \registers[24][14] , \registers[24][13] , \registers[24][12] ,
         \registers[24][11] , \registers[24][10] , \registers[24][9] ,
         \registers[24][8] , \registers[24][7] , \registers[24][6] ,
         \registers[24][5] , \registers[24][4] , \registers[24][3] ,
         \registers[24][2] , \registers[24][1] , \registers[24][0] ,
         \registers[25][31] , \registers[25][30] , \registers[25][29] ,
         \registers[25][28] , \registers[25][27] , \registers[25][26] ,
         \registers[25][25] , \registers[25][24] , \registers[25][23] ,
         \registers[25][22] , \registers[25][21] , \registers[25][20] ,
         \registers[25][19] , \registers[25][18] , \registers[25][17] ,
         \registers[25][16] , \registers[25][15] , \registers[25][14] ,
         \registers[25][13] , \registers[25][12] , \registers[25][11] ,
         \registers[25][10] , \registers[25][9] , \registers[25][8] ,
         \registers[25][7] , \registers[25][6] , \registers[25][5] ,
         \registers[25][4] , \registers[25][3] , \registers[25][2] ,
         \registers[25][1] , \registers[25][0] , \registers[28][31] ,
         \registers[28][30] , \registers[28][29] , \registers[28][28] ,
         \registers[28][27] , \registers[28][26] , \registers[28][25] ,
         \registers[28][24] , \registers[28][23] , \registers[28][22] ,
         \registers[28][21] , \registers[28][20] , \registers[28][19] ,
         \registers[28][18] , \registers[28][17] , \registers[28][16] ,
         \registers[28][15] , \registers[28][14] , \registers[28][13] ,
         \registers[28][12] , \registers[28][11] , \registers[28][10] ,
         \registers[28][9] , \registers[28][8] , \registers[28][7] ,
         \registers[28][6] , \registers[28][5] , \registers[28][4] ,
         \registers[28][3] , \registers[28][2] , \registers[28][1] ,
         \registers[28][0] , \registers[29][31] , \registers[29][30] ,
         \registers[29][29] , \registers[29][28] , \registers[29][27] ,
         \registers[29][26] , \registers[29][25] , \registers[29][24] ,
         \registers[29][23] , \registers[29][22] , \registers[29][21] ,
         \registers[29][20] , \registers[29][19] , \registers[29][18] ,
         \registers[29][17] , \registers[29][16] , \registers[29][15] ,
         \registers[29][14] , \registers[29][13] , \registers[29][12] ,
         \registers[29][11] , \registers[29][10] , \registers[29][9] ,
         \registers[29][8] , \registers[29][7] , \registers[29][6] ,
         \registers[29][5] , \registers[29][4] , \registers[29][3] ,
         \registers[29][2] , \registers[29][1] , \registers[29][0] , N82, N185,
         N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1113, n1115, n1117, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1156, n1157, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1432, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1112, n1114, n1116, n1118, n1155, n1158,
         n1225, n1226, n1361, n1362, n1429, n1430, n1431, n1433, n1500, n1501,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844;

  DFFR_X1 \registers_reg[1][31]  ( .D(n3513), .CK(CLK), .RN(n3305), .Q(
        \registers[1][31] ) );
  DFFR_X1 \registers_reg[1][30]  ( .D(n3512), .CK(CLK), .RN(n3305), .Q(
        \registers[1][30] ) );
  DFFR_X1 \registers_reg[1][29]  ( .D(n3511), .CK(CLK), .RN(n3304), .Q(
        \registers[1][29] ) );
  DFFR_X1 \registers_reg[1][28]  ( .D(n3510), .CK(CLK), .RN(n3304), .Q(
        \registers[1][28] ) );
  DFFR_X1 \registers_reg[1][27]  ( .D(n3509), .CK(CLK), .RN(n3304), .Q(
        \registers[1][27] ) );
  DFFR_X1 \registers_reg[1][26]  ( .D(n3508), .CK(CLK), .RN(n3304), .Q(
        \registers[1][26] ) );
  DFFR_X1 \registers_reg[1][25]  ( .D(n3507), .CK(CLK), .RN(n3304), .Q(
        \registers[1][25] ) );
  DFFR_X1 \registers_reg[1][24]  ( .D(n3506), .CK(CLK), .RN(n3304), .Q(
        \registers[1][24] ) );
  DFFR_X1 \registers_reg[1][23]  ( .D(n3505), .CK(CLK), .RN(n3304), .Q(
        \registers[1][23] ) );
  DFFR_X1 \registers_reg[1][22]  ( .D(n3504), .CK(CLK), .RN(n3304), .Q(
        \registers[1][22] ) );
  DFFR_X1 \registers_reg[1][21]  ( .D(n3503), .CK(CLK), .RN(n3304), .Q(
        \registers[1][21] ) );
  DFFR_X1 \registers_reg[1][20]  ( .D(n3502), .CK(CLK), .RN(n3304), .Q(
        \registers[1][20] ) );
  DFFR_X1 \registers_reg[1][19]  ( .D(n3501), .CK(CLK), .RN(n3304), .Q(
        \registers[1][19] ) );
  DFFR_X1 \registers_reg[1][18]  ( .D(n3500), .CK(CLK), .RN(n3303), .Q(
        \registers[1][18] ) );
  DFFR_X1 \registers_reg[1][17]  ( .D(n3499), .CK(CLK), .RN(n3303), .Q(
        \registers[1][17] ) );
  DFFR_X1 \registers_reg[1][16]  ( .D(n3498), .CK(CLK), .RN(n3303), .Q(
        \registers[1][16] ) );
  DFFR_X1 \registers_reg[1][15]  ( .D(n3497), .CK(CLK), .RN(n3303), .Q(
        \registers[1][15] ) );
  DFFR_X1 \registers_reg[1][14]  ( .D(n3496), .CK(CLK), .RN(n3303), .Q(
        \registers[1][14] ) );
  DFFR_X1 \registers_reg[1][13]  ( .D(n3495), .CK(CLK), .RN(n3303), .Q(
        \registers[1][13] ) );
  DFFR_X1 \registers_reg[1][12]  ( .D(n3494), .CK(CLK), .RN(n3303), .Q(
        \registers[1][12] ) );
  DFFR_X1 \registers_reg[1][11]  ( .D(n3493), .CK(CLK), .RN(n3303), .Q(
        \registers[1][11] ) );
  DFFR_X1 \registers_reg[1][10]  ( .D(n3492), .CK(CLK), .RN(n3303), .Q(
        \registers[1][10] ) );
  DFFR_X1 \registers_reg[1][9]  ( .D(n3491), .CK(CLK), .RN(n3303), .Q(
        \registers[1][9] ) );
  DFFR_X1 \registers_reg[1][8]  ( .D(n3490), .CK(CLK), .RN(n3303), .Q(
        \registers[1][8] ) );
  DFFR_X1 \registers_reg[1][7]  ( .D(n3489), .CK(CLK), .RN(n3302), .Q(
        \registers[1][7] ) );
  DFFR_X1 \registers_reg[1][6]  ( .D(n3488), .CK(CLK), .RN(n3302), .Q(
        \registers[1][6] ) );
  DFFR_X1 \registers_reg[1][5]  ( .D(n3487), .CK(CLK), .RN(n3302), .Q(
        \registers[1][5] ) );
  DFFR_X1 \registers_reg[1][4]  ( .D(n3486), .CK(CLK), .RN(n3302), .Q(
        \registers[1][4] ) );
  DFFR_X1 \registers_reg[1][3]  ( .D(n3485), .CK(CLK), .RN(n3302), .Q(
        \registers[1][3] ) );
  DFFR_X1 \registers_reg[1][2]  ( .D(n3484), .CK(CLK), .RN(n3302), .Q(
        \registers[1][2] ) );
  DFFR_X1 \registers_reg[1][1]  ( .D(n3483), .CK(CLK), .RN(n3302), .Q(
        \registers[1][1] ) );
  DFFR_X1 \registers_reg[1][0]  ( .D(n3482), .CK(CLK), .RN(n3302), .Q(
        \registers[1][0] ) );
  DFFR_X1 \registers_reg[2][31]  ( .D(n3284), .CK(CLK), .RN(n3302), .QN(n33)
         );
  DFFR_X1 \registers_reg[2][30]  ( .D(n3283), .CK(CLK), .RN(n3302), .QN(n34)
         );
  DFFR_X1 \registers_reg[2][29]  ( .D(n3282), .CK(CLK), .RN(n3302), .QN(n35)
         );
  DFFR_X1 \registers_reg[2][28]  ( .D(n3281), .CK(CLK), .RN(n3301), .QN(n36)
         );
  DFFR_X1 \registers_reg[2][27]  ( .D(n3280), .CK(CLK), .RN(n3301), .QN(n37)
         );
  DFFR_X1 \registers_reg[2][26]  ( .D(n3279), .CK(CLK), .RN(n3301), .QN(n38)
         );
  DFFR_X1 \registers_reg[2][25]  ( .D(n3278), .CK(CLK), .RN(n3301), .QN(n39)
         );
  DFFR_X1 \registers_reg[2][24]  ( .D(n3277), .CK(CLK), .RN(n3301), .QN(n40)
         );
  DFFR_X1 \registers_reg[2][23]  ( .D(n3276), .CK(CLK), .RN(n3301), .QN(n41)
         );
  DFFR_X1 \registers_reg[2][22]  ( .D(n3275), .CK(CLK), .RN(n3301), .QN(n42)
         );
  DFFR_X1 \registers_reg[2][21]  ( .D(n3274), .CK(CLK), .RN(n3301), .QN(n43)
         );
  DFFR_X1 \registers_reg[2][20]  ( .D(n3273), .CK(CLK), .RN(n3301), .QN(n44)
         );
  DFFR_X1 \registers_reg[2][19]  ( .D(n3272), .CK(CLK), .RN(n3301), .QN(n45)
         );
  DFFR_X1 \registers_reg[2][18]  ( .D(n3271), .CK(CLK), .RN(n3301), .QN(n46)
         );
  DFFR_X1 \registers_reg[2][17]  ( .D(n3270), .CK(CLK), .RN(n3300), .QN(n47)
         );
  DFFR_X1 \registers_reg[2][16]  ( .D(n3269), .CK(CLK), .RN(n3300), .QN(n48)
         );
  DFFR_X1 \registers_reg[2][15]  ( .D(n3268), .CK(CLK), .RN(n3300), .QN(n49)
         );
  DFFR_X1 \registers_reg[2][14]  ( .D(n3267), .CK(CLK), .RN(n3300), .QN(n50)
         );
  DFFR_X1 \registers_reg[2][13]  ( .D(n3266), .CK(CLK), .RN(n3300), .QN(n51)
         );
  DFFR_X1 \registers_reg[2][12]  ( .D(n3265), .CK(CLK), .RN(n3300), .QN(n52)
         );
  DFFR_X1 \registers_reg[2][11]  ( .D(n3264), .CK(CLK), .RN(n3300), .QN(n53)
         );
  DFFR_X1 \registers_reg[2][10]  ( .D(n3263), .CK(CLK), .RN(n3300), .QN(n54)
         );
  DFFR_X1 \registers_reg[2][9]  ( .D(n3262), .CK(CLK), .RN(n3300), .QN(n55) );
  DFFR_X1 \registers_reg[2][8]  ( .D(n3261), .CK(CLK), .RN(n3300), .QN(n56) );
  DFFR_X1 \registers_reg[2][7]  ( .D(n3260), .CK(CLK), .RN(n3300), .QN(n57) );
  DFFR_X1 \registers_reg[2][6]  ( .D(n3259), .CK(CLK), .RN(n3299), .QN(n58) );
  DFFR_X1 \registers_reg[2][5]  ( .D(n3258), .CK(CLK), .RN(n3299), .QN(n59) );
  DFFR_X1 \registers_reg[2][4]  ( .D(n3257), .CK(CLK), .RN(n3299), .QN(n60) );
  DFFR_X1 \registers_reg[2][3]  ( .D(n3256), .CK(CLK), .RN(n3299), .QN(n61) );
  DFFR_X1 \registers_reg[2][2]  ( .D(n3255), .CK(CLK), .RN(n3299), .QN(n62) );
  DFFR_X1 \registers_reg[2][1]  ( .D(n3254), .CK(CLK), .RN(n3299), .QN(n63) );
  DFFR_X1 \registers_reg[2][0]  ( .D(n3253), .CK(CLK), .RN(n3299), .QN(n64) );
  DFFR_X1 \registers_reg[3][31]  ( .D(n3252), .CK(CLK), .RN(n3299), .QN(n65)
         );
  DFFR_X1 \registers_reg[3][30]  ( .D(n3251), .CK(CLK), .RN(n3299), .QN(n66)
         );
  DFFR_X1 \registers_reg[3][29]  ( .D(n3250), .CK(CLK), .RN(n3299), .QN(n67)
         );
  DFFR_X1 \registers_reg[3][28]  ( .D(n3249), .CK(CLK), .RN(n3299), .QN(n68)
         );
  DFFR_X1 \registers_reg[3][27]  ( .D(n3248), .CK(CLK), .RN(n3298), .QN(n69)
         );
  DFFR_X1 \registers_reg[3][26]  ( .D(n3247), .CK(CLK), .RN(n3298), .QN(n70)
         );
  DFFR_X1 \registers_reg[3][25]  ( .D(n3246), .CK(CLK), .RN(n3298), .QN(n71)
         );
  DFFR_X1 \registers_reg[3][24]  ( .D(n3245), .CK(CLK), .RN(n3298), .QN(n72)
         );
  DFFR_X1 \registers_reg[3][23]  ( .D(n3244), .CK(CLK), .RN(n3298), .QN(n73)
         );
  DFFR_X1 \registers_reg[3][22]  ( .D(n3243), .CK(CLK), .RN(n3298), .QN(n74)
         );
  DFFR_X1 \registers_reg[3][21]  ( .D(n3242), .CK(CLK), .RN(n3298), .QN(n75)
         );
  DFFR_X1 \registers_reg[3][20]  ( .D(n3241), .CK(CLK), .RN(n3298), .QN(n76)
         );
  DFFR_X1 \registers_reg[3][19]  ( .D(n3240), .CK(CLK), .RN(n3298), .QN(n77)
         );
  DFFR_X1 \registers_reg[3][18]  ( .D(n3239), .CK(CLK), .RN(n3298), .QN(n78)
         );
  DFFR_X1 \registers_reg[3][17]  ( .D(n3238), .CK(CLK), .RN(n3298), .QN(n79)
         );
  DFFR_X1 \registers_reg[3][16]  ( .D(n3237), .CK(CLK), .RN(n3297), .QN(n80)
         );
  DFFR_X1 \registers_reg[3][15]  ( .D(n3236), .CK(CLK), .RN(n3297), .QN(n81)
         );
  DFFR_X1 \registers_reg[3][14]  ( .D(n3235), .CK(CLK), .RN(n3297), .QN(n82)
         );
  DFFR_X1 \registers_reg[3][13]  ( .D(n3234), .CK(CLK), .RN(n3297), .QN(n83)
         );
  DFFR_X1 \registers_reg[3][12]  ( .D(n3233), .CK(CLK), .RN(n3297), .QN(n84)
         );
  DFFR_X1 \registers_reg[3][11]  ( .D(n3232), .CK(CLK), .RN(n3297), .QN(n85)
         );
  DFFR_X1 \registers_reg[3][10]  ( .D(n3231), .CK(CLK), .RN(n3297), .QN(n86)
         );
  DFFR_X1 \registers_reg[3][9]  ( .D(n3230), .CK(CLK), .RN(n3297), .QN(n87) );
  DFFR_X1 \registers_reg[3][8]  ( .D(n3229), .CK(CLK), .RN(n3297), .QN(n88) );
  DFFR_X1 \registers_reg[3][7]  ( .D(n3228), .CK(CLK), .RN(n3297), .QN(n89) );
  DFFR_X1 \registers_reg[3][6]  ( .D(n3227), .CK(CLK), .RN(n3297), .QN(n90) );
  DFFR_X1 \registers_reg[3][5]  ( .D(n3226), .CK(CLK), .RN(n3296), .QN(n91) );
  DFFR_X1 \registers_reg[3][4]  ( .D(n3225), .CK(CLK), .RN(n3296), .QN(n92) );
  DFFR_X1 \registers_reg[3][3]  ( .D(n3224), .CK(CLK), .RN(n3296), .QN(n93) );
  DFFR_X1 \registers_reg[3][2]  ( .D(n3223), .CK(CLK), .RN(n3296), .QN(n94) );
  DFFR_X1 \registers_reg[3][1]  ( .D(n3222), .CK(CLK), .RN(n3296), .QN(n95) );
  DFFR_X1 \registers_reg[3][0]  ( .D(n3221), .CK(CLK), .RN(n3296), .QN(n96) );
  DFFR_X1 \registers_reg[4][31]  ( .D(n3220), .CK(CLK), .RN(n3296), .QN(n97)
         );
  DFFR_X1 \registers_reg[4][30]  ( .D(n3219), .CK(CLK), .RN(n3296), .QN(n98)
         );
  DFFR_X1 \registers_reg[4][29]  ( .D(n3218), .CK(CLK), .RN(n3296), .QN(n99)
         );
  DFFR_X1 \registers_reg[4][28]  ( .D(n3217), .CK(CLK), .RN(n3296), .QN(n100)
         );
  DFFR_X1 \registers_reg[4][27]  ( .D(n3216), .CK(CLK), .RN(n3296), .QN(n101)
         );
  DFFR_X1 \registers_reg[4][26]  ( .D(n3215), .CK(CLK), .RN(n3295), .QN(n102)
         );
  DFFR_X1 \registers_reg[4][25]  ( .D(n3214), .CK(CLK), .RN(n3295), .QN(n103)
         );
  DFFR_X1 \registers_reg[4][24]  ( .D(n3213), .CK(CLK), .RN(n3295), .QN(n104)
         );
  DFFR_X1 \registers_reg[4][23]  ( .D(n3212), .CK(CLK), .RN(n3295), .QN(n105)
         );
  DFFR_X1 \registers_reg[4][22]  ( .D(n3211), .CK(CLK), .RN(n3295), .QN(n106)
         );
  DFFR_X1 \registers_reg[4][21]  ( .D(n3210), .CK(CLK), .RN(n3295), .QN(n107)
         );
  DFFR_X1 \registers_reg[4][20]  ( .D(n3209), .CK(CLK), .RN(n3295), .QN(n108)
         );
  DFFR_X1 \registers_reg[4][19]  ( .D(n3208), .CK(CLK), .RN(n3295), .QN(n109)
         );
  DFFR_X1 \registers_reg[4][18]  ( .D(n3207), .CK(CLK), .RN(n3295), .QN(n110)
         );
  DFFR_X1 \registers_reg[4][17]  ( .D(n3206), .CK(CLK), .RN(n3295), .QN(n111)
         );
  DFFR_X1 \registers_reg[4][16]  ( .D(n3205), .CK(CLK), .RN(n3295), .QN(n112)
         );
  DFFR_X1 \registers_reg[4][15]  ( .D(n3204), .CK(CLK), .RN(n3294), .QN(n113)
         );
  DFFR_X1 \registers_reg[4][14]  ( .D(n3203), .CK(CLK), .RN(n3294), .QN(n114)
         );
  DFFR_X1 \registers_reg[4][13]  ( .D(n3202), .CK(CLK), .RN(n3294), .QN(n115)
         );
  DFFR_X1 \registers_reg[4][12]  ( .D(n3201), .CK(CLK), .RN(n3294), .QN(n116)
         );
  DFFR_X1 \registers_reg[4][11]  ( .D(n3200), .CK(CLK), .RN(n3294), .QN(n117)
         );
  DFFR_X1 \registers_reg[4][10]  ( .D(n3199), .CK(CLK), .RN(n3294), .QN(n118)
         );
  DFFR_X1 \registers_reg[4][9]  ( .D(n3198), .CK(CLK), .RN(n3294), .QN(n119)
         );
  DFFR_X1 \registers_reg[4][8]  ( .D(n3197), .CK(CLK), .RN(n3294), .QN(n120)
         );
  DFFR_X1 \registers_reg[4][7]  ( .D(n3196), .CK(CLK), .RN(n3294), .QN(n121)
         );
  DFFR_X1 \registers_reg[4][6]  ( .D(n3195), .CK(CLK), .RN(n3294), .QN(n122)
         );
  DFFR_X1 \registers_reg[4][5]  ( .D(n3194), .CK(CLK), .RN(n3294), .QN(n123)
         );
  DFFR_X1 \registers_reg[4][4]  ( .D(n3193), .CK(CLK), .RN(n3293), .QN(n124)
         );
  DFFR_X1 \registers_reg[4][3]  ( .D(n3192), .CK(CLK), .RN(n3293), .QN(n125)
         );
  DFFR_X1 \registers_reg[4][2]  ( .D(n3191), .CK(CLK), .RN(n3293), .QN(n126)
         );
  DFFR_X1 \registers_reg[4][1]  ( .D(n3190), .CK(CLK), .RN(n3293), .QN(n127)
         );
  DFFR_X1 \registers_reg[4][0]  ( .D(n3189), .CK(CLK), .RN(n3293), .QN(n128)
         );
  DFFR_X1 \registers_reg[5][31]  ( .D(n3188), .CK(CLK), .RN(n3293), .QN(n129)
         );
  DFFR_X1 \registers_reg[5][30]  ( .D(n3187), .CK(CLK), .RN(n3293), .QN(n130)
         );
  DFFR_X1 \registers_reg[5][29]  ( .D(n3186), .CK(CLK), .RN(n3293), .QN(n131)
         );
  DFFR_X1 \registers_reg[5][28]  ( .D(n3185), .CK(CLK), .RN(n3293), .QN(n132)
         );
  DFFR_X1 \registers_reg[5][27]  ( .D(n3184), .CK(CLK), .RN(n3293), .QN(n133)
         );
  DFFR_X1 \registers_reg[5][26]  ( .D(n3183), .CK(CLK), .RN(n3293), .QN(n134)
         );
  DFFR_X1 \registers_reg[5][25]  ( .D(n3182), .CK(CLK), .RN(n3292), .QN(n135)
         );
  DFFR_X1 \registers_reg[5][24]  ( .D(n3181), .CK(CLK), .RN(n3292), .QN(n136)
         );
  DFFR_X1 \registers_reg[5][23]  ( .D(n3180), .CK(CLK), .RN(n3292), .QN(n137)
         );
  DFFR_X1 \registers_reg[5][22]  ( .D(n3179), .CK(CLK), .RN(n3292), .QN(n138)
         );
  DFFR_X1 \registers_reg[5][21]  ( .D(n3178), .CK(CLK), .RN(n3292), .QN(n139)
         );
  DFFR_X1 \registers_reg[5][20]  ( .D(n3177), .CK(CLK), .RN(n3292), .QN(n140)
         );
  DFFR_X1 \registers_reg[5][19]  ( .D(n3176), .CK(CLK), .RN(n3292), .QN(n141)
         );
  DFFR_X1 \registers_reg[5][18]  ( .D(n3175), .CK(CLK), .RN(n3292), .QN(n142)
         );
  DFFR_X1 \registers_reg[5][17]  ( .D(n3174), .CK(CLK), .RN(n3292), .QN(n143)
         );
  DFFR_X1 \registers_reg[5][16]  ( .D(n3173), .CK(CLK), .RN(n3292), .QN(n144)
         );
  DFFR_X1 \registers_reg[5][15]  ( .D(n3172), .CK(CLK), .RN(n3292), .QN(n145)
         );
  DFFR_X1 \registers_reg[5][14]  ( .D(n3171), .CK(CLK), .RN(n3291), .QN(n146)
         );
  DFFR_X1 \registers_reg[5][13]  ( .D(n3170), .CK(CLK), .RN(n3291), .QN(n147)
         );
  DFFR_X1 \registers_reg[5][12]  ( .D(n3169), .CK(CLK), .RN(n3291), .QN(n148)
         );
  DFFR_X1 \registers_reg[5][11]  ( .D(n3168), .CK(CLK), .RN(n3291), .QN(n149)
         );
  DFFR_X1 \registers_reg[5][10]  ( .D(n3167), .CK(CLK), .RN(n3291), .QN(n150)
         );
  DFFR_X1 \registers_reg[5][9]  ( .D(n3166), .CK(CLK), .RN(n3291), .QN(n151)
         );
  DFFR_X1 \registers_reg[5][8]  ( .D(n3165), .CK(CLK), .RN(n3291), .QN(n152)
         );
  DFFR_X1 \registers_reg[5][7]  ( .D(n3164), .CK(CLK), .RN(n3291), .QN(n153)
         );
  DFFR_X1 \registers_reg[5][6]  ( .D(n3163), .CK(CLK), .RN(n3291), .QN(n154)
         );
  DFFR_X1 \registers_reg[5][5]  ( .D(n3162), .CK(CLK), .RN(n3291), .QN(n155)
         );
  DFFR_X1 \registers_reg[5][4]  ( .D(n3161), .CK(CLK), .RN(n3291), .QN(n156)
         );
  DFFR_X1 \registers_reg[5][3]  ( .D(n3160), .CK(CLK), .RN(n3290), .QN(n157)
         );
  DFFR_X1 \registers_reg[5][2]  ( .D(n3159), .CK(CLK), .RN(n3290), .QN(n158)
         );
  DFFR_X1 \registers_reg[5][1]  ( .D(n3158), .CK(CLK), .RN(n3290), .QN(n159)
         );
  DFFR_X1 \registers_reg[5][0]  ( .D(n3157), .CK(CLK), .RN(n3290), .QN(n160)
         );
  DFFR_X1 \registers_reg[6][31]  ( .D(n3545), .CK(CLK), .RN(n3290), .Q(
        \registers[6][31] ) );
  DFFR_X1 \registers_reg[6][30]  ( .D(n3544), .CK(CLK), .RN(n3290), .Q(
        \registers[6][30] ) );
  DFFR_X1 \registers_reg[6][29]  ( .D(n3543), .CK(CLK), .RN(n3290), .Q(
        \registers[6][29] ) );
  DFFR_X1 \registers_reg[6][28]  ( .D(n3542), .CK(CLK), .RN(n3290), .Q(
        \registers[6][28] ) );
  DFFR_X1 \registers_reg[6][27]  ( .D(n3541), .CK(CLK), .RN(n3290), .Q(
        \registers[6][27] ) );
  DFFR_X1 \registers_reg[6][26]  ( .D(n3540), .CK(CLK), .RN(n3290), .Q(
        \registers[6][26] ) );
  DFFR_X1 \registers_reg[6][25]  ( .D(n3539), .CK(CLK), .RN(n3290), .Q(
        \registers[6][25] ) );
  DFFR_X1 \registers_reg[6][24]  ( .D(n3538), .CK(CLK), .RN(n3289), .Q(
        \registers[6][24] ) );
  DFFR_X1 \registers_reg[6][23]  ( .D(n3537), .CK(CLK), .RN(n3289), .Q(
        \registers[6][23] ) );
  DFFR_X1 \registers_reg[6][22]  ( .D(n3536), .CK(CLK), .RN(n3289), .Q(
        \registers[6][22] ) );
  DFFR_X1 \registers_reg[6][21]  ( .D(n3535), .CK(CLK), .RN(n3289), .Q(
        \registers[6][21] ) );
  DFFR_X1 \registers_reg[6][20]  ( .D(n3534), .CK(CLK), .RN(n3289), .Q(
        \registers[6][20] ) );
  DFFR_X1 \registers_reg[6][19]  ( .D(n3533), .CK(CLK), .RN(n3289), .Q(
        \registers[6][19] ) );
  DFFR_X1 \registers_reg[6][18]  ( .D(n3532), .CK(CLK), .RN(n3289), .Q(
        \registers[6][18] ) );
  DFFR_X1 \registers_reg[6][17]  ( .D(n3531), .CK(CLK), .RN(n3289), .Q(
        \registers[6][17] ) );
  DFFR_X1 \registers_reg[6][16]  ( .D(n3530), .CK(CLK), .RN(n3289), .Q(
        \registers[6][16] ) );
  DFFR_X1 \registers_reg[6][15]  ( .D(n3529), .CK(CLK), .RN(n3289), .Q(
        \registers[6][15] ) );
  DFFR_X1 \registers_reg[6][14]  ( .D(n3528), .CK(CLK), .RN(n3289), .Q(
        \registers[6][14] ) );
  DFFR_X1 \registers_reg[6][13]  ( .D(n3527), .CK(CLK), .RN(n3288), .Q(
        \registers[6][13] ) );
  DFFR_X1 \registers_reg[6][12]  ( .D(n3526), .CK(CLK), .RN(n3288), .Q(
        \registers[6][12] ) );
  DFFR_X1 \registers_reg[6][11]  ( .D(n3525), .CK(CLK), .RN(n3288), .Q(
        \registers[6][11] ) );
  DFFR_X1 \registers_reg[6][10]  ( .D(n3524), .CK(CLK), .RN(n3288), .Q(
        \registers[6][10] ) );
  DFFR_X1 \registers_reg[6][9]  ( .D(n3523), .CK(CLK), .RN(n3288), .Q(
        \registers[6][9] ) );
  DFFR_X1 \registers_reg[6][8]  ( .D(n3522), .CK(CLK), .RN(n3288), .Q(
        \registers[6][8] ) );
  DFFR_X1 \registers_reg[6][7]  ( .D(n3521), .CK(CLK), .RN(n3288), .Q(
        \registers[6][7] ) );
  DFFR_X1 \registers_reg[6][6]  ( .D(n3520), .CK(CLK), .RN(n3288), .Q(
        \registers[6][6] ) );
  DFFR_X1 \registers_reg[6][5]  ( .D(n3519), .CK(CLK), .RN(n3288), .Q(
        \registers[6][5] ) );
  DFFR_X1 \registers_reg[6][4]  ( .D(n3518), .CK(CLK), .RN(n3288), .Q(
        \registers[6][4] ) );
  DFFR_X1 \registers_reg[6][3]  ( .D(n3517), .CK(CLK), .RN(n3288), .Q(
        \registers[6][3] ) );
  DFFR_X1 \registers_reg[6][2]  ( .D(n3516), .CK(CLK), .RN(n3287), .Q(
        \registers[6][2] ) );
  DFFR_X1 \registers_reg[6][1]  ( .D(n3515), .CK(CLK), .RN(n3287), .Q(
        \registers[6][1] ) );
  DFFR_X1 \registers_reg[6][0]  ( .D(n3514), .CK(CLK), .RN(n3287), .Q(
        \registers[6][0] ) );
  DFFR_X1 \registers_reg[7][31]  ( .D(n3458), .CK(CLK), .RN(n3287), .Q(
        \registers[7][31] ) );
  DFFR_X1 \registers_reg[7][30]  ( .D(n3457), .CK(CLK), .RN(n3287), .Q(
        \registers[7][30] ) );
  DFFR_X1 \registers_reg[7][29]  ( .D(n3456), .CK(CLK), .RN(n3287), .Q(
        \registers[7][29] ) );
  DFFR_X1 \registers_reg[7][28]  ( .D(n3455), .CK(CLK), .RN(n3287), .Q(
        \registers[7][28] ) );
  DFFR_X1 \registers_reg[7][27]  ( .D(n3454), .CK(CLK), .RN(n3287), .Q(
        \registers[7][27] ) );
  DFFR_X1 \registers_reg[7][26]  ( .D(n3453), .CK(CLK), .RN(n3287), .Q(
        \registers[7][26] ) );
  DFFR_X1 \registers_reg[7][25]  ( .D(n3452), .CK(CLK), .RN(n3287), .Q(
        \registers[7][25] ) );
  DFFR_X1 \registers_reg[7][24]  ( .D(n3451), .CK(CLK), .RN(n3287), .Q(
        \registers[7][24] ) );
  DFFR_X1 \registers_reg[7][23]  ( .D(n3450), .CK(CLK), .RN(n3286), .Q(
        \registers[7][23] ) );
  DFFR_X1 \registers_reg[7][22]  ( .D(n3481), .CK(CLK), .RN(n3286), .Q(
        \registers[7][22] ) );
  DFFR_X1 \registers_reg[7][21]  ( .D(n3480), .CK(CLK), .RN(n3286), .Q(
        \registers[7][21] ) );
  DFFR_X1 \registers_reg[7][20]  ( .D(n3479), .CK(CLK), .RN(n3286), .Q(
        \registers[7][20] ) );
  DFFR_X1 \registers_reg[7][19]  ( .D(n3478), .CK(CLK), .RN(n3286), .Q(
        \registers[7][19] ) );
  DFFR_X1 \registers_reg[7][18]  ( .D(n3477), .CK(CLK), .RN(n3286), .Q(
        \registers[7][18] ) );
  DFFR_X1 \registers_reg[7][17]  ( .D(n3476), .CK(CLK), .RN(n3286), .Q(
        \registers[7][17] ) );
  DFFR_X1 \registers_reg[7][16]  ( .D(n3475), .CK(CLK), .RN(n3286), .Q(
        \registers[7][16] ) );
  DFFR_X1 \registers_reg[7][15]  ( .D(n3474), .CK(CLK), .RN(n3286), .Q(
        \registers[7][15] ) );
  DFFR_X1 \registers_reg[7][14]  ( .D(n3473), .CK(CLK), .RN(n3286), .Q(
        \registers[7][14] ) );
  DFFR_X1 \registers_reg[7][13]  ( .D(n3472), .CK(CLK), .RN(n3286), .Q(
        \registers[7][13] ) );
  DFFR_X1 \registers_reg[7][12]  ( .D(n3471), .CK(CLK), .RN(n3285), .Q(
        \registers[7][12] ) );
  DFFR_X1 \registers_reg[7][11]  ( .D(n3470), .CK(CLK), .RN(n3285), .Q(
        \registers[7][11] ) );
  DFFR_X1 \registers_reg[7][10]  ( .D(n3469), .CK(CLK), .RN(n3285), .Q(
        \registers[7][10] ) );
  DFFR_X1 \registers_reg[7][9]  ( .D(n3468), .CK(CLK), .RN(n3285), .Q(
        \registers[7][9] ) );
  DFFR_X1 \registers_reg[7][8]  ( .D(n3467), .CK(CLK), .RN(n3285), .Q(
        \registers[7][8] ) );
  DFFR_X1 \registers_reg[7][7]  ( .D(n3466), .CK(CLK), .RN(n3285), .Q(
        \registers[7][7] ) );
  DFFR_X1 \registers_reg[7][6]  ( .D(n3465), .CK(CLK), .RN(n3285), .Q(
        \registers[7][6] ) );
  DFFR_X1 \registers_reg[7][5]  ( .D(n3464), .CK(CLK), .RN(n3285), .Q(
        \registers[7][5] ) );
  DFFR_X1 \registers_reg[7][4]  ( .D(n3463), .CK(CLK), .RN(n3285), .Q(
        \registers[7][4] ) );
  DFFR_X1 \registers_reg[7][3]  ( .D(n3462), .CK(CLK), .RN(n3285), .Q(
        \registers[7][3] ) );
  DFFR_X1 \registers_reg[7][2]  ( .D(n3461), .CK(CLK), .RN(n3285), .Q(
        \registers[7][2] ) );
  DFFR_X1 \registers_reg[7][1]  ( .D(n3460), .CK(CLK), .RN(n1501), .Q(
        \registers[7][1] ) );
  DFFR_X1 \registers_reg[7][0]  ( .D(n3459), .CK(CLK), .RN(n1501), .Q(
        \registers[7][0] ) );
  DFFR_X1 \registers_reg[8][31]  ( .D(n3353), .CK(CLK), .RN(n1501), .Q(
        \registers[8][31] ) );
  DFFR_X1 \registers_reg[8][30]  ( .D(n3352), .CK(CLK), .RN(n1501), .Q(
        \registers[8][30] ) );
  DFFR_X1 \registers_reg[8][29]  ( .D(n3351), .CK(CLK), .RN(n1501), .Q(
        \registers[8][29] ) );
  DFFR_X1 \registers_reg[8][28]  ( .D(n3350), .CK(CLK), .RN(n1501), .Q(
        \registers[8][28] ) );
  DFFR_X1 \registers_reg[8][27]  ( .D(n3349), .CK(CLK), .RN(n1501), .Q(
        \registers[8][27] ) );
  DFFR_X1 \registers_reg[8][26]  ( .D(n3348), .CK(CLK), .RN(n1501), .Q(
        \registers[8][26] ) );
  DFFR_X1 \registers_reg[8][25]  ( .D(n3347), .CK(CLK), .RN(n1501), .Q(
        \registers[8][25] ) );
  DFFR_X1 \registers_reg[8][24]  ( .D(n3346), .CK(CLK), .RN(n1501), .Q(
        \registers[8][24] ) );
  DFFR_X1 \registers_reg[8][23]  ( .D(n3345), .CK(CLK), .RN(n1501), .Q(
        \registers[8][23] ) );
  DFFR_X1 \registers_reg[8][22]  ( .D(n3344), .CK(CLK), .RN(n1500), .Q(
        \registers[8][22] ) );
  DFFR_X1 \registers_reg[8][21]  ( .D(n3343), .CK(CLK), .RN(n1500), .Q(
        \registers[8][21] ) );
  DFFR_X1 \registers_reg[8][20]  ( .D(n3342), .CK(CLK), .RN(n1500), .Q(
        \registers[8][20] ) );
  DFFR_X1 \registers_reg[8][19]  ( .D(n3341), .CK(CLK), .RN(n1500), .Q(
        \registers[8][19] ) );
  DFFR_X1 \registers_reg[8][18]  ( .D(n3340), .CK(CLK), .RN(n1500), .Q(
        \registers[8][18] ) );
  DFFR_X1 \registers_reg[8][17]  ( .D(n3339), .CK(CLK), .RN(n1500), .Q(
        \registers[8][17] ) );
  DFFR_X1 \registers_reg[8][16]  ( .D(n3338), .CK(CLK), .RN(n1500), .Q(
        \registers[8][16] ) );
  DFFR_X1 \registers_reg[8][15]  ( .D(n3337), .CK(CLK), .RN(n1500), .Q(
        \registers[8][15] ) );
  DFFR_X1 \registers_reg[8][14]  ( .D(n3336), .CK(CLK), .RN(n1500), .Q(
        \registers[8][14] ) );
  DFFR_X1 \registers_reg[8][13]  ( .D(n3335), .CK(CLK), .RN(n1500), .Q(
        \registers[8][13] ) );
  DFFR_X1 \registers_reg[8][12]  ( .D(n3334), .CK(CLK), .RN(n1500), .Q(
        \registers[8][12] ) );
  DFFR_X1 \registers_reg[8][11]  ( .D(n3333), .CK(CLK), .RN(n1433), .Q(
        \registers[8][11] ) );
  DFFR_X1 \registers_reg[8][10]  ( .D(n3332), .CK(CLK), .RN(n1433), .Q(
        \registers[8][10] ) );
  DFFR_X1 \registers_reg[8][9]  ( .D(n3331), .CK(CLK), .RN(n1433), .Q(
        \registers[8][9] ) );
  DFFR_X1 \registers_reg[8][8]  ( .D(n3330), .CK(CLK), .RN(n1433), .Q(
        \registers[8][8] ) );
  DFFR_X1 \registers_reg[8][7]  ( .D(n3329), .CK(CLK), .RN(n1433), .Q(
        \registers[8][7] ) );
  DFFR_X1 \registers_reg[8][6]  ( .D(n3328), .CK(CLK), .RN(n1433), .Q(
        \registers[8][6] ) );
  DFFR_X1 \registers_reg[8][5]  ( .D(n3327), .CK(CLK), .RN(n1433), .Q(
        \registers[8][5] ) );
  DFFR_X1 \registers_reg[8][4]  ( .D(n3326), .CK(CLK), .RN(n1433), .Q(
        \registers[8][4] ) );
  DFFR_X1 \registers_reg[8][3]  ( .D(n3325), .CK(CLK), .RN(n1433), .Q(
        \registers[8][3] ) );
  DFFR_X1 \registers_reg[8][2]  ( .D(n3324), .CK(CLK), .RN(n1433), .Q(
        \registers[8][2] ) );
  DFFR_X1 \registers_reg[8][1]  ( .D(n3323), .CK(CLK), .RN(n1433), .Q(
        \registers[8][1] ) );
  DFFR_X1 \registers_reg[8][0]  ( .D(n3322), .CK(CLK), .RN(n1431), .Q(
        \registers[8][0] ) );
  DFFR_X1 \registers_reg[9][31]  ( .D(n3385), .CK(CLK), .RN(n1431), .Q(
        \registers[9][31] ) );
  DFFR_X1 \registers_reg[9][30]  ( .D(n3384), .CK(CLK), .RN(n1431), .Q(
        \registers[9][30] ) );
  DFFR_X1 \registers_reg[9][29]  ( .D(n3383), .CK(CLK), .RN(n1431), .Q(
        \registers[9][29] ) );
  DFFR_X1 \registers_reg[9][28]  ( .D(n3382), .CK(CLK), .RN(n1431), .Q(
        \registers[9][28] ) );
  DFFR_X1 \registers_reg[9][27]  ( .D(n3381), .CK(CLK), .RN(n1431), .Q(
        \registers[9][27] ) );
  DFFR_X1 \registers_reg[9][26]  ( .D(n3380), .CK(CLK), .RN(n1431), .Q(
        \registers[9][26] ) );
  DFFR_X1 \registers_reg[9][25]  ( .D(n3379), .CK(CLK), .RN(n1431), .Q(
        \registers[9][25] ) );
  DFFR_X1 \registers_reg[9][24]  ( .D(n3378), .CK(CLK), .RN(n1431), .Q(
        \registers[9][24] ) );
  DFFR_X1 \registers_reg[9][23]  ( .D(n3377), .CK(CLK), .RN(n1431), .Q(
        \registers[9][23] ) );
  DFFR_X1 \registers_reg[9][22]  ( .D(n3376), .CK(CLK), .RN(n1431), .Q(
        \registers[9][22] ) );
  DFFR_X1 \registers_reg[9][21]  ( .D(n3375), .CK(CLK), .RN(n1430), .Q(
        \registers[9][21] ) );
  DFFR_X1 \registers_reg[9][20]  ( .D(n3374), .CK(CLK), .RN(n1430), .Q(
        \registers[9][20] ) );
  DFFR_X1 \registers_reg[9][19]  ( .D(n3373), .CK(CLK), .RN(n1430), .Q(
        \registers[9][19] ) );
  DFFR_X1 \registers_reg[9][18]  ( .D(n3372), .CK(CLK), .RN(n1430), .Q(
        \registers[9][18] ) );
  DFFR_X1 \registers_reg[9][17]  ( .D(n3371), .CK(CLK), .RN(n1430), .Q(
        \registers[9][17] ) );
  DFFR_X1 \registers_reg[9][16]  ( .D(n3370), .CK(CLK), .RN(n1430), .Q(
        \registers[9][16] ) );
  DFFR_X1 \registers_reg[9][15]  ( .D(n3369), .CK(CLK), .RN(n1430), .Q(
        \registers[9][15] ) );
  DFFR_X1 \registers_reg[9][14]  ( .D(n3368), .CK(CLK), .RN(n1430), .Q(
        \registers[9][14] ) );
  DFFR_X1 \registers_reg[9][13]  ( .D(n3367), .CK(CLK), .RN(n1430), .Q(
        \registers[9][13] ) );
  DFFR_X1 \registers_reg[9][12]  ( .D(n3366), .CK(CLK), .RN(n1430), .Q(
        \registers[9][12] ) );
  DFFR_X1 \registers_reg[9][11]  ( .D(n3365), .CK(CLK), .RN(n1430), .Q(
        \registers[9][11] ) );
  DFFR_X1 \registers_reg[9][10]  ( .D(n3364), .CK(CLK), .RN(n1429), .Q(
        \registers[9][10] ) );
  DFFR_X1 \registers_reg[9][9]  ( .D(n3363), .CK(CLK), .RN(n1429), .Q(
        \registers[9][9] ) );
  DFFR_X1 \registers_reg[9][8]  ( .D(n3362), .CK(CLK), .RN(n1429), .Q(
        \registers[9][8] ) );
  DFFR_X1 \registers_reg[9][7]  ( .D(n3361), .CK(CLK), .RN(n1429), .Q(
        \registers[9][7] ) );
  DFFR_X1 \registers_reg[9][6]  ( .D(n3360), .CK(CLK), .RN(n1429), .Q(
        \registers[9][6] ) );
  DFFR_X1 \registers_reg[9][5]  ( .D(n3359), .CK(CLK), .RN(n1429), .Q(
        \registers[9][5] ) );
  DFFR_X1 \registers_reg[9][4]  ( .D(n3358), .CK(CLK), .RN(n1429), .Q(
        \registers[9][4] ) );
  DFFR_X1 \registers_reg[9][3]  ( .D(n3357), .CK(CLK), .RN(n1429), .Q(
        \registers[9][3] ) );
  DFFR_X1 \registers_reg[9][2]  ( .D(n3356), .CK(CLK), .RN(n1429), .Q(
        \registers[9][2] ) );
  DFFR_X1 \registers_reg[9][1]  ( .D(n3355), .CK(CLK), .RN(n1429), .Q(
        \registers[9][1] ) );
  DFFR_X1 \registers_reg[9][0]  ( .D(n3354), .CK(CLK), .RN(n1429), .Q(
        \registers[9][0] ) );
  DFFR_X1 \registers_reg[10][31]  ( .D(n3156), .CK(CLK), .RN(n1362), .QN(n289)
         );
  DFFR_X1 \registers_reg[10][30]  ( .D(n3155), .CK(CLK), .RN(n1362), .QN(n290)
         );
  DFFR_X1 \registers_reg[10][29]  ( .D(n3154), .CK(CLK), .RN(n1362), .QN(n291)
         );
  DFFR_X1 \registers_reg[10][28]  ( .D(n3153), .CK(CLK), .RN(n1362), .QN(n292)
         );
  DFFR_X1 \registers_reg[10][27]  ( .D(n3152), .CK(CLK), .RN(n1362), .QN(n293)
         );
  DFFR_X1 \registers_reg[10][26]  ( .D(n3151), .CK(CLK), .RN(n1362), .QN(n294)
         );
  DFFR_X1 \registers_reg[10][25]  ( .D(n3150), .CK(CLK), .RN(n1362), .QN(n295)
         );
  DFFR_X1 \registers_reg[10][24]  ( .D(n3149), .CK(CLK), .RN(n1362), .QN(n296)
         );
  DFFR_X1 \registers_reg[10][23]  ( .D(n3148), .CK(CLK), .RN(n1362), .QN(n297)
         );
  DFFR_X1 \registers_reg[10][22]  ( .D(n3147), .CK(CLK), .RN(n1362), .QN(n298)
         );
  DFFR_X1 \registers_reg[10][21]  ( .D(n3146), .CK(CLK), .RN(n1362), .QN(n299)
         );
  DFFR_X1 \registers_reg[10][20]  ( .D(n3145), .CK(CLK), .RN(n1361), .QN(n300)
         );
  DFFR_X1 \registers_reg[10][19]  ( .D(n3144), .CK(CLK), .RN(n1361), .QN(n301)
         );
  DFFR_X1 \registers_reg[10][18]  ( .D(n3143), .CK(CLK), .RN(n1361), .QN(n302)
         );
  DFFR_X1 \registers_reg[10][17]  ( .D(n3142), .CK(CLK), .RN(n1361), .QN(n303)
         );
  DFFR_X1 \registers_reg[10][16]  ( .D(n3141), .CK(CLK), .RN(n1361), .QN(n304)
         );
  DFFR_X1 \registers_reg[10][15]  ( .D(n3140), .CK(CLK), .RN(n1361), .QN(n305)
         );
  DFFR_X1 \registers_reg[10][14]  ( .D(n3139), .CK(CLK), .RN(n1361), .QN(n306)
         );
  DFFR_X1 \registers_reg[10][13]  ( .D(n3138), .CK(CLK), .RN(n1361), .QN(n307)
         );
  DFFR_X1 \registers_reg[10][12]  ( .D(n3137), .CK(CLK), .RN(n1361), .QN(n308)
         );
  DFFR_X1 \registers_reg[10][11]  ( .D(n3136), .CK(CLK), .RN(n1361), .QN(n309)
         );
  DFFR_X1 \registers_reg[10][10]  ( .D(n3135), .CK(CLK), .RN(n1361), .QN(n310)
         );
  DFFR_X1 \registers_reg[10][9]  ( .D(n3134), .CK(CLK), .RN(n1226), .QN(n311)
         );
  DFFR_X1 \registers_reg[10][8]  ( .D(n3133), .CK(CLK), .RN(n1226), .QN(n312)
         );
  DFFR_X1 \registers_reg[10][7]  ( .D(n3132), .CK(CLK), .RN(n1226), .QN(n313)
         );
  DFFR_X1 \registers_reg[10][6]  ( .D(n3131), .CK(CLK), .RN(n1226), .QN(n314)
         );
  DFFR_X1 \registers_reg[10][5]  ( .D(n3130), .CK(CLK), .RN(n1226), .QN(n315)
         );
  DFFR_X1 \registers_reg[10][4]  ( .D(n3129), .CK(CLK), .RN(n1226), .QN(n316)
         );
  DFFR_X1 \registers_reg[10][3]  ( .D(n3128), .CK(CLK), .RN(n1226), .QN(n317)
         );
  DFFR_X1 \registers_reg[10][2]  ( .D(n3127), .CK(CLK), .RN(n1226), .QN(n318)
         );
  DFFR_X1 \registers_reg[10][1]  ( .D(n3126), .CK(CLK), .RN(n1226), .QN(n319)
         );
  DFFR_X1 \registers_reg[10][0]  ( .D(n3125), .CK(CLK), .RN(n1226), .QN(n320)
         );
  DFFR_X1 \registers_reg[11][31]  ( .D(n3124), .CK(CLK), .RN(n1226), .QN(n321)
         );
  DFFR_X1 \registers_reg[11][30]  ( .D(n3123), .CK(CLK), .RN(n1225), .QN(n322)
         );
  DFFR_X1 \registers_reg[11][29]  ( .D(n3122), .CK(CLK), .RN(n1225), .QN(n323)
         );
  DFFR_X1 \registers_reg[11][28]  ( .D(n3121), .CK(CLK), .RN(n1225), .QN(n324)
         );
  DFFR_X1 \registers_reg[11][27]  ( .D(n3120), .CK(CLK), .RN(n1225), .QN(n325)
         );
  DFFR_X1 \registers_reg[11][26]  ( .D(n3119), .CK(CLK), .RN(n1225), .QN(n326)
         );
  DFFR_X1 \registers_reg[11][25]  ( .D(n3118), .CK(CLK), .RN(n1225), .QN(n327)
         );
  DFFR_X1 \registers_reg[11][24]  ( .D(n3117), .CK(CLK), .RN(n1225), .QN(n328)
         );
  DFFR_X1 \registers_reg[11][23]  ( .D(n3116), .CK(CLK), .RN(n1225), .QN(n329)
         );
  DFFR_X1 \registers_reg[11][22]  ( .D(n3115), .CK(CLK), .RN(n1225), .QN(n330)
         );
  DFFR_X1 \registers_reg[11][21]  ( .D(n3114), .CK(CLK), .RN(n1225), .QN(n331)
         );
  DFFR_X1 \registers_reg[11][20]  ( .D(n3113), .CK(CLK), .RN(n1225), .QN(n332)
         );
  DFFR_X1 \registers_reg[11][19]  ( .D(n3112), .CK(CLK), .RN(n1158), .QN(n333)
         );
  DFFR_X1 \registers_reg[11][18]  ( .D(n3111), .CK(CLK), .RN(n1158), .QN(n334)
         );
  DFFR_X1 \registers_reg[11][17]  ( .D(n3110), .CK(CLK), .RN(n1158), .QN(n335)
         );
  DFFR_X1 \registers_reg[11][16]  ( .D(n3109), .CK(CLK), .RN(n1158), .QN(n336)
         );
  DFFR_X1 \registers_reg[11][15]  ( .D(n3108), .CK(CLK), .RN(n1158), .QN(n337)
         );
  DFFR_X1 \registers_reg[11][14]  ( .D(n3107), .CK(CLK), .RN(n1158), .QN(n338)
         );
  DFFR_X1 \registers_reg[11][13]  ( .D(n3106), .CK(CLK), .RN(n1158), .QN(n339)
         );
  DFFR_X1 \registers_reg[11][12]  ( .D(n3105), .CK(CLK), .RN(n1158), .QN(n340)
         );
  DFFR_X1 \registers_reg[11][11]  ( .D(n3104), .CK(CLK), .RN(n1158), .QN(n341)
         );
  DFFR_X1 \registers_reg[11][10]  ( .D(n3103), .CK(CLK), .RN(n1158), .QN(n342)
         );
  DFFR_X1 \registers_reg[11][9]  ( .D(n3102), .CK(CLK), .RN(n1158), .QN(n343)
         );
  DFFR_X1 \registers_reg[11][8]  ( .D(n3101), .CK(CLK), .RN(n1155), .QN(n344)
         );
  DFFR_X1 \registers_reg[11][7]  ( .D(n3100), .CK(CLK), .RN(n1155), .QN(n345)
         );
  DFFR_X1 \registers_reg[11][6]  ( .D(n3099), .CK(CLK), .RN(n1155), .QN(n346)
         );
  DFFR_X1 \registers_reg[11][5]  ( .D(n3098), .CK(CLK), .RN(n1155), .QN(n347)
         );
  DFFR_X1 \registers_reg[11][4]  ( .D(n3097), .CK(CLK), .RN(n1155), .QN(n348)
         );
  DFFR_X1 \registers_reg[11][3]  ( .D(n3096), .CK(CLK), .RN(n1155), .QN(n349)
         );
  DFFR_X1 \registers_reg[11][2]  ( .D(n3095), .CK(CLK), .RN(n1155), .QN(n350)
         );
  DFFR_X1 \registers_reg[11][1]  ( .D(n3094), .CK(CLK), .RN(n1155), .QN(n351)
         );
  DFFR_X1 \registers_reg[11][0]  ( .D(n3093), .CK(CLK), .RN(n1155), .QN(n352)
         );
  DFFR_X1 \registers_reg[12][31]  ( .D(n3417), .CK(CLK), .RN(n1155), .Q(
        \registers[12][31] ) );
  DFFR_X1 \registers_reg[12][30]  ( .D(n3416), .CK(CLK), .RN(n1155), .Q(
        \registers[12][30] ) );
  DFFR_X1 \registers_reg[12][29]  ( .D(n3415), .CK(CLK), .RN(n1118), .Q(
        \registers[12][29] ) );
  DFFR_X1 \registers_reg[12][28]  ( .D(n3414), .CK(CLK), .RN(n1118), .Q(
        \registers[12][28] ) );
  DFFR_X1 \registers_reg[12][27]  ( .D(n3413), .CK(CLK), .RN(n1118), .Q(
        \registers[12][27] ) );
  DFFR_X1 \registers_reg[12][26]  ( .D(n3412), .CK(CLK), .RN(n1118), .Q(
        \registers[12][26] ) );
  DFFR_X1 \registers_reg[12][25]  ( .D(n3411), .CK(CLK), .RN(n1118), .Q(
        \registers[12][25] ) );
  DFFR_X1 \registers_reg[12][24]  ( .D(n3410), .CK(CLK), .RN(n1118), .Q(
        \registers[12][24] ) );
  DFFR_X1 \registers_reg[12][23]  ( .D(n3409), .CK(CLK), .RN(n1118), .Q(
        \registers[12][23] ) );
  DFFR_X1 \registers_reg[12][22]  ( .D(n3408), .CK(CLK), .RN(n1118), .Q(
        \registers[12][22] ) );
  DFFR_X1 \registers_reg[12][21]  ( .D(n3407), .CK(CLK), .RN(n1118), .Q(
        \registers[12][21] ) );
  DFFR_X1 \registers_reg[12][20]  ( .D(n3406), .CK(CLK), .RN(n1118), .Q(
        \registers[12][20] ) );
  DFFR_X1 \registers_reg[12][19]  ( .D(n3405), .CK(CLK), .RN(n1118), .Q(
        \registers[12][19] ) );
  DFFR_X1 \registers_reg[12][18]  ( .D(n3404), .CK(CLK), .RN(n1116), .Q(
        \registers[12][18] ) );
  DFFR_X1 \registers_reg[12][17]  ( .D(n3403), .CK(CLK), .RN(n1116), .Q(
        \registers[12][17] ) );
  DFFR_X1 \registers_reg[12][16]  ( .D(n3402), .CK(CLK), .RN(n1116), .Q(
        \registers[12][16] ) );
  DFFR_X1 \registers_reg[12][15]  ( .D(n3401), .CK(CLK), .RN(n1116), .Q(
        \registers[12][15] ) );
  DFFR_X1 \registers_reg[12][14]  ( .D(n3400), .CK(CLK), .RN(n1116), .Q(
        \registers[12][14] ) );
  DFFR_X1 \registers_reg[12][13]  ( .D(n3399), .CK(CLK), .RN(n1116), .Q(
        \registers[12][13] ) );
  DFFR_X1 \registers_reg[12][12]  ( .D(n3398), .CK(CLK), .RN(n1116), .Q(
        \registers[12][12] ) );
  DFFR_X1 \registers_reg[12][11]  ( .D(n3397), .CK(CLK), .RN(n1116), .Q(
        \registers[12][11] ) );
  DFFR_X1 \registers_reg[12][10]  ( .D(n3396), .CK(CLK), .RN(n1116), .Q(
        \registers[12][10] ) );
  DFFR_X1 \registers_reg[12][9]  ( .D(n3395), .CK(CLK), .RN(n1116), .Q(
        \registers[12][9] ) );
  DFFR_X1 \registers_reg[12][8]  ( .D(n3394), .CK(CLK), .RN(n1116), .Q(
        \registers[12][8] ) );
  DFFR_X1 \registers_reg[12][7]  ( .D(n3393), .CK(CLK), .RN(n1114), .Q(
        \registers[12][7] ) );
  DFFR_X1 \registers_reg[12][6]  ( .D(n3392), .CK(CLK), .RN(n1114), .Q(
        \registers[12][6] ) );
  DFFR_X1 \registers_reg[12][5]  ( .D(n3391), .CK(CLK), .RN(n1114), .Q(
        \registers[12][5] ) );
  DFFR_X1 \registers_reg[12][4]  ( .D(n3390), .CK(CLK), .RN(n1114), .Q(
        \registers[12][4] ) );
  DFFR_X1 \registers_reg[12][3]  ( .D(n3389), .CK(CLK), .RN(n1114), .Q(
        \registers[12][3] ) );
  DFFR_X1 \registers_reg[12][2]  ( .D(n3388), .CK(CLK), .RN(n1114), .Q(
        \registers[12][2] ) );
  DFFR_X1 \registers_reg[12][1]  ( .D(n3387), .CK(CLK), .RN(n1114), .Q(
        \registers[12][1] ) );
  DFFR_X1 \registers_reg[12][0]  ( .D(n3386), .CK(CLK), .RN(n1114), .Q(
        \registers[12][0] ) );
  DFFR_X1 \registers_reg[13][31]  ( .D(n3449), .CK(CLK), .RN(n1114), .Q(
        \registers[13][31] ) );
  DFFR_X1 \registers_reg[13][30]  ( .D(n3448), .CK(CLK), .RN(n1114), .Q(
        \registers[13][30] ) );
  DFFR_X1 \registers_reg[13][29]  ( .D(n3447), .CK(CLK), .RN(n1114), .Q(
        \registers[13][29] ) );
  DFFR_X1 \registers_reg[13][28]  ( .D(n3446), .CK(CLK), .RN(n1112), .Q(
        \registers[13][28] ) );
  DFFR_X1 \registers_reg[13][27]  ( .D(n3445), .CK(CLK), .RN(n1112), .Q(
        \registers[13][27] ) );
  DFFR_X1 \registers_reg[13][26]  ( .D(n3444), .CK(CLK), .RN(n1112), .Q(
        \registers[13][26] ) );
  DFFR_X1 \registers_reg[13][25]  ( .D(n3443), .CK(CLK), .RN(n1112), .Q(
        \registers[13][25] ) );
  DFFR_X1 \registers_reg[13][24]  ( .D(n3442), .CK(CLK), .RN(n1112), .Q(
        \registers[13][24] ) );
  DFFR_X1 \registers_reg[13][23]  ( .D(n3441), .CK(CLK), .RN(n1112), .Q(
        \registers[13][23] ) );
  DFFR_X1 \registers_reg[13][22]  ( .D(n3440), .CK(CLK), .RN(n1112), .Q(
        \registers[13][22] ) );
  DFFR_X1 \registers_reg[13][21]  ( .D(n3439), .CK(CLK), .RN(n1112), .Q(
        \registers[13][21] ) );
  DFFR_X1 \registers_reg[13][20]  ( .D(n3438), .CK(CLK), .RN(n1112), .Q(
        \registers[13][20] ) );
  DFFR_X1 \registers_reg[13][19]  ( .D(n3437), .CK(CLK), .RN(n1112), .Q(
        \registers[13][19] ) );
  DFFR_X1 \registers_reg[13][18]  ( .D(n3436), .CK(CLK), .RN(n1112), .Q(
        \registers[13][18] ) );
  DFFR_X1 \registers_reg[13][17]  ( .D(n3435), .CK(CLK), .RN(n1066), .Q(
        \registers[13][17] ) );
  DFFR_X1 \registers_reg[13][16]  ( .D(n3434), .CK(CLK), .RN(n1066), .Q(
        \registers[13][16] ) );
  DFFR_X1 \registers_reg[13][15]  ( .D(n3433), .CK(CLK), .RN(n1066), .Q(
        \registers[13][15] ) );
  DFFR_X1 \registers_reg[13][14]  ( .D(n3432), .CK(CLK), .RN(n1066), .Q(
        \registers[13][14] ) );
  DFFR_X1 \registers_reg[13][13]  ( .D(n3431), .CK(CLK), .RN(n1066), .Q(
        \registers[13][13] ) );
  DFFR_X1 \registers_reg[13][12]  ( .D(n3430), .CK(CLK), .RN(n1066), .Q(
        \registers[13][12] ) );
  DFFR_X1 \registers_reg[13][11]  ( .D(n3429), .CK(CLK), .RN(n1066), .Q(
        \registers[13][11] ) );
  DFFR_X1 \registers_reg[13][10]  ( .D(n3428), .CK(CLK), .RN(n1066), .Q(
        \registers[13][10] ) );
  DFFR_X1 \registers_reg[13][9]  ( .D(n3427), .CK(CLK), .RN(n1066), .Q(
        \registers[13][9] ) );
  DFFR_X1 \registers_reg[13][8]  ( .D(n3426), .CK(CLK), .RN(n1066), .Q(
        \registers[13][8] ) );
  DFFR_X1 \registers_reg[13][7]  ( .D(n3425), .CK(CLK), .RN(n1066), .Q(
        \registers[13][7] ) );
  DFFR_X1 \registers_reg[13][6]  ( .D(n3424), .CK(CLK), .RN(n1065), .Q(
        \registers[13][6] ) );
  DFFR_X1 \registers_reg[13][5]  ( .D(n3423), .CK(CLK), .RN(n1065), .Q(
        \registers[13][5] ) );
  DFFR_X1 \registers_reg[13][4]  ( .D(n3422), .CK(CLK), .RN(n1065), .Q(
        \registers[13][4] ) );
  DFFR_X1 \registers_reg[13][3]  ( .D(n3421), .CK(CLK), .RN(n1065), .Q(
        \registers[13][3] ) );
  DFFR_X1 \registers_reg[13][2]  ( .D(n3420), .CK(CLK), .RN(n1065), .Q(
        \registers[13][2] ) );
  DFFR_X1 \registers_reg[13][1]  ( .D(n3419), .CK(CLK), .RN(n1065), .Q(
        \registers[13][1] ) );
  DFFR_X1 \registers_reg[13][0]  ( .D(n3418), .CK(CLK), .RN(n1065), .Q(
        \registers[13][0] ) );
  DFFR_X1 \registers_reg[14][31]  ( .D(n3092), .CK(CLK), .RN(n1065), .QN(n417)
         );
  DFFR_X1 \registers_reg[14][30]  ( .D(n3091), .CK(CLK), .RN(n1065), .QN(n418)
         );
  DFFR_X1 \registers_reg[14][29]  ( .D(n3090), .CK(CLK), .RN(n1065), .QN(n419)
         );
  DFFR_X1 \registers_reg[14][28]  ( .D(n3089), .CK(CLK), .RN(n1065), .QN(n420)
         );
  DFFR_X1 \registers_reg[14][27]  ( .D(n3088), .CK(CLK), .RN(n1064), .QN(n421)
         );
  DFFR_X1 \registers_reg[14][26]  ( .D(n3087), .CK(CLK), .RN(n1064), .QN(n422)
         );
  DFFR_X1 \registers_reg[14][25]  ( .D(n3086), .CK(CLK), .RN(n1064), .QN(n423)
         );
  DFFR_X1 \registers_reg[14][24]  ( .D(n3085), .CK(CLK), .RN(n1064), .QN(n424)
         );
  DFFR_X1 \registers_reg[14][23]  ( .D(n3084), .CK(CLK), .RN(n1064), .QN(n425)
         );
  DFFR_X1 \registers_reg[14][22]  ( .D(n3083), .CK(CLK), .RN(n1064), .QN(n426)
         );
  DFFR_X1 \registers_reg[14][21]  ( .D(n3082), .CK(CLK), .RN(n1064), .QN(n427)
         );
  DFFR_X1 \registers_reg[14][20]  ( .D(n3081), .CK(CLK), .RN(n1064), .QN(n428)
         );
  DFFR_X1 \registers_reg[14][19]  ( .D(n3080), .CK(CLK), .RN(n1064), .QN(n429)
         );
  DFFR_X1 \registers_reg[14][18]  ( .D(n3079), .CK(CLK), .RN(n1064), .QN(n430)
         );
  DFFR_X1 \registers_reg[14][17]  ( .D(n3078), .CK(CLK), .RN(n1064), .QN(n431)
         );
  DFFR_X1 \registers_reg[14][16]  ( .D(n3077), .CK(CLK), .RN(n1063), .QN(n432)
         );
  DFFR_X1 \registers_reg[14][15]  ( .D(n3076), .CK(CLK), .RN(n1063), .QN(n433)
         );
  DFFR_X1 \registers_reg[14][14]  ( .D(n3075), .CK(CLK), .RN(n1063), .QN(n434)
         );
  DFFR_X1 \registers_reg[14][13]  ( .D(n3074), .CK(CLK), .RN(n1063), .QN(n435)
         );
  DFFR_X1 \registers_reg[14][12]  ( .D(n3073), .CK(CLK), .RN(n1063), .QN(n436)
         );
  DFFR_X1 \registers_reg[14][11]  ( .D(n3072), .CK(CLK), .RN(n1063), .QN(n437)
         );
  DFFR_X1 \registers_reg[14][10]  ( .D(n3071), .CK(CLK), .RN(n1063), .QN(n438)
         );
  DFFR_X1 \registers_reg[14][9]  ( .D(n3070), .CK(CLK), .RN(n1063), .QN(n439)
         );
  DFFR_X1 \registers_reg[14][8]  ( .D(n3069), .CK(CLK), .RN(n1063), .QN(n440)
         );
  DFFR_X1 \registers_reg[14][7]  ( .D(n3068), .CK(CLK), .RN(n1063), .QN(n441)
         );
  DFFR_X1 \registers_reg[14][6]  ( .D(n3067), .CK(CLK), .RN(n1063), .QN(n442)
         );
  DFFR_X1 \registers_reg[14][5]  ( .D(n3066), .CK(CLK), .RN(n1062), .QN(n443)
         );
  DFFR_X1 \registers_reg[14][4]  ( .D(n3065), .CK(CLK), .RN(n1062), .QN(n444)
         );
  DFFR_X1 \registers_reg[14][3]  ( .D(n3064), .CK(CLK), .RN(n1062), .QN(n445)
         );
  DFFR_X1 \registers_reg[14][2]  ( .D(n3063), .CK(CLK), .RN(n1062), .QN(n446)
         );
  DFFR_X1 \registers_reg[14][1]  ( .D(n3062), .CK(CLK), .RN(n1062), .QN(n447)
         );
  DFFR_X1 \registers_reg[14][0]  ( .D(n3061), .CK(CLK), .RN(n1062), .QN(n448)
         );
  DFFR_X1 \registers_reg[15][31]  ( .D(n3060), .CK(CLK), .RN(n1062), .QN(n449)
         );
  DFFR_X1 \registers_reg[15][30]  ( .D(n3059), .CK(CLK), .RN(n1062), .QN(n450)
         );
  DFFR_X1 \registers_reg[15][29]  ( .D(n3058), .CK(CLK), .RN(n1062), .QN(n451)
         );
  DFFR_X1 \registers_reg[15][28]  ( .D(n3057), .CK(CLK), .RN(n1062), .QN(n452)
         );
  DFFR_X1 \registers_reg[15][27]  ( .D(n3056), .CK(CLK), .RN(n1062), .QN(n453)
         );
  DFFR_X1 \registers_reg[15][26]  ( .D(n3055), .CK(CLK), .RN(n1061), .QN(n454)
         );
  DFFR_X1 \registers_reg[15][25]  ( .D(n3054), .CK(CLK), .RN(n1061), .QN(n455)
         );
  DFFR_X1 \registers_reg[15][24]  ( .D(n3053), .CK(CLK), .RN(n1061), .QN(n456)
         );
  DFFR_X1 \registers_reg[15][23]  ( .D(n3052), .CK(CLK), .RN(n1061), .QN(n457)
         );
  DFFR_X1 \registers_reg[15][22]  ( .D(n3051), .CK(CLK), .RN(n1061), .QN(n458)
         );
  DFFR_X1 \registers_reg[15][21]  ( .D(n3050), .CK(CLK), .RN(n1061), .QN(n459)
         );
  DFFR_X1 \registers_reg[15][20]  ( .D(n3049), .CK(CLK), .RN(n1061), .QN(n460)
         );
  DFFR_X1 \registers_reg[15][19]  ( .D(n3048), .CK(CLK), .RN(n1061), .QN(n461)
         );
  DFFR_X1 \registers_reg[15][18]  ( .D(n3047), .CK(CLK), .RN(n1061), .QN(n462)
         );
  DFFR_X1 \registers_reg[15][17]  ( .D(n3046), .CK(CLK), .RN(n1061), .QN(n463)
         );
  DFFR_X1 \registers_reg[15][16]  ( .D(n3045), .CK(CLK), .RN(n1061), .QN(n464)
         );
  DFFR_X1 \registers_reg[15][15]  ( .D(n3044), .CK(CLK), .RN(n1060), .QN(n465)
         );
  DFFR_X1 \registers_reg[15][14]  ( .D(n3043), .CK(CLK), .RN(n1060), .QN(n466)
         );
  DFFR_X1 \registers_reg[15][13]  ( .D(n3042), .CK(CLK), .RN(n1060), .QN(n467)
         );
  DFFR_X1 \registers_reg[15][12]  ( .D(n3041), .CK(CLK), .RN(n1060), .QN(n468)
         );
  DFFR_X1 \registers_reg[15][11]  ( .D(n3040), .CK(CLK), .RN(n1060), .QN(n469)
         );
  DFFR_X1 \registers_reg[15][10]  ( .D(n3039), .CK(CLK), .RN(n1060), .QN(n470)
         );
  DFFR_X1 \registers_reg[15][9]  ( .D(n3038), .CK(CLK), .RN(n1060), .QN(n471)
         );
  DFFR_X1 \registers_reg[15][8]  ( .D(n3037), .CK(CLK), .RN(n1060), .QN(n472)
         );
  DFFR_X1 \registers_reg[15][7]  ( .D(n3036), .CK(CLK), .RN(n1060), .QN(n473)
         );
  DFFR_X1 \registers_reg[15][6]  ( .D(n3035), .CK(CLK), .RN(n1060), .QN(n474)
         );
  DFFR_X1 \registers_reg[15][5]  ( .D(n3034), .CK(CLK), .RN(n1060), .QN(n475)
         );
  DFFR_X1 \registers_reg[15][4]  ( .D(n3033), .CK(CLK), .RN(n1059), .QN(n476)
         );
  DFFR_X1 \registers_reg[15][3]  ( .D(n3032), .CK(CLK), .RN(n1059), .QN(n477)
         );
  DFFR_X1 \registers_reg[15][2]  ( .D(n3031), .CK(CLK), .RN(n1059), .QN(n478)
         );
  DFFR_X1 \registers_reg[15][1]  ( .D(n3030), .CK(CLK), .RN(n1059), .QN(n479)
         );
  DFFR_X1 \registers_reg[15][0]  ( .D(n3029), .CK(CLK), .RN(n1059), .QN(n480)
         );
  DFFR_X1 \registers_reg[16][31]  ( .D(n3028), .CK(CLK), .RN(n1059), .QN(n481)
         );
  DFFR_X1 \registers_reg[16][30]  ( .D(n3027), .CK(CLK), .RN(n1059), .QN(n482)
         );
  DFFR_X1 \registers_reg[16][29]  ( .D(n3026), .CK(CLK), .RN(n1059), .QN(n483)
         );
  DFFR_X1 \registers_reg[16][28]  ( .D(n3025), .CK(CLK), .RN(n1059), .QN(n484)
         );
  DFFR_X1 \registers_reg[16][27]  ( .D(n3024), .CK(CLK), .RN(n1059), .QN(n485)
         );
  DFFR_X1 \registers_reg[16][26]  ( .D(n3023), .CK(CLK), .RN(n1059), .QN(n486)
         );
  DFFR_X1 \registers_reg[16][25]  ( .D(n3022), .CK(CLK), .RN(n1058), .QN(n487)
         );
  DFFR_X1 \registers_reg[16][24]  ( .D(n3021), .CK(CLK), .RN(n1058), .QN(n488)
         );
  DFFR_X1 \registers_reg[16][23]  ( .D(n3020), .CK(CLK), .RN(n1058), .QN(n489)
         );
  DFFR_X1 \registers_reg[16][22]  ( .D(n3019), .CK(CLK), .RN(n1058), .QN(n490)
         );
  DFFR_X1 \registers_reg[16][21]  ( .D(n3018), .CK(CLK), .RN(n1058), .QN(n491)
         );
  DFFR_X1 \registers_reg[16][20]  ( .D(n3017), .CK(CLK), .RN(n1058), .QN(n492)
         );
  DFFR_X1 \registers_reg[16][19]  ( .D(n3016), .CK(CLK), .RN(n1058), .QN(n493)
         );
  DFFR_X1 \registers_reg[16][18]  ( .D(n3015), .CK(CLK), .RN(n1058), .QN(n494)
         );
  DFFR_X1 \registers_reg[16][17]  ( .D(n3014), .CK(CLK), .RN(n1058), .QN(n495)
         );
  DFFR_X1 \registers_reg[16][16]  ( .D(n3013), .CK(CLK), .RN(n1058), .QN(n496)
         );
  DFFR_X1 \registers_reg[16][15]  ( .D(n3012), .CK(CLK), .RN(n1058), .QN(n497)
         );
  DFFR_X1 \registers_reg[16][14]  ( .D(n3011), .CK(CLK), .RN(n1057), .QN(n498)
         );
  DFFR_X1 \registers_reg[16][13]  ( .D(n3010), .CK(CLK), .RN(n1057), .QN(n499)
         );
  DFFR_X1 \registers_reg[16][12]  ( .D(n3009), .CK(CLK), .RN(n1057), .QN(n500)
         );
  DFFR_X1 \registers_reg[16][11]  ( .D(n3008), .CK(CLK), .RN(n1057), .QN(n501)
         );
  DFFR_X1 \registers_reg[16][10]  ( .D(n3007), .CK(CLK), .RN(n1057), .QN(n502)
         );
  DFFR_X1 \registers_reg[16][9]  ( .D(n3006), .CK(CLK), .RN(n1057), .QN(n503)
         );
  DFFR_X1 \registers_reg[16][8]  ( .D(n3005), .CK(CLK), .RN(n1057), .QN(n504)
         );
  DFFR_X1 \registers_reg[16][7]  ( .D(n3004), .CK(CLK), .RN(n1057), .QN(n505)
         );
  DFFR_X1 \registers_reg[16][6]  ( .D(n3003), .CK(CLK), .RN(n1057), .QN(n506)
         );
  DFFR_X1 \registers_reg[16][5]  ( .D(n3002), .CK(CLK), .RN(n1057), .QN(n507)
         );
  DFFR_X1 \registers_reg[16][4]  ( .D(n3001), .CK(CLK), .RN(n1057), .QN(n508)
         );
  DFFR_X1 \registers_reg[16][3]  ( .D(n3000), .CK(CLK), .RN(n1056), .QN(n509)
         );
  DFFR_X1 \registers_reg[16][2]  ( .D(n2999), .CK(CLK), .RN(n1056), .QN(n510)
         );
  DFFR_X1 \registers_reg[16][1]  ( .D(n2998), .CK(CLK), .RN(n1056), .QN(n511)
         );
  DFFR_X1 \registers_reg[16][0]  ( .D(n2997), .CK(CLK), .RN(n1056), .QN(n512)
         );
  DFFR_X1 \registers_reg[17][31]  ( .D(n2996), .CK(CLK), .RN(n1056), .QN(n513)
         );
  DFFR_X1 \registers_reg[17][30]  ( .D(n2995), .CK(CLK), .RN(n1056), .QN(n514)
         );
  DFFR_X1 \registers_reg[17][29]  ( .D(n2994), .CK(CLK), .RN(n1056), .QN(n515)
         );
  DFFR_X1 \registers_reg[17][28]  ( .D(n2993), .CK(CLK), .RN(n1056), .QN(n516)
         );
  DFFR_X1 \registers_reg[17][27]  ( .D(n2992), .CK(CLK), .RN(n1056), .QN(n517)
         );
  DFFR_X1 \registers_reg[17][26]  ( .D(n2991), .CK(CLK), .RN(n1056), .QN(n518)
         );
  DFFR_X1 \registers_reg[17][25]  ( .D(n2990), .CK(CLK), .RN(n1056), .QN(n519)
         );
  DFFR_X1 \registers_reg[17][24]  ( .D(n2989), .CK(CLK), .RN(n1055), .QN(n520)
         );
  DFFR_X1 \registers_reg[17][23]  ( .D(n2988), .CK(CLK), .RN(n1055), .QN(n521)
         );
  DFFR_X1 \registers_reg[17][22]  ( .D(n2987), .CK(CLK), .RN(n1055), .QN(n522)
         );
  DFFR_X1 \registers_reg[17][21]  ( .D(n2986), .CK(CLK), .RN(n1055), .QN(n523)
         );
  DFFR_X1 \registers_reg[17][20]  ( .D(n2985), .CK(CLK), .RN(n1055), .QN(n524)
         );
  DFFR_X1 \registers_reg[17][19]  ( .D(n2984), .CK(CLK), .RN(n1055), .QN(n525)
         );
  DFFR_X1 \registers_reg[17][18]  ( .D(n2983), .CK(CLK), .RN(n1055), .QN(n526)
         );
  DFFR_X1 \registers_reg[17][17]  ( .D(n2982), .CK(CLK), .RN(n1055), .QN(n527)
         );
  DFFR_X1 \registers_reg[17][16]  ( .D(n2981), .CK(CLK), .RN(n1055), .QN(n528)
         );
  DFFR_X1 \registers_reg[17][15]  ( .D(n2980), .CK(CLK), .RN(n1055), .QN(n529)
         );
  DFFR_X1 \registers_reg[17][14]  ( .D(n2979), .CK(CLK), .RN(n1055), .QN(n530)
         );
  DFFR_X1 \registers_reg[17][13]  ( .D(n2978), .CK(CLK), .RN(n1054), .QN(n531)
         );
  DFFR_X1 \registers_reg[17][12]  ( .D(n2977), .CK(CLK), .RN(n1054), .QN(n532)
         );
  DFFR_X1 \registers_reg[17][11]  ( .D(n2976), .CK(CLK), .RN(n1054), .QN(n533)
         );
  DFFR_X1 \registers_reg[17][10]  ( .D(n2975), .CK(CLK), .RN(n1054), .QN(n534)
         );
  DFFR_X1 \registers_reg[17][9]  ( .D(n2974), .CK(CLK), .RN(n1054), .QN(n535)
         );
  DFFR_X1 \registers_reg[17][8]  ( .D(n2973), .CK(CLK), .RN(n1054), .QN(n536)
         );
  DFFR_X1 \registers_reg[17][7]  ( .D(n2972), .CK(CLK), .RN(n1054), .QN(n537)
         );
  DFFR_X1 \registers_reg[17][6]  ( .D(n2971), .CK(CLK), .RN(n1054), .QN(n538)
         );
  DFFR_X1 \registers_reg[17][5]  ( .D(n2970), .CK(CLK), .RN(n1054), .QN(n539)
         );
  DFFR_X1 \registers_reg[17][4]  ( .D(n2969), .CK(CLK), .RN(n1054), .QN(n540)
         );
  DFFR_X1 \registers_reg[17][3]  ( .D(n2968), .CK(CLK), .RN(n1054), .QN(n541)
         );
  DFFR_X1 \registers_reg[17][2]  ( .D(n2967), .CK(CLK), .RN(n1053), .QN(n542)
         );
  DFFR_X1 \registers_reg[17][1]  ( .D(n2966), .CK(CLK), .RN(n1053), .QN(n543)
         );
  DFFR_X1 \registers_reg[17][0]  ( .D(n2965), .CK(CLK), .RN(n1053), .QN(n544)
         );
  DFFR_X1 \registers_reg[18][31]  ( .D(n3578), .CK(CLK), .RN(n1053), .Q(
        \registers[18][31] ) );
  DFFR_X1 \registers_reg[18][30]  ( .D(n3577), .CK(CLK), .RN(n1053), .Q(
        \registers[18][30] ) );
  DFFR_X1 \registers_reg[18][29]  ( .D(n3576), .CK(CLK), .RN(n1053), .Q(
        \registers[18][29] ) );
  DFFR_X1 \registers_reg[18][28]  ( .D(n3575), .CK(CLK), .RN(n1053), .Q(
        \registers[18][28] ) );
  DFFR_X1 \registers_reg[18][27]  ( .D(n3574), .CK(CLK), .RN(n1053), .Q(
        \registers[18][27] ) );
  DFFR_X1 \registers_reg[18][26]  ( .D(n3573), .CK(CLK), .RN(n1053), .Q(
        \registers[18][26] ) );
  DFFR_X1 \registers_reg[18][25]  ( .D(n3572), .CK(CLK), .RN(n1053), .Q(
        \registers[18][25] ) );
  DFFR_X1 \registers_reg[18][24]  ( .D(n3571), .CK(CLK), .RN(n1053), .Q(
        \registers[18][24] ) );
  DFFR_X1 \registers_reg[18][23]  ( .D(n3570), .CK(CLK), .RN(n1052), .Q(
        \registers[18][23] ) );
  DFFR_X1 \registers_reg[18][22]  ( .D(n3569), .CK(CLK), .RN(n1052), .Q(
        \registers[18][22] ) );
  DFFR_X1 \registers_reg[18][21]  ( .D(n3568), .CK(CLK), .RN(n1052), .Q(
        \registers[18][21] ) );
  DFFR_X1 \registers_reg[18][20]  ( .D(n3567), .CK(CLK), .RN(n1052), .Q(
        \registers[18][20] ) );
  DFFR_X1 \registers_reg[18][19]  ( .D(n3566), .CK(CLK), .RN(n1052), .Q(
        \registers[18][19] ) );
  DFFR_X1 \registers_reg[18][18]  ( .D(n3565), .CK(CLK), .RN(n1052), .Q(
        \registers[18][18] ) );
  DFFR_X1 \registers_reg[18][17]  ( .D(n3564), .CK(CLK), .RN(n1052), .Q(
        \registers[18][17] ) );
  DFFR_X1 \registers_reg[18][16]  ( .D(n3563), .CK(CLK), .RN(n1052), .Q(
        \registers[18][16] ) );
  DFFR_X1 \registers_reg[18][15]  ( .D(n3562), .CK(CLK), .RN(n1052), .Q(
        \registers[18][15] ) );
  DFFR_X1 \registers_reg[18][14]  ( .D(n3561), .CK(CLK), .RN(n1052), .Q(
        \registers[18][14] ) );
  DFFR_X1 \registers_reg[18][13]  ( .D(n3560), .CK(CLK), .RN(n1052), .Q(
        \registers[18][13] ) );
  DFFR_X1 \registers_reg[18][12]  ( .D(n3559), .CK(CLK), .RN(n1051), .Q(
        \registers[18][12] ) );
  DFFR_X1 \registers_reg[18][11]  ( .D(n3558), .CK(CLK), .RN(n1051), .Q(
        \registers[18][11] ) );
  DFFR_X1 \registers_reg[18][10]  ( .D(n3557), .CK(CLK), .RN(n1051), .Q(
        \registers[18][10] ) );
  DFFR_X1 \registers_reg[18][9]  ( .D(n3556), .CK(CLK), .RN(n1051), .Q(
        \registers[18][9] ) );
  DFFR_X1 \registers_reg[18][8]  ( .D(n3555), .CK(CLK), .RN(n1051), .Q(
        \registers[18][8] ) );
  DFFR_X1 \registers_reg[18][7]  ( .D(n3554), .CK(CLK), .RN(n1051), .Q(
        \registers[18][7] ) );
  DFFR_X1 \registers_reg[18][6]  ( .D(n3553), .CK(CLK), .RN(n1051), .Q(
        \registers[18][6] ) );
  DFFR_X1 \registers_reg[18][5]  ( .D(n3552), .CK(CLK), .RN(n1051), .Q(
        \registers[18][5] ) );
  DFFR_X1 \registers_reg[18][4]  ( .D(n3551), .CK(CLK), .RN(n1051), .Q(
        \registers[18][4] ) );
  DFFR_X1 \registers_reg[18][3]  ( .D(n3550), .CK(CLK), .RN(n1051), .Q(
        \registers[18][3] ) );
  DFFR_X1 \registers_reg[18][2]  ( .D(n3549), .CK(CLK), .RN(n1051), .Q(
        \registers[18][2] ) );
  DFFR_X1 \registers_reg[18][1]  ( .D(n3548), .CK(CLK), .RN(n1050), .Q(
        \registers[18][1] ) );
  DFFR_X1 \registers_reg[18][0]  ( .D(n3547), .CK(CLK), .RN(n1050), .Q(
        \registers[18][0] ) );
  DFFR_X1 \registers_reg[19][31]  ( .D(n3610), .CK(CLK), .RN(n1050), .Q(
        \registers[19][31] ) );
  DFFR_X1 \registers_reg[19][30]  ( .D(n3609), .CK(CLK), .RN(n1050), .Q(
        \registers[19][30] ) );
  DFFR_X1 \registers_reg[19][29]  ( .D(n3608), .CK(CLK), .RN(n1050), .Q(
        \registers[19][29] ) );
  DFFR_X1 \registers_reg[19][28]  ( .D(n3607), .CK(CLK), .RN(n1050), .Q(
        \registers[19][28] ) );
  DFFR_X1 \registers_reg[19][27]  ( .D(n3606), .CK(CLK), .RN(n1050), .Q(
        \registers[19][27] ) );
  DFFR_X1 \registers_reg[19][26]  ( .D(n3605), .CK(CLK), .RN(n1050), .Q(
        \registers[19][26] ) );
  DFFR_X1 \registers_reg[19][25]  ( .D(n3604), .CK(CLK), .RN(n1050), .Q(
        \registers[19][25] ) );
  DFFR_X1 \registers_reg[19][24]  ( .D(n3603), .CK(CLK), .RN(n1050), .Q(
        \registers[19][24] ) );
  DFFR_X1 \registers_reg[19][23]  ( .D(n3602), .CK(CLK), .RN(n1050), .Q(
        \registers[19][23] ) );
  DFFR_X1 \registers_reg[19][22]  ( .D(n3601), .CK(CLK), .RN(n1049), .Q(
        \registers[19][22] ) );
  DFFR_X1 \registers_reg[19][21]  ( .D(n3600), .CK(CLK), .RN(n1049), .Q(
        \registers[19][21] ) );
  DFFR_X1 \registers_reg[19][20]  ( .D(n3599), .CK(CLK), .RN(n1049), .Q(
        \registers[19][20] ) );
  DFFR_X1 \registers_reg[19][19]  ( .D(n3598), .CK(CLK), .RN(n1049), .Q(
        \registers[19][19] ) );
  DFFR_X1 \registers_reg[19][18]  ( .D(n3597), .CK(CLK), .RN(n1049), .Q(
        \registers[19][18] ) );
  DFFR_X1 \registers_reg[19][17]  ( .D(n3596), .CK(CLK), .RN(n1049), .Q(
        \registers[19][17] ) );
  DFFR_X1 \registers_reg[19][16]  ( .D(n3595), .CK(CLK), .RN(n1049), .Q(
        \registers[19][16] ) );
  DFFR_X1 \registers_reg[19][15]  ( .D(n3594), .CK(CLK), .RN(n1049), .Q(
        \registers[19][15] ) );
  DFFR_X1 \registers_reg[19][14]  ( .D(n3593), .CK(CLK), .RN(n1049), .Q(
        \registers[19][14] ) );
  DFFR_X1 \registers_reg[19][13]  ( .D(n3592), .CK(CLK), .RN(n1049), .Q(
        \registers[19][13] ) );
  DFFR_X1 \registers_reg[19][12]  ( .D(n3591), .CK(CLK), .RN(n1049), .Q(
        \registers[19][12] ) );
  DFFR_X1 \registers_reg[19][11]  ( .D(n3590), .CK(CLK), .RN(n1048), .Q(
        \registers[19][11] ) );
  DFFR_X1 \registers_reg[19][10]  ( .D(n3589), .CK(CLK), .RN(n1048), .Q(
        \registers[19][10] ) );
  DFFR_X1 \registers_reg[19][9]  ( .D(n3588), .CK(CLK), .RN(n1048), .Q(
        \registers[19][9] ) );
  DFFR_X1 \registers_reg[19][8]  ( .D(n3587), .CK(CLK), .RN(n1048), .Q(
        \registers[19][8] ) );
  DFFR_X1 \registers_reg[19][7]  ( .D(n3586), .CK(CLK), .RN(n1048), .Q(
        \registers[19][7] ) );
  DFFR_X1 \registers_reg[19][6]  ( .D(n3585), .CK(CLK), .RN(n1048), .Q(
        \registers[19][6] ) );
  DFFR_X1 \registers_reg[19][5]  ( .D(n3584), .CK(CLK), .RN(n1048), .Q(
        \registers[19][5] ) );
  DFFR_X1 \registers_reg[19][4]  ( .D(n3583), .CK(CLK), .RN(n1048), .Q(
        \registers[19][4] ) );
  DFFR_X1 \registers_reg[19][3]  ( .D(n3582), .CK(CLK), .RN(n1048), .Q(
        \registers[19][3] ) );
  DFFR_X1 \registers_reg[19][2]  ( .D(n3581), .CK(CLK), .RN(n1048), .Q(
        \registers[19][2] ) );
  DFFR_X1 \registers_reg[19][1]  ( .D(n3580), .CK(CLK), .RN(n1048), .Q(
        \registers[19][1] ) );
  DFFR_X1 \registers_reg[19][0]  ( .D(n3579), .CK(CLK), .RN(n1047), .Q(
        \registers[19][0] ) );
  DFFR_X1 \registers_reg[20][31]  ( .D(n2964), .CK(CLK), .RN(n1047), .QN(n609)
         );
  DFFR_X1 \registers_reg[20][30]  ( .D(n2963), .CK(CLK), .RN(n1047), .QN(n610)
         );
  DFFR_X1 \registers_reg[20][29]  ( .D(n2962), .CK(CLK), .RN(n1047), .QN(n611)
         );
  DFFR_X1 \registers_reg[20][28]  ( .D(n2961), .CK(CLK), .RN(n1047), .QN(n612)
         );
  DFFR_X1 \registers_reg[20][27]  ( .D(n2960), .CK(CLK), .RN(n1047), .QN(n613)
         );
  DFFR_X1 \registers_reg[20][26]  ( .D(n2959), .CK(CLK), .RN(n1047), .QN(n614)
         );
  DFFR_X1 \registers_reg[20][25]  ( .D(n2958), .CK(CLK), .RN(n1047), .QN(n615)
         );
  DFFR_X1 \registers_reg[20][24]  ( .D(n2957), .CK(CLK), .RN(n1047), .QN(n616)
         );
  DFFR_X1 \registers_reg[20][23]  ( .D(n2956), .CK(CLK), .RN(n1047), .QN(n617)
         );
  DFFR_X1 \registers_reg[20][22]  ( .D(n2955), .CK(CLK), .RN(n1047), .QN(n618)
         );
  DFFR_X1 \registers_reg[20][21]  ( .D(n2954), .CK(CLK), .RN(n1046), .QN(n619)
         );
  DFFR_X1 \registers_reg[20][20]  ( .D(n2953), .CK(CLK), .RN(n1046), .QN(n620)
         );
  DFFR_X1 \registers_reg[20][19]  ( .D(n2952), .CK(CLK), .RN(n1046), .QN(n621)
         );
  DFFR_X1 \registers_reg[20][18]  ( .D(n2951), .CK(CLK), .RN(n1046), .QN(n622)
         );
  DFFR_X1 \registers_reg[20][17]  ( .D(n2950), .CK(CLK), .RN(n1046), .QN(n623)
         );
  DFFR_X1 \registers_reg[20][16]  ( .D(n2949), .CK(CLK), .RN(n1046), .QN(n624)
         );
  DFFR_X1 \registers_reg[20][15]  ( .D(n2948), .CK(CLK), .RN(n1046), .QN(n625)
         );
  DFFR_X1 \registers_reg[20][14]  ( .D(n2947), .CK(CLK), .RN(n1046), .QN(n626)
         );
  DFFR_X1 \registers_reg[20][13]  ( .D(n2946), .CK(CLK), .RN(n1046), .QN(n627)
         );
  DFFR_X1 \registers_reg[20][12]  ( .D(n2945), .CK(CLK), .RN(n1046), .QN(n628)
         );
  DFFR_X1 \registers_reg[20][11]  ( .D(n2944), .CK(CLK), .RN(n1046), .QN(n629)
         );
  DFFR_X1 \registers_reg[20][10]  ( .D(n2943), .CK(CLK), .RN(n1045), .QN(n630)
         );
  DFFR_X1 \registers_reg[20][9]  ( .D(n2942), .CK(CLK), .RN(n1045), .QN(n631)
         );
  DFFR_X1 \registers_reg[20][8]  ( .D(n2941), .CK(CLK), .RN(n1045), .QN(n632)
         );
  DFFR_X1 \registers_reg[20][7]  ( .D(n2940), .CK(CLK), .RN(n1045), .QN(n633)
         );
  DFFR_X1 \registers_reg[20][6]  ( .D(n2939), .CK(CLK), .RN(n1045), .QN(n634)
         );
  DFFR_X1 \registers_reg[20][5]  ( .D(n2938), .CK(CLK), .RN(n1045), .QN(n635)
         );
  DFFR_X1 \registers_reg[20][4]  ( .D(n2937), .CK(CLK), .RN(n1045), .QN(n636)
         );
  DFFR_X1 \registers_reg[20][3]  ( .D(n2936), .CK(CLK), .RN(n1045), .QN(n637)
         );
  DFFR_X1 \registers_reg[20][2]  ( .D(n2935), .CK(CLK), .RN(n1045), .QN(n638)
         );
  DFFR_X1 \registers_reg[20][1]  ( .D(n2934), .CK(CLK), .RN(n1045), .QN(n639)
         );
  DFFR_X1 \registers_reg[20][0]  ( .D(n2933), .CK(CLK), .RN(n1045), .QN(n640)
         );
  DFFR_X1 \registers_reg[21][31]  ( .D(n2932), .CK(CLK), .RN(n1044), .QN(n641)
         );
  DFFR_X1 \registers_reg[21][30]  ( .D(n2931), .CK(CLK), .RN(n1044), .QN(n642)
         );
  DFFR_X1 \registers_reg[21][29]  ( .D(n2930), .CK(CLK), .RN(n1044), .QN(n643)
         );
  DFFR_X1 \registers_reg[21][28]  ( .D(n2929), .CK(CLK), .RN(n1044), .QN(n644)
         );
  DFFR_X1 \registers_reg[21][27]  ( .D(n2928), .CK(CLK), .RN(n1044), .QN(n645)
         );
  DFFR_X1 \registers_reg[21][26]  ( .D(n2927), .CK(CLK), .RN(n1044), .QN(n646)
         );
  DFFR_X1 \registers_reg[21][25]  ( .D(n2926), .CK(CLK), .RN(n1044), .QN(n647)
         );
  DFFR_X1 \registers_reg[21][24]  ( .D(n2925), .CK(CLK), .RN(n1044), .QN(n648)
         );
  DFFR_X1 \registers_reg[21][23]  ( .D(n2924), .CK(CLK), .RN(n1044), .QN(n649)
         );
  DFFR_X1 \registers_reg[21][22]  ( .D(n2923), .CK(CLK), .RN(n1044), .QN(n650)
         );
  DFFR_X1 \registers_reg[21][21]  ( .D(n2922), .CK(CLK), .RN(n1044), .QN(n651)
         );
  DFFR_X1 \registers_reg[21][20]  ( .D(n2921), .CK(CLK), .RN(n1043), .QN(n652)
         );
  DFFR_X1 \registers_reg[21][19]  ( .D(n2920), .CK(CLK), .RN(n1043), .QN(n653)
         );
  DFFR_X1 \registers_reg[21][18]  ( .D(n2919), .CK(CLK), .RN(n1043), .QN(n654)
         );
  DFFR_X1 \registers_reg[21][17]  ( .D(n2918), .CK(CLK), .RN(n1043), .QN(n655)
         );
  DFFR_X1 \registers_reg[21][16]  ( .D(n2917), .CK(CLK), .RN(n1043), .QN(n656)
         );
  DFFR_X1 \registers_reg[21][15]  ( .D(n2916), .CK(CLK), .RN(n1043), .QN(n657)
         );
  DFFR_X1 \registers_reg[21][14]  ( .D(n2915), .CK(CLK), .RN(n1043), .QN(n658)
         );
  DFFR_X1 \registers_reg[21][13]  ( .D(n2914), .CK(CLK), .RN(n1043), .QN(n659)
         );
  DFFR_X1 \registers_reg[21][12]  ( .D(n2913), .CK(CLK), .RN(n1043), .QN(n660)
         );
  DFFR_X1 \registers_reg[21][11]  ( .D(n2912), .CK(CLK), .RN(n1043), .QN(n661)
         );
  DFFR_X1 \registers_reg[21][10]  ( .D(n2911), .CK(CLK), .RN(n1043), .QN(n662)
         );
  DFFR_X1 \registers_reg[21][9]  ( .D(n2910), .CK(CLK), .RN(n1042), .QN(n663)
         );
  DFFR_X1 \registers_reg[21][8]  ( .D(n2909), .CK(CLK), .RN(n1042), .QN(n664)
         );
  DFFR_X1 \registers_reg[21][7]  ( .D(n2908), .CK(CLK), .RN(n1042), .QN(n665)
         );
  DFFR_X1 \registers_reg[21][6]  ( .D(n2907), .CK(CLK), .RN(n1042), .QN(n666)
         );
  DFFR_X1 \registers_reg[21][5]  ( .D(n2906), .CK(CLK), .RN(n1042), .QN(n667)
         );
  DFFR_X1 \registers_reg[21][4]  ( .D(n2905), .CK(CLK), .RN(n1042), .QN(n668)
         );
  DFFR_X1 \registers_reg[21][3]  ( .D(n2904), .CK(CLK), .RN(n1042), .QN(n669)
         );
  DFFR_X1 \registers_reg[21][2]  ( .D(n2903), .CK(CLK), .RN(n1042), .QN(n670)
         );
  DFFR_X1 \registers_reg[21][1]  ( .D(n2902), .CK(CLK), .RN(n1042), .QN(n671)
         );
  DFFR_X1 \registers_reg[21][0]  ( .D(n2901), .CK(CLK), .RN(n1042), .QN(n672)
         );
  DFFR_X1 \registers_reg[22][31]  ( .D(n3642), .CK(CLK), .RN(n1042), .Q(
        \registers[22][31] ) );
  DFFR_X1 \registers_reg[22][30]  ( .D(n3641), .CK(CLK), .RN(n1041), .Q(
        \registers[22][30] ) );
  DFFR_X1 \registers_reg[22][29]  ( .D(n3640), .CK(CLK), .RN(n1041), .Q(
        \registers[22][29] ) );
  DFFR_X1 \registers_reg[22][28]  ( .D(n3639), .CK(CLK), .RN(n1041), .Q(
        \registers[22][28] ) );
  DFFR_X1 \registers_reg[22][27]  ( .D(n3638), .CK(CLK), .RN(n1041), .Q(
        \registers[22][27] ) );
  DFFR_X1 \registers_reg[22][26]  ( .D(n3637), .CK(CLK), .RN(n1041), .Q(
        \registers[22][26] ) );
  DFFR_X1 \registers_reg[22][25]  ( .D(n3636), .CK(CLK), .RN(n1041), .Q(
        \registers[22][25] ) );
  DFFR_X1 \registers_reg[22][24]  ( .D(n3635), .CK(CLK), .RN(n1041), .Q(
        \registers[22][24] ) );
  DFFR_X1 \registers_reg[22][23]  ( .D(n3634), .CK(CLK), .RN(n1041), .Q(
        \registers[22][23] ) );
  DFFR_X1 \registers_reg[22][22]  ( .D(n3633), .CK(CLK), .RN(n1041), .Q(
        \registers[22][22] ) );
  DFFR_X1 \registers_reg[22][21]  ( .D(n3632), .CK(CLK), .RN(n1041), .Q(
        \registers[22][21] ) );
  DFFR_X1 \registers_reg[22][20]  ( .D(n3631), .CK(CLK), .RN(n1041), .Q(
        \registers[22][20] ) );
  DFFR_X1 \registers_reg[22][19]  ( .D(n3630), .CK(CLK), .RN(n1040), .Q(
        \registers[22][19] ) );
  DFFR_X1 \registers_reg[22][18]  ( .D(n3629), .CK(CLK), .RN(n1040), .Q(
        \registers[22][18] ) );
  DFFR_X1 \registers_reg[22][17]  ( .D(n3628), .CK(CLK), .RN(n1040), .Q(
        \registers[22][17] ) );
  DFFR_X1 \registers_reg[22][16]  ( .D(n3627), .CK(CLK), .RN(n1040), .Q(
        \registers[22][16] ) );
  DFFR_X1 \registers_reg[22][15]  ( .D(n3626), .CK(CLK), .RN(n1040), .Q(
        \registers[22][15] ) );
  DFFR_X1 \registers_reg[22][14]  ( .D(n3625), .CK(CLK), .RN(n1040), .Q(
        \registers[22][14] ) );
  DFFR_X1 \registers_reg[22][13]  ( .D(n3624), .CK(CLK), .RN(n1040), .Q(
        \registers[22][13] ) );
  DFFR_X1 \registers_reg[22][12]  ( .D(n3623), .CK(CLK), .RN(n1040), .Q(
        \registers[22][12] ) );
  DFFR_X1 \registers_reg[22][11]  ( .D(n3622), .CK(CLK), .RN(n1040), .Q(
        \registers[22][11] ) );
  DFFR_X1 \registers_reg[22][10]  ( .D(n3621), .CK(CLK), .RN(n1040), .Q(
        \registers[22][10] ) );
  DFFR_X1 \registers_reg[22][9]  ( .D(n3620), .CK(CLK), .RN(n1040), .Q(
        \registers[22][9] ) );
  DFFR_X1 \registers_reg[22][8]  ( .D(n3619), .CK(CLK), .RN(n1039), .Q(
        \registers[22][8] ) );
  DFFR_X1 \registers_reg[22][7]  ( .D(n3618), .CK(CLK), .RN(n1039), .Q(
        \registers[22][7] ) );
  DFFR_X1 \registers_reg[22][6]  ( .D(n3617), .CK(CLK), .RN(n1039), .Q(
        \registers[22][6] ) );
  DFFR_X1 \registers_reg[22][5]  ( .D(n3616), .CK(CLK), .RN(n1039), .Q(
        \registers[22][5] ) );
  DFFR_X1 \registers_reg[22][4]  ( .D(n3615), .CK(CLK), .RN(n1039), .Q(
        \registers[22][4] ) );
  DFFR_X1 \registers_reg[22][3]  ( .D(n3614), .CK(CLK), .RN(n1039), .Q(
        \registers[22][3] ) );
  DFFR_X1 \registers_reg[22][2]  ( .D(n3613), .CK(CLK), .RN(n1039), .Q(
        \registers[22][2] ) );
  DFFR_X1 \registers_reg[22][1]  ( .D(n3612), .CK(CLK), .RN(n1039), .Q(
        \registers[22][1] ) );
  DFFR_X1 \registers_reg[22][0]  ( .D(n3611), .CK(CLK), .RN(n1039), .Q(
        \registers[22][0] ) );
  DFFR_X1 \registers_reg[23][31]  ( .D(n3674), .CK(CLK), .RN(n1039), .Q(
        \registers[23][31] ) );
  DFFR_X1 \registers_reg[23][30]  ( .D(n3673), .CK(CLK), .RN(n1039), .Q(
        \registers[23][30] ) );
  DFFR_X1 \registers_reg[23][29]  ( .D(n3672), .CK(CLK), .RN(n1038), .Q(
        \registers[23][29] ) );
  DFFR_X1 \registers_reg[23][28]  ( .D(n3671), .CK(CLK), .RN(n1038), .Q(
        \registers[23][28] ) );
  DFFR_X1 \registers_reg[23][27]  ( .D(n3670), .CK(CLK), .RN(n1038), .Q(
        \registers[23][27] ) );
  DFFR_X1 \registers_reg[23][26]  ( .D(n3669), .CK(CLK), .RN(n1038), .Q(
        \registers[23][26] ) );
  DFFR_X1 \registers_reg[23][25]  ( .D(n3668), .CK(CLK), .RN(n1038), .Q(
        \registers[23][25] ) );
  DFFR_X1 \registers_reg[23][24]  ( .D(n3667), .CK(CLK), .RN(n1038), .Q(
        \registers[23][24] ) );
  DFFR_X1 \registers_reg[23][23]  ( .D(n3666), .CK(CLK), .RN(n1038), .Q(
        \registers[23][23] ) );
  DFFR_X1 \registers_reg[23][22]  ( .D(n3665), .CK(CLK), .RN(n1038), .Q(
        \registers[23][22] ) );
  DFFR_X1 \registers_reg[23][21]  ( .D(n3664), .CK(CLK), .RN(n1038), .Q(
        \registers[23][21] ) );
  DFFR_X1 \registers_reg[23][20]  ( .D(n3663), .CK(CLK), .RN(n1038), .Q(
        \registers[23][20] ) );
  DFFR_X1 \registers_reg[23][19]  ( .D(n3662), .CK(CLK), .RN(n1038), .Q(
        \registers[23][19] ) );
  DFFR_X1 \registers_reg[23][18]  ( .D(n3661), .CK(CLK), .RN(n1037), .Q(
        \registers[23][18] ) );
  DFFR_X1 \registers_reg[23][17]  ( .D(n3660), .CK(CLK), .RN(n1037), .Q(
        \registers[23][17] ) );
  DFFR_X1 \registers_reg[23][16]  ( .D(n3659), .CK(CLK), .RN(n1037), .Q(
        \registers[23][16] ) );
  DFFR_X1 \registers_reg[23][15]  ( .D(n3658), .CK(CLK), .RN(n1037), .Q(
        \registers[23][15] ) );
  DFFR_X1 \registers_reg[23][14]  ( .D(n3657), .CK(CLK), .RN(n1037), .Q(
        \registers[23][14] ) );
  DFFR_X1 \registers_reg[23][13]  ( .D(n3656), .CK(CLK), .RN(n1037), .Q(
        \registers[23][13] ) );
  DFFR_X1 \registers_reg[23][12]  ( .D(n3655), .CK(CLK), .RN(n1037), .Q(
        \registers[23][12] ) );
  DFFR_X1 \registers_reg[23][11]  ( .D(n3654), .CK(CLK), .RN(n1037), .Q(
        \registers[23][11] ) );
  DFFR_X1 \registers_reg[23][10]  ( .D(n3653), .CK(CLK), .RN(n1037), .Q(
        \registers[23][10] ) );
  DFFR_X1 \registers_reg[23][9]  ( .D(n3652), .CK(CLK), .RN(n1037), .Q(
        \registers[23][9] ) );
  DFFR_X1 \registers_reg[23][8]  ( .D(n3651), .CK(CLK), .RN(n1037), .Q(
        \registers[23][8] ) );
  DFFR_X1 \registers_reg[23][7]  ( .D(n3650), .CK(CLK), .RN(n1036), .Q(
        \registers[23][7] ) );
  DFFR_X1 \registers_reg[23][6]  ( .D(n3649), .CK(CLK), .RN(n1036), .Q(
        \registers[23][6] ) );
  DFFR_X1 \registers_reg[23][5]  ( .D(n3648), .CK(CLK), .RN(n1036), .Q(
        \registers[23][5] ) );
  DFFR_X1 \registers_reg[23][4]  ( .D(n3647), .CK(CLK), .RN(n1036), .Q(
        \registers[23][4] ) );
  DFFR_X1 \registers_reg[23][3]  ( .D(n3646), .CK(CLK), .RN(n1036), .Q(
        \registers[23][3] ) );
  DFFR_X1 \registers_reg[23][2]  ( .D(n3645), .CK(CLK), .RN(n1036), .Q(
        \registers[23][2] ) );
  DFFR_X1 \registers_reg[23][1]  ( .D(n3644), .CK(CLK), .RN(n1036), .Q(
        \registers[23][1] ) );
  DFFR_X1 \registers_reg[23][0]  ( .D(n3643), .CK(CLK), .RN(n1036), .Q(
        \registers[23][0] ) );
  DFFR_X1 \registers_reg[24][31]  ( .D(n3706), .CK(CLK), .RN(n1036), .Q(
        \registers[24][31] ) );
  DFFR_X1 \registers_reg[24][30]  ( .D(n3705), .CK(CLK), .RN(n1036), .Q(
        \registers[24][30] ) );
  DFFR_X1 \registers_reg[24][29]  ( .D(n3704), .CK(CLK), .RN(n1036), .Q(
        \registers[24][29] ) );
  DFFR_X1 \registers_reg[24][28]  ( .D(n3703), .CK(CLK), .RN(n1035), .Q(
        \registers[24][28] ) );
  DFFR_X1 \registers_reg[24][27]  ( .D(n3702), .CK(CLK), .RN(n1035), .Q(
        \registers[24][27] ) );
  DFFR_X1 \registers_reg[24][26]  ( .D(n3701), .CK(CLK), .RN(n1035), .Q(
        \registers[24][26] ) );
  DFFR_X1 \registers_reg[24][25]  ( .D(n3700), .CK(CLK), .RN(n1035), .Q(
        \registers[24][25] ) );
  DFFR_X1 \registers_reg[24][24]  ( .D(n3699), .CK(CLK), .RN(n1035), .Q(
        \registers[24][24] ) );
  DFFR_X1 \registers_reg[24][23]  ( .D(n3698), .CK(CLK), .RN(n1035), .Q(
        \registers[24][23] ) );
  DFFR_X1 \registers_reg[24][22]  ( .D(n3697), .CK(CLK), .RN(n1035), .Q(
        \registers[24][22] ) );
  DFFR_X1 \registers_reg[24][21]  ( .D(n3696), .CK(CLK), .RN(n1035), .Q(
        \registers[24][21] ) );
  DFFR_X1 \registers_reg[24][20]  ( .D(n3695), .CK(CLK), .RN(n1035), .Q(
        \registers[24][20] ) );
  DFFR_X1 \registers_reg[24][19]  ( .D(n3694), .CK(CLK), .RN(n1035), .Q(
        \registers[24][19] ) );
  DFFR_X1 \registers_reg[24][18]  ( .D(n3693), .CK(CLK), .RN(n1035), .Q(
        \registers[24][18] ) );
  DFFR_X1 \registers_reg[24][17]  ( .D(n3692), .CK(CLK), .RN(n1034), .Q(
        \registers[24][17] ) );
  DFFR_X1 \registers_reg[24][16]  ( .D(n3691), .CK(CLK), .RN(n1034), .Q(
        \registers[24][16] ) );
  DFFR_X1 \registers_reg[24][15]  ( .D(n3690), .CK(CLK), .RN(n1034), .Q(
        \registers[24][15] ) );
  DFFR_X1 \registers_reg[24][14]  ( .D(n3689), .CK(CLK), .RN(n1034), .Q(
        \registers[24][14] ) );
  DFFR_X1 \registers_reg[24][13]  ( .D(n3688), .CK(CLK), .RN(n1034), .Q(
        \registers[24][13] ) );
  DFFR_X1 \registers_reg[24][12]  ( .D(n3687), .CK(CLK), .RN(n1034), .Q(
        \registers[24][12] ) );
  DFFR_X1 \registers_reg[24][11]  ( .D(n3686), .CK(CLK), .RN(n1034), .Q(
        \registers[24][11] ) );
  DFFR_X1 \registers_reg[24][10]  ( .D(n3685), .CK(CLK), .RN(n1034), .Q(
        \registers[24][10] ) );
  DFFR_X1 \registers_reg[24][9]  ( .D(n3684), .CK(CLK), .RN(n1034), .Q(
        \registers[24][9] ) );
  DFFR_X1 \registers_reg[24][8]  ( .D(n3683), .CK(CLK), .RN(n1034), .Q(
        \registers[24][8] ) );
  DFFR_X1 \registers_reg[24][7]  ( .D(n3682), .CK(CLK), .RN(n1034), .Q(
        \registers[24][7] ) );
  DFFR_X1 \registers_reg[24][6]  ( .D(n3681), .CK(CLK), .RN(n1033), .Q(
        \registers[24][6] ) );
  DFFR_X1 \registers_reg[24][5]  ( .D(n3680), .CK(CLK), .RN(n1033), .Q(
        \registers[24][5] ) );
  DFFR_X1 \registers_reg[24][4]  ( .D(n3679), .CK(CLK), .RN(n1033), .Q(
        \registers[24][4] ) );
  DFFR_X1 \registers_reg[24][3]  ( .D(n3678), .CK(CLK), .RN(n1033), .Q(
        \registers[24][3] ) );
  DFFR_X1 \registers_reg[24][2]  ( .D(n3677), .CK(CLK), .RN(n1033), .Q(
        \registers[24][2] ) );
  DFFR_X1 \registers_reg[24][1]  ( .D(n3676), .CK(CLK), .RN(n1033), .Q(
        \registers[24][1] ) );
  DFFR_X1 \registers_reg[24][0]  ( .D(n3675), .CK(CLK), .RN(n1033), .Q(
        \registers[24][0] ) );
  DFFR_X1 \registers_reg[25][31]  ( .D(n3738), .CK(CLK), .RN(n1033), .Q(
        \registers[25][31] ) );
  DFFR_X1 \registers_reg[25][30]  ( .D(n3737), .CK(CLK), .RN(n1033), .Q(
        \registers[25][30] ) );
  DFFR_X1 \registers_reg[25][29]  ( .D(n3736), .CK(CLK), .RN(n1033), .Q(
        \registers[25][29] ) );
  DFFR_X1 \registers_reg[25][28]  ( .D(n3735), .CK(CLK), .RN(n1033), .Q(
        \registers[25][28] ) );
  DFFR_X1 \registers_reg[25][27]  ( .D(n3734), .CK(CLK), .RN(n1032), .Q(
        \registers[25][27] ) );
  DFFR_X1 \registers_reg[25][26]  ( .D(n3733), .CK(CLK), .RN(n1032), .Q(
        \registers[25][26] ) );
  DFFR_X1 \registers_reg[25][25]  ( .D(n3732), .CK(CLK), .RN(n1032), .Q(
        \registers[25][25] ) );
  DFFR_X1 \registers_reg[25][24]  ( .D(n3731), .CK(CLK), .RN(n1032), .Q(
        \registers[25][24] ) );
  DFFR_X1 \registers_reg[25][23]  ( .D(n3730), .CK(CLK), .RN(n1032), .Q(
        \registers[25][23] ) );
  DFFR_X1 \registers_reg[25][22]  ( .D(n3729), .CK(CLK), .RN(n1032), .Q(
        \registers[25][22] ) );
  DFFR_X1 \registers_reg[25][21]  ( .D(n3728), .CK(CLK), .RN(n1032), .Q(
        \registers[25][21] ) );
  DFFR_X1 \registers_reg[25][20]  ( .D(n3727), .CK(CLK), .RN(n1032), .Q(
        \registers[25][20] ) );
  DFFR_X1 \registers_reg[25][19]  ( .D(n3726), .CK(CLK), .RN(n1032), .Q(
        \registers[25][19] ) );
  DFFR_X1 \registers_reg[25][18]  ( .D(n3725), .CK(CLK), .RN(n1032), .Q(
        \registers[25][18] ) );
  DFFR_X1 \registers_reg[25][17]  ( .D(n3724), .CK(CLK), .RN(n1032), .Q(
        \registers[25][17] ) );
  DFFR_X1 \registers_reg[25][16]  ( .D(n3723), .CK(CLK), .RN(n1031), .Q(
        \registers[25][16] ) );
  DFFR_X1 \registers_reg[25][15]  ( .D(n3722), .CK(CLK), .RN(n1031), .Q(
        \registers[25][15] ) );
  DFFR_X1 \registers_reg[25][14]  ( .D(n3721), .CK(CLK), .RN(n1031), .Q(
        \registers[25][14] ) );
  DFFR_X1 \registers_reg[25][13]  ( .D(n3720), .CK(CLK), .RN(n1031), .Q(
        \registers[25][13] ) );
  DFFR_X1 \registers_reg[25][12]  ( .D(n3719), .CK(CLK), .RN(n1031), .Q(
        \registers[25][12] ) );
  DFFR_X1 \registers_reg[25][11]  ( .D(n3718), .CK(CLK), .RN(n1031), .Q(
        \registers[25][11] ) );
  DFFR_X1 \registers_reg[25][10]  ( .D(n3717), .CK(CLK), .RN(n1031), .Q(
        \registers[25][10] ) );
  DFFR_X1 \registers_reg[25][9]  ( .D(n3716), .CK(CLK), .RN(n1031), .Q(
        \registers[25][9] ) );
  DFFR_X1 \registers_reg[25][8]  ( .D(n3715), .CK(CLK), .RN(n1031), .Q(
        \registers[25][8] ) );
  DFFR_X1 \registers_reg[25][7]  ( .D(n3714), .CK(CLK), .RN(n1031), .Q(
        \registers[25][7] ) );
  DFFR_X1 \registers_reg[25][6]  ( .D(n3713), .CK(CLK), .RN(n1031), .Q(
        \registers[25][6] ) );
  DFFR_X1 \registers_reg[25][5]  ( .D(n3712), .CK(CLK), .RN(n1030), .Q(
        \registers[25][5] ) );
  DFFR_X1 \registers_reg[25][4]  ( .D(n3711), .CK(CLK), .RN(n1030), .Q(
        \registers[25][4] ) );
  DFFR_X1 \registers_reg[25][3]  ( .D(n3710), .CK(CLK), .RN(n1030), .Q(
        \registers[25][3] ) );
  DFFR_X1 \registers_reg[25][2]  ( .D(n3709), .CK(CLK), .RN(n1030), .Q(
        \registers[25][2] ) );
  DFFR_X1 \registers_reg[25][1]  ( .D(n3708), .CK(CLK), .RN(n1030), .Q(
        \registers[25][1] ) );
  DFFR_X1 \registers_reg[25][0]  ( .D(n3707), .CK(CLK), .RN(n1030), .Q(
        \registers[25][0] ) );
  DFFR_X1 \registers_reg[26][31]  ( .D(n2900), .CK(CLK), .RN(n1030), .QN(n801)
         );
  DFFR_X1 \registers_reg[26][30]  ( .D(n2899), .CK(CLK), .RN(n1030), .QN(n802)
         );
  DFFR_X1 \registers_reg[26][29]  ( .D(n2898), .CK(CLK), .RN(n1030), .QN(n803)
         );
  DFFR_X1 \registers_reg[26][28]  ( .D(n2897), .CK(CLK), .RN(n1030), .QN(n804)
         );
  DFFR_X1 \registers_reg[26][27]  ( .D(n2896), .CK(CLK), .RN(n1030), .QN(n805)
         );
  DFFR_X1 \registers_reg[26][26]  ( .D(n2895), .CK(CLK), .RN(n1029), .QN(n806)
         );
  DFFR_X1 \registers_reg[26][25]  ( .D(n2894), .CK(CLK), .RN(n1029), .QN(n807)
         );
  DFFR_X1 \registers_reg[26][24]  ( .D(n2893), .CK(CLK), .RN(n1029), .QN(n808)
         );
  DFFR_X1 \registers_reg[26][23]  ( .D(n2892), .CK(CLK), .RN(n1029), .QN(n809)
         );
  DFFR_X1 \registers_reg[26][22]  ( .D(n2891), .CK(CLK), .RN(n1029), .QN(n810)
         );
  DFFR_X1 \registers_reg[26][21]  ( .D(n2890), .CK(CLK), .RN(n1029), .QN(n811)
         );
  DFFR_X1 \registers_reg[26][20]  ( .D(n2889), .CK(CLK), .RN(n1029), .QN(n812)
         );
  DFFR_X1 \registers_reg[26][19]  ( .D(n2888), .CK(CLK), .RN(n1029), .QN(n813)
         );
  DFFR_X1 \registers_reg[26][18]  ( .D(n2887), .CK(CLK), .RN(n1029), .QN(n814)
         );
  DFFR_X1 \registers_reg[26][17]  ( .D(n2886), .CK(CLK), .RN(n1029), .QN(n815)
         );
  DFFR_X1 \registers_reg[26][16]  ( .D(n2885), .CK(CLK), .RN(n1029), .QN(n816)
         );
  DFFR_X1 \registers_reg[26][15]  ( .D(n2884), .CK(CLK), .RN(n1028), .QN(n817)
         );
  DFFR_X1 \registers_reg[26][14]  ( .D(n2883), .CK(CLK), .RN(n1028), .QN(n818)
         );
  DFFR_X1 \registers_reg[26][13]  ( .D(n2882), .CK(CLK), .RN(n1028), .QN(n819)
         );
  DFFR_X1 \registers_reg[26][12]  ( .D(n2881), .CK(CLK), .RN(n1028), .QN(n820)
         );
  DFFR_X1 \registers_reg[26][11]  ( .D(n2880), .CK(CLK), .RN(n1028), .QN(n821)
         );
  DFFR_X1 \registers_reg[26][10]  ( .D(n2879), .CK(CLK), .RN(n1028), .QN(n822)
         );
  DFFR_X1 \registers_reg[26][9]  ( .D(n2878), .CK(CLK), .RN(n1028), .QN(n823)
         );
  DFFR_X1 \registers_reg[26][8]  ( .D(n2877), .CK(CLK), .RN(n1028), .QN(n824)
         );
  DFFR_X1 \registers_reg[26][7]  ( .D(n2876), .CK(CLK), .RN(n1028), .QN(n825)
         );
  DFFR_X1 \registers_reg[26][6]  ( .D(n2875), .CK(CLK), .RN(n1028), .QN(n826)
         );
  DFFR_X1 \registers_reg[26][5]  ( .D(n2874), .CK(CLK), .RN(n1028), .QN(n827)
         );
  DFFR_X1 \registers_reg[26][4]  ( .D(n2873), .CK(CLK), .RN(n1027), .QN(n828)
         );
  DFFR_X1 \registers_reg[26][3]  ( .D(n2872), .CK(CLK), .RN(n1027), .QN(n829)
         );
  DFFR_X1 \registers_reg[26][2]  ( .D(n2871), .CK(CLK), .RN(n1027), .QN(n830)
         );
  DFFR_X1 \registers_reg[26][1]  ( .D(n2870), .CK(CLK), .RN(n1027), .QN(n831)
         );
  DFFR_X1 \registers_reg[26][0]  ( .D(n2869), .CK(CLK), .RN(n1027), .QN(n832)
         );
  DFFR_X1 \registers_reg[27][31]  ( .D(n2868), .CK(CLK), .RN(n1027), .QN(n833)
         );
  DFFR_X1 \registers_reg[27][30]  ( .D(n2867), .CK(CLK), .RN(n1027), .QN(n834)
         );
  DFFR_X1 \registers_reg[27][29]  ( .D(n2866), .CK(CLK), .RN(n1027), .QN(n835)
         );
  DFFR_X1 \registers_reg[27][28]  ( .D(n2865), .CK(CLK), .RN(n1027), .QN(n836)
         );
  DFFR_X1 \registers_reg[27][27]  ( .D(n2864), .CK(CLK), .RN(n1027), .QN(n837)
         );
  DFFR_X1 \registers_reg[27][26]  ( .D(n2863), .CK(CLK), .RN(n1027), .QN(n838)
         );
  DFFR_X1 \registers_reg[27][25]  ( .D(n2862), .CK(CLK), .RN(n1026), .QN(n839)
         );
  DFFR_X1 \registers_reg[27][24]  ( .D(n2861), .CK(CLK), .RN(n1026), .QN(n840)
         );
  DFFR_X1 \registers_reg[27][23]  ( .D(n2860), .CK(CLK), .RN(n1026), .QN(n841)
         );
  DFFR_X1 \registers_reg[27][22]  ( .D(n2859), .CK(CLK), .RN(n1026), .QN(n842)
         );
  DFFR_X1 \registers_reg[27][21]  ( .D(n2858), .CK(CLK), .RN(n1026), .QN(n843)
         );
  DFFR_X1 \registers_reg[27][20]  ( .D(n2857), .CK(CLK), .RN(n1026), .QN(n844)
         );
  DFFR_X1 \registers_reg[27][19]  ( .D(n2856), .CK(CLK), .RN(n1026), .QN(n845)
         );
  DFFR_X1 \registers_reg[27][18]  ( .D(n2855), .CK(CLK), .RN(n1026), .QN(n846)
         );
  DFFR_X1 \registers_reg[27][17]  ( .D(n2854), .CK(CLK), .RN(n1026), .QN(n847)
         );
  DFFR_X1 \registers_reg[27][16]  ( .D(n2853), .CK(CLK), .RN(n1026), .QN(n848)
         );
  DFFR_X1 \registers_reg[27][15]  ( .D(n2852), .CK(CLK), .RN(n1026), .QN(n849)
         );
  DFFR_X1 \registers_reg[27][14]  ( .D(n2851), .CK(CLK), .RN(n1025), .QN(n850)
         );
  DFFR_X1 \registers_reg[27][13]  ( .D(n2850), .CK(CLK), .RN(n1025), .QN(n851)
         );
  DFFR_X1 \registers_reg[27][12]  ( .D(n2849), .CK(CLK), .RN(n1025), .QN(n852)
         );
  DFFR_X1 \registers_reg[27][11]  ( .D(n2848), .CK(CLK), .RN(n1025), .QN(n853)
         );
  DFFR_X1 \registers_reg[27][10]  ( .D(n2847), .CK(CLK), .RN(n1025), .QN(n854)
         );
  DFFR_X1 \registers_reg[27][9]  ( .D(n2846), .CK(CLK), .RN(n1025), .QN(n855)
         );
  DFFR_X1 \registers_reg[27][8]  ( .D(n2845), .CK(CLK), .RN(n1025), .QN(n856)
         );
  DFFR_X1 \registers_reg[27][7]  ( .D(n2844), .CK(CLK), .RN(n1025), .QN(n857)
         );
  DFFR_X1 \registers_reg[27][6]  ( .D(n2843), .CK(CLK), .RN(n1025), .QN(n858)
         );
  DFFR_X1 \registers_reg[27][5]  ( .D(n2842), .CK(CLK), .RN(n1025), .QN(n859)
         );
  DFFR_X1 \registers_reg[27][4]  ( .D(n2841), .CK(CLK), .RN(n1025), .QN(n860)
         );
  DFFR_X1 \registers_reg[27][3]  ( .D(n2840), .CK(CLK), .RN(n1024), .QN(n861)
         );
  DFFR_X1 \registers_reg[27][2]  ( .D(n2839), .CK(CLK), .RN(n1024), .QN(n862)
         );
  DFFR_X1 \registers_reg[27][1]  ( .D(n2838), .CK(CLK), .RN(n1024), .QN(n863)
         );
  DFFR_X1 \registers_reg[27][0]  ( .D(n2837), .CK(CLK), .RN(n1024), .QN(n864)
         );
  DFFR_X1 \registers_reg[28][31]  ( .D(n3770), .CK(CLK), .RN(n1024), .Q(
        \registers[28][31] ) );
  DFFR_X1 \registers_reg[28][30]  ( .D(n3769), .CK(CLK), .RN(n1024), .Q(
        \registers[28][30] ) );
  DFFR_X1 \registers_reg[28][29]  ( .D(n3768), .CK(CLK), .RN(n1024), .Q(
        \registers[28][29] ) );
  DFFR_X1 \registers_reg[28][28]  ( .D(n3767), .CK(CLK), .RN(n1024), .Q(
        \registers[28][28] ) );
  DFFR_X1 \registers_reg[28][27]  ( .D(n3766), .CK(CLK), .RN(n1024), .Q(
        \registers[28][27] ) );
  DFFR_X1 \registers_reg[28][26]  ( .D(n3765), .CK(CLK), .RN(n1024), .Q(
        \registers[28][26] ) );
  DFFR_X1 \registers_reg[28][25]  ( .D(n3764), .CK(CLK), .RN(n1024), .Q(
        \registers[28][25] ) );
  DFFR_X1 \registers_reg[28][24]  ( .D(n3763), .CK(CLK), .RN(n1023), .Q(
        \registers[28][24] ) );
  DFFR_X1 \registers_reg[28][23]  ( .D(n3762), .CK(CLK), .RN(n1023), .Q(
        \registers[28][23] ) );
  DFFR_X1 \registers_reg[28][22]  ( .D(n3761), .CK(CLK), .RN(n1023), .Q(
        \registers[28][22] ) );
  DFFR_X1 \registers_reg[28][21]  ( .D(n3760), .CK(CLK), .RN(n1023), .Q(
        \registers[28][21] ) );
  DFFR_X1 \registers_reg[28][20]  ( .D(n3759), .CK(CLK), .RN(n1023), .Q(
        \registers[28][20] ) );
  DFFR_X1 \registers_reg[28][19]  ( .D(n3758), .CK(CLK), .RN(n1023), .Q(
        \registers[28][19] ) );
  DFFR_X1 \registers_reg[28][18]  ( .D(n3757), .CK(CLK), .RN(n1023), .Q(
        \registers[28][18] ) );
  DFFR_X1 \registers_reg[28][17]  ( .D(n3756), .CK(CLK), .RN(n1023), .Q(
        \registers[28][17] ) );
  DFFR_X1 \registers_reg[28][16]  ( .D(n3755), .CK(CLK), .RN(n1023), .Q(
        \registers[28][16] ) );
  DFFR_X1 \registers_reg[28][15]  ( .D(n3754), .CK(CLK), .RN(n1023), .Q(
        \registers[28][15] ) );
  DFFR_X1 \registers_reg[28][14]  ( .D(n3753), .CK(CLK), .RN(n1023), .Q(
        \registers[28][14] ) );
  DFFR_X1 \registers_reg[28][13]  ( .D(n3752), .CK(CLK), .RN(n1022), .Q(
        \registers[28][13] ) );
  DFFR_X1 \registers_reg[28][12]  ( .D(n3751), .CK(CLK), .RN(n1022), .Q(
        \registers[28][12] ) );
  DFFR_X1 \registers_reg[28][11]  ( .D(n3750), .CK(CLK), .RN(n1022), .Q(
        \registers[28][11] ) );
  DFFR_X1 \registers_reg[28][10]  ( .D(n3749), .CK(CLK), .RN(n1022), .Q(
        \registers[28][10] ) );
  DFFR_X1 \registers_reg[28][9]  ( .D(n3748), .CK(CLK), .RN(n1022), .Q(
        \registers[28][9] ) );
  DFFR_X1 \registers_reg[28][8]  ( .D(n3747), .CK(CLK), .RN(n1022), .Q(
        \registers[28][8] ) );
  DFFR_X1 \registers_reg[28][7]  ( .D(n3746), .CK(CLK), .RN(n1022), .Q(
        \registers[28][7] ) );
  DFFR_X1 \registers_reg[28][6]  ( .D(n3745), .CK(CLK), .RN(n1022), .Q(
        \registers[28][6] ) );
  DFFR_X1 \registers_reg[28][5]  ( .D(n3744), .CK(CLK), .RN(n1022), .Q(
        \registers[28][5] ) );
  DFFR_X1 \registers_reg[28][4]  ( .D(n3743), .CK(CLK), .RN(n1022), .Q(
        \registers[28][4] ) );
  DFFR_X1 \registers_reg[28][3]  ( .D(n3742), .CK(CLK), .RN(n1022), .Q(
        \registers[28][3] ) );
  DFFR_X1 \registers_reg[28][2]  ( .D(n3741), .CK(CLK), .RN(n1021), .Q(
        \registers[28][2] ) );
  DFFR_X1 \registers_reg[28][1]  ( .D(n3740), .CK(CLK), .RN(n1021), .Q(
        \registers[28][1] ) );
  DFFR_X1 \registers_reg[28][0]  ( .D(n3739), .CK(CLK), .RN(n1021), .Q(
        \registers[28][0] ) );
  DFFR_X1 \registers_reg[29][31]  ( .D(n3802), .CK(CLK), .RN(n1021), .Q(
        \registers[29][31] ) );
  DFFR_X1 \registers_reg[29][30]  ( .D(n3801), .CK(CLK), .RN(n1021), .Q(
        \registers[29][30] ) );
  DFFR_X1 \registers_reg[29][29]  ( .D(n3800), .CK(CLK), .RN(n1021), .Q(
        \registers[29][29] ) );
  DFFR_X1 \registers_reg[29][28]  ( .D(n3799), .CK(CLK), .RN(n1021), .Q(
        \registers[29][28] ) );
  DFFR_X1 \registers_reg[29][27]  ( .D(n3798), .CK(CLK), .RN(n1021), .Q(
        \registers[29][27] ) );
  DFFR_X1 \registers_reg[29][26]  ( .D(n3797), .CK(CLK), .RN(n1021), .Q(
        \registers[29][26] ) );
  DFFR_X1 \registers_reg[29][25]  ( .D(n3796), .CK(CLK), .RN(n1021), .Q(
        \registers[29][25] ) );
  DFFR_X1 \registers_reg[29][24]  ( .D(n3795), .CK(CLK), .RN(n1021), .Q(
        \registers[29][24] ) );
  DFFR_X1 \registers_reg[29][23]  ( .D(n3794), .CK(CLK), .RN(n1020), .Q(
        \registers[29][23] ) );
  DFFR_X1 \registers_reg[29][22]  ( .D(n3793), .CK(CLK), .RN(n1020), .Q(
        \registers[29][22] ) );
  DFFR_X1 \registers_reg[29][21]  ( .D(n3792), .CK(CLK), .RN(n1020), .Q(
        \registers[29][21] ) );
  DFFR_X1 \registers_reg[29][20]  ( .D(n3791), .CK(CLK), .RN(n1020), .Q(
        \registers[29][20] ) );
  DFFR_X1 \registers_reg[29][19]  ( .D(n3790), .CK(CLK), .RN(n1020), .Q(
        \registers[29][19] ) );
  DFFR_X1 \registers_reg[29][18]  ( .D(n3789), .CK(CLK), .RN(n1020), .Q(
        \registers[29][18] ) );
  DFFR_X1 \registers_reg[29][17]  ( .D(n3788), .CK(CLK), .RN(n1020), .Q(
        \registers[29][17] ) );
  DFFR_X1 \registers_reg[29][16]  ( .D(n3787), .CK(CLK), .RN(n1020), .Q(
        \registers[29][16] ) );
  DFFR_X1 \registers_reg[29][15]  ( .D(n3786), .CK(CLK), .RN(n1020), .Q(
        \registers[29][15] ) );
  DFFR_X1 \registers_reg[29][14]  ( .D(n3785), .CK(CLK), .RN(n1020), .Q(
        \registers[29][14] ) );
  DFFR_X1 \registers_reg[29][13]  ( .D(n3784), .CK(CLK), .RN(n1020), .Q(
        \registers[29][13] ) );
  DFFR_X1 \registers_reg[29][12]  ( .D(n3783), .CK(CLK), .RN(n1019), .Q(
        \registers[29][12] ) );
  DFFR_X1 \registers_reg[29][11]  ( .D(n3782), .CK(CLK), .RN(n1019), .Q(
        \registers[29][11] ) );
  DFFR_X1 \registers_reg[29][10]  ( .D(n3781), .CK(CLK), .RN(n1019), .Q(
        \registers[29][10] ) );
  DFFR_X1 \registers_reg[29][9]  ( .D(n3780), .CK(CLK), .RN(n1019), .Q(
        \registers[29][9] ) );
  DFFR_X1 \registers_reg[29][8]  ( .D(n3779), .CK(CLK), .RN(n1019), .Q(
        \registers[29][8] ) );
  DFFR_X1 \registers_reg[29][7]  ( .D(n3778), .CK(CLK), .RN(n1019), .Q(
        \registers[29][7] ) );
  DFFR_X1 \registers_reg[29][6]  ( .D(n3777), .CK(CLK), .RN(n1019), .Q(
        \registers[29][6] ) );
  DFFR_X1 \registers_reg[29][5]  ( .D(n3776), .CK(CLK), .RN(n1019), .Q(
        \registers[29][5] ) );
  DFFR_X1 \registers_reg[29][4]  ( .D(n3775), .CK(CLK), .RN(n1019), .Q(
        \registers[29][4] ) );
  DFFR_X1 \registers_reg[29][3]  ( .D(n3774), .CK(CLK), .RN(n1019), .Q(
        \registers[29][3] ) );
  DFFR_X1 \registers_reg[29][2]  ( .D(n3773), .CK(CLK), .RN(n1019), .Q(
        \registers[29][2] ) );
  DFFR_X1 \registers_reg[29][1]  ( .D(n3772), .CK(CLK), .RN(n1018), .Q(
        \registers[29][1] ) );
  DFFR_X1 \registers_reg[29][0]  ( .D(n3771), .CK(CLK), .RN(n1018), .Q(
        \registers[29][0] ) );
  DFFR_X1 \registers_reg[30][31]  ( .D(n2836), .CK(CLK), .RN(n1018), .QN(n929)
         );
  DFFR_X1 \registers_reg[30][30]  ( .D(n2835), .CK(CLK), .RN(n1018), .QN(n930)
         );
  DFFR_X1 \registers_reg[30][29]  ( .D(n2834), .CK(CLK), .RN(n1018), .QN(n931)
         );
  DFFR_X1 \registers_reg[30][28]  ( .D(n2833), .CK(CLK), .RN(n1018), .QN(n932)
         );
  DFFR_X1 \registers_reg[30][27]  ( .D(n2832), .CK(CLK), .RN(n1018), .QN(n933)
         );
  DFFR_X1 \registers_reg[30][26]  ( .D(n2831), .CK(CLK), .RN(n1018), .QN(n934)
         );
  DFFR_X1 \registers_reg[30][25]  ( .D(n2830), .CK(CLK), .RN(n1018), .QN(n935)
         );
  DFFR_X1 \registers_reg[30][24]  ( .D(n2829), .CK(CLK), .RN(n1018), .QN(n936)
         );
  DFFR_X1 \registers_reg[30][23]  ( .D(n2828), .CK(CLK), .RN(n1018), .QN(n937)
         );
  DFFR_X1 \registers_reg[30][22]  ( .D(n2827), .CK(CLK), .RN(n1017), .QN(n938)
         );
  DFFR_X1 \registers_reg[30][21]  ( .D(n2826), .CK(CLK), .RN(n1017), .QN(n939)
         );
  DFFR_X1 \registers_reg[30][20]  ( .D(n2825), .CK(CLK), .RN(n1017), .QN(n940)
         );
  DFFR_X1 \registers_reg[30][19]  ( .D(n2824), .CK(CLK), .RN(n1017), .QN(n941)
         );
  DFFR_X1 \registers_reg[30][18]  ( .D(n2823), .CK(CLK), .RN(n1017), .QN(n942)
         );
  DFFR_X1 \registers_reg[30][17]  ( .D(n2822), .CK(CLK), .RN(n1017), .QN(n943)
         );
  DFFR_X1 \registers_reg[30][16]  ( .D(n2821), .CK(CLK), .RN(n1017), .QN(n944)
         );
  DFFR_X1 \registers_reg[30][15]  ( .D(n2820), .CK(CLK), .RN(n1017), .QN(n945)
         );
  DFFR_X1 \registers_reg[30][14]  ( .D(n2819), .CK(CLK), .RN(n1017), .QN(n946)
         );
  DFFR_X1 \registers_reg[30][13]  ( .D(n2818), .CK(CLK), .RN(n1017), .QN(n947)
         );
  DFFR_X1 \registers_reg[30][12]  ( .D(n2817), .CK(CLK), .RN(n1017), .QN(n948)
         );
  DFFR_X1 \registers_reg[30][11]  ( .D(n2816), .CK(CLK), .RN(n1016), .QN(n949)
         );
  DFFR_X1 \registers_reg[30][10]  ( .D(n2815), .CK(CLK), .RN(n1016), .QN(n950)
         );
  DFFR_X1 \registers_reg[30][9]  ( .D(n2814), .CK(CLK), .RN(n1016), .QN(n951)
         );
  DFFR_X1 \registers_reg[30][8]  ( .D(n2813), .CK(CLK), .RN(n1016), .QN(n952)
         );
  DFFR_X1 \registers_reg[30][7]  ( .D(n2812), .CK(CLK), .RN(n1016), .QN(n953)
         );
  DFFR_X1 \registers_reg[30][6]  ( .D(n2811), .CK(CLK), .RN(n1016), .QN(n954)
         );
  DFFR_X1 \registers_reg[30][5]  ( .D(n2810), .CK(CLK), .RN(n1016), .QN(n955)
         );
  DFFR_X1 \registers_reg[30][4]  ( .D(n2809), .CK(CLK), .RN(n1016), .QN(n956)
         );
  DFFR_X1 \registers_reg[30][3]  ( .D(n2808), .CK(CLK), .RN(n1016), .QN(n957)
         );
  DFFR_X1 \registers_reg[30][2]  ( .D(n2807), .CK(CLK), .RN(n1016), .QN(n958)
         );
  DFFR_X1 \registers_reg[30][1]  ( .D(n2806), .CK(CLK), .RN(n1016), .QN(n959)
         );
  DFFR_X1 \registers_reg[30][0]  ( .D(n2805), .CK(CLK), .RN(n1015), .QN(n960)
         );
  DFFR_X1 \registers_reg[31][31]  ( .D(n2804), .CK(CLK), .RN(n1015), .QN(n961)
         );
  DFFR_X1 \registers_reg[31][30]  ( .D(n2803), .CK(CLK), .RN(n1015), .QN(n962)
         );
  DFFR_X1 \registers_reg[31][29]  ( .D(n2802), .CK(CLK), .RN(n1015), .QN(n963)
         );
  DFFR_X1 \registers_reg[31][28]  ( .D(n2801), .CK(CLK), .RN(n1015), .QN(n964)
         );
  DFFR_X1 \registers_reg[31][27]  ( .D(n2800), .CK(CLK), .RN(n1015), .QN(n965)
         );
  DFFR_X1 \registers_reg[31][26]  ( .D(n2799), .CK(CLK), .RN(n1015), .QN(n966)
         );
  DFFR_X1 \registers_reg[31][25]  ( .D(n2798), .CK(CLK), .RN(n1015), .QN(n967)
         );
  DFFR_X1 \registers_reg[31][24]  ( .D(n2797), .CK(CLK), .RN(n1015), .QN(n968)
         );
  DFFR_X1 \registers_reg[31][23]  ( .D(n2796), .CK(CLK), .RN(n1015), .QN(n969)
         );
  DFFR_X1 \registers_reg[31][22]  ( .D(n2795), .CK(CLK), .RN(n1015), .QN(n970)
         );
  DFFR_X1 \registers_reg[31][21]  ( .D(n2794), .CK(CLK), .RN(n1014), .QN(n971)
         );
  DFFR_X1 \registers_reg[31][20]  ( .D(n2793), .CK(CLK), .RN(n1014), .QN(n972)
         );
  DFFR_X1 \registers_reg[31][19]  ( .D(n2792), .CK(CLK), .RN(n1014), .QN(n973)
         );
  DFFR_X1 \registers_reg[31][18]  ( .D(n2791), .CK(CLK), .RN(n1014), .QN(n974)
         );
  DFFR_X1 \registers_reg[31][17]  ( .D(n2790), .CK(CLK), .RN(n1014), .QN(n975)
         );
  DFFR_X1 \registers_reg[31][16]  ( .D(n2789), .CK(CLK), .RN(n1014), .QN(n976)
         );
  DFFR_X1 \registers_reg[31][15]  ( .D(n2788), .CK(CLK), .RN(n1014), .QN(n977)
         );
  DFFR_X1 \registers_reg[31][14]  ( .D(n2787), .CK(CLK), .RN(n1014), .QN(n978)
         );
  DFFR_X1 \registers_reg[31][13]  ( .D(n2786), .CK(CLK), .RN(n1014), .QN(n979)
         );
  DFFR_X1 \registers_reg[31][12]  ( .D(n2785), .CK(CLK), .RN(n1014), .QN(n980)
         );
  DFFR_X1 \registers_reg[31][11]  ( .D(n2784), .CK(CLK), .RN(n1014), .QN(n981)
         );
  DFFR_X1 \registers_reg[31][10]  ( .D(n2783), .CK(CLK), .RN(n1013), .QN(n982)
         );
  DFFR_X1 \registers_reg[31][9]  ( .D(n2782), .CK(CLK), .RN(n1013), .QN(n983)
         );
  DFFR_X1 \registers_reg[31][8]  ( .D(n2781), .CK(CLK), .RN(n1013), .QN(n984)
         );
  DFFR_X1 \registers_reg[31][7]  ( .D(n2780), .CK(CLK), .RN(n1013), .QN(n985)
         );
  DFFR_X1 \registers_reg[31][6]  ( .D(n2779), .CK(CLK), .RN(n1013), .QN(n986)
         );
  DFFR_X1 \registers_reg[31][5]  ( .D(n2778), .CK(CLK), .RN(n1013), .QN(n987)
         );
  DFFR_X1 \registers_reg[31][4]  ( .D(n2777), .CK(CLK), .RN(n1013), .QN(n988)
         );
  DFFR_X1 \registers_reg[31][3]  ( .D(n2776), .CK(CLK), .RN(n1013), .QN(n989)
         );
  DFFR_X1 \registers_reg[31][2]  ( .D(n2775), .CK(CLK), .RN(n1013), .QN(n990)
         );
  DFFR_X1 \registers_reg[31][1]  ( .D(n2774), .CK(CLK), .RN(n1013), .QN(n991)
         );
  DFFR_X1 \registers_reg[31][0]  ( .D(n2773), .CK(CLK), .RN(n1013), .QN(n992)
         );
  DLH_X1 \OUT1_reg[31]  ( .G(n998), .D(N216), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n998), .D(N215), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n998), .D(N214), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n998), .D(N213), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n998), .D(N212), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n998), .D(N211), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n998), .D(N210), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n998), .D(N209), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n998), .D(N208), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n998), .D(N207), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n999), .D(N206), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n999), .D(N205), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n999), .D(N204), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n999), .D(N203), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n999), .D(N202), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n999), .D(N201), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n999), .D(N200), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n999), .D(N199), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n999), .D(N198), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n999), .D(N197), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n1000), .D(N196), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n1000), .D(N195), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n1000), .D(N194), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n1000), .D(N193), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n1000), .D(N192), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n1000), .D(N191), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n1000), .D(N190), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n1000), .D(N189), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n1000), .D(N188), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n1000), .D(N187), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n1001), .D(N186), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n1001), .D(N185), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(n994), .D(N351), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n994), .D(N350), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n994), .D(N349), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n994), .D(N348), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n994), .D(N347), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n994), .D(N346), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n994), .D(N345), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n994), .D(N344), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n994), .D(N343), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n994), .D(N342), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n995), .D(N341), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n995), .D(N340), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n995), .D(N339), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n995), .D(N338), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n995), .D(N337), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n995), .D(N336), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n995), .D(N335), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n995), .D(N334), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n995), .D(N333), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n995), .D(N332), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n996), .D(N331), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n996), .D(N330), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n996), .D(N329), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n996), .D(N328), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n996), .D(N327), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n996), .D(N326), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n996), .D(N325), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n996), .D(N324), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n996), .D(N323), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n996), .D(N322), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n997), .D(N321), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n997), .D(N320), .Q(OUT2[0]) );
  NOR2_X1 U2 ( .A1(n3811), .A2(ADD_RD2[2]), .ZN(n2159) );
  NOR2_X1 U3 ( .A1(n3808), .A2(ADD_RD1[2]), .ZN(n2750) );
  INV_X1 U4 ( .A(n784), .ZN(n777) );
  INV_X1 U5 ( .A(n784), .ZN(n776) );
  INV_X1 U6 ( .A(n775), .ZN(n768) );
  INV_X1 U7 ( .A(n775), .ZN(n767) );
  INV_X1 U8 ( .A(n748), .ZN(n741) );
  INV_X1 U9 ( .A(n748), .ZN(n740) );
  INV_X1 U10 ( .A(n739), .ZN(n732) );
  INV_X1 U11 ( .A(n739), .ZN(n731) );
  INV_X1 U12 ( .A(n730), .ZN(n723) );
  INV_X1 U13 ( .A(n730), .ZN(n722) );
  INV_X1 U14 ( .A(n721), .ZN(n714) );
  INV_X1 U15 ( .A(n721), .ZN(n713) );
  INV_X1 U16 ( .A(n694), .ZN(n687) );
  INV_X1 U17 ( .A(n694), .ZN(n686) );
  INV_X1 U18 ( .A(n685), .ZN(n678) );
  INV_X1 U19 ( .A(n685), .ZN(n677) );
  INV_X1 U20 ( .A(n576), .ZN(n569) );
  INV_X1 U21 ( .A(n576), .ZN(n568) );
  INV_X1 U22 ( .A(n567), .ZN(n560) );
  INV_X1 U23 ( .A(n567), .ZN(n559) );
  INV_X1 U24 ( .A(n412), .ZN(n405) );
  INV_X1 U25 ( .A(n412), .ZN(n404) );
  INV_X1 U26 ( .A(n403), .ZN(n396) );
  INV_X1 U27 ( .A(n403), .ZN(n395) );
  INV_X1 U28 ( .A(n875), .ZN(n868) );
  INV_X1 U29 ( .A(n875), .ZN(n867) );
  INV_X1 U30 ( .A(n866), .ZN(n795) );
  INV_X1 U31 ( .A(n866), .ZN(n794) );
  INV_X1 U32 ( .A(n793), .ZN(n786) );
  INV_X1 U33 ( .A(n793), .ZN(n785) );
  INV_X1 U34 ( .A(n766), .ZN(n759) );
  INV_X1 U35 ( .A(n766), .ZN(n758) );
  INV_X1 U36 ( .A(n757), .ZN(n750) );
  INV_X1 U37 ( .A(n757), .ZN(n749) );
  INV_X1 U38 ( .A(n712), .ZN(n705) );
  INV_X1 U39 ( .A(n712), .ZN(n704) );
  INV_X1 U40 ( .A(n703), .ZN(n696) );
  INV_X1 U41 ( .A(n703), .ZN(n695) );
  INV_X1 U42 ( .A(n676), .ZN(n605) );
  INV_X1 U43 ( .A(n676), .ZN(n604) );
  INV_X1 U44 ( .A(n603), .ZN(n596) );
  INV_X1 U45 ( .A(n603), .ZN(n595) );
  INV_X1 U46 ( .A(n594), .ZN(n587) );
  INV_X1 U47 ( .A(n594), .ZN(n586) );
  INV_X1 U48 ( .A(n585), .ZN(n578) );
  INV_X1 U49 ( .A(n585), .ZN(n577) );
  INV_X1 U50 ( .A(n558), .ZN(n551) );
  INV_X1 U51 ( .A(n558), .ZN(n550) );
  INV_X1 U52 ( .A(n549), .ZN(n414) );
  INV_X1 U53 ( .A(n549), .ZN(n413) );
  INV_X1 U54 ( .A(n911), .ZN(n904) );
  INV_X1 U55 ( .A(n911), .ZN(n903) );
  INV_X1 U56 ( .A(n902), .ZN(n895) );
  INV_X1 U57 ( .A(n902), .ZN(n894) );
  INV_X1 U58 ( .A(n893), .ZN(n886) );
  INV_X1 U59 ( .A(n893), .ZN(n885) );
  INV_X1 U60 ( .A(n884), .ZN(n877) );
  INV_X1 U61 ( .A(n884), .ZN(n876) );
  INV_X1 U62 ( .A(n920), .ZN(n912) );
  INV_X1 U63 ( .A(n920), .ZN(n913) );
  INV_X1 U64 ( .A(n993), .ZN(n922) );
  INV_X1 U65 ( .A(n993), .ZN(n921) );
  BUF_X1 U66 ( .A(n1068), .Z(n993) );
  BUF_X1 U67 ( .A(n1), .Z(n905) );
  BUF_X1 U68 ( .A(n1), .Z(n906) );
  BUF_X1 U69 ( .A(n1), .Z(n907) );
  BUF_X1 U70 ( .A(n1), .Z(n908) );
  BUF_X1 U71 ( .A(n1), .Z(n909) );
  BUF_X1 U72 ( .A(n1), .Z(n910) );
  BUF_X1 U73 ( .A(n2), .Z(n896) );
  BUF_X1 U74 ( .A(n2), .Z(n897) );
  BUF_X1 U75 ( .A(n2), .Z(n898) );
  BUF_X1 U76 ( .A(n2), .Z(n899) );
  BUF_X1 U77 ( .A(n2), .Z(n900) );
  BUF_X1 U78 ( .A(n2), .Z(n901) );
  BUF_X1 U79 ( .A(n3), .Z(n887) );
  BUF_X1 U80 ( .A(n3), .Z(n888) );
  BUF_X1 U81 ( .A(n3), .Z(n889) );
  BUF_X1 U82 ( .A(n3), .Z(n890) );
  BUF_X1 U83 ( .A(n3), .Z(n891) );
  BUF_X1 U84 ( .A(n3), .Z(n892) );
  BUF_X1 U85 ( .A(n4), .Z(n878) );
  BUF_X1 U86 ( .A(n4), .Z(n879) );
  BUF_X1 U87 ( .A(n4), .Z(n880) );
  BUF_X1 U88 ( .A(n4), .Z(n881) );
  BUF_X1 U89 ( .A(n4), .Z(n882) );
  BUF_X1 U90 ( .A(n4), .Z(n883) );
  BUF_X1 U91 ( .A(n5), .Z(n796) );
  BUF_X1 U92 ( .A(n5), .Z(n797) );
  BUF_X1 U93 ( .A(n5), .Z(n798) );
  BUF_X1 U94 ( .A(n5), .Z(n799) );
  BUF_X1 U95 ( .A(n5), .Z(n800) );
  BUF_X1 U96 ( .A(n5), .Z(n865) );
  BUF_X1 U97 ( .A(n6), .Z(n787) );
  BUF_X1 U98 ( .A(n6), .Z(n788) );
  BUF_X1 U99 ( .A(n6), .Z(n789) );
  BUF_X1 U100 ( .A(n6), .Z(n790) );
  BUF_X1 U101 ( .A(n6), .Z(n791) );
  BUF_X1 U102 ( .A(n6), .Z(n792) );
  BUF_X1 U103 ( .A(n7), .Z(n760) );
  BUF_X1 U104 ( .A(n7), .Z(n761) );
  BUF_X1 U105 ( .A(n7), .Z(n762) );
  BUF_X1 U106 ( .A(n7), .Z(n763) );
  BUF_X1 U107 ( .A(n7), .Z(n764) );
  BUF_X1 U108 ( .A(n7), .Z(n765) );
  BUF_X1 U109 ( .A(n8), .Z(n751) );
  BUF_X1 U110 ( .A(n8), .Z(n752) );
  BUF_X1 U111 ( .A(n8), .Z(n753) );
  BUF_X1 U112 ( .A(n8), .Z(n754) );
  BUF_X1 U113 ( .A(n8), .Z(n755) );
  BUF_X1 U114 ( .A(n8), .Z(n756) );
  BUF_X1 U115 ( .A(n9), .Z(n706) );
  BUF_X1 U116 ( .A(n9), .Z(n707) );
  BUF_X1 U117 ( .A(n9), .Z(n708) );
  BUF_X1 U118 ( .A(n9), .Z(n709) );
  BUF_X1 U119 ( .A(n9), .Z(n710) );
  BUF_X1 U120 ( .A(n9), .Z(n711) );
  BUF_X1 U121 ( .A(n10), .Z(n697) );
  BUF_X1 U122 ( .A(n10), .Z(n698) );
  BUF_X1 U123 ( .A(n10), .Z(n699) );
  BUF_X1 U124 ( .A(n10), .Z(n700) );
  BUF_X1 U125 ( .A(n10), .Z(n701) );
  BUF_X1 U126 ( .A(n10), .Z(n702) );
  BUF_X1 U127 ( .A(n11), .Z(n606) );
  BUF_X1 U128 ( .A(n11), .Z(n607) );
  BUF_X1 U129 ( .A(n11), .Z(n608) );
  BUF_X1 U130 ( .A(n11), .Z(n673) );
  BUF_X1 U131 ( .A(n11), .Z(n674) );
  BUF_X1 U132 ( .A(n11), .Z(n675) );
  BUF_X1 U133 ( .A(n12), .Z(n588) );
  BUF_X1 U134 ( .A(n12), .Z(n589) );
  BUF_X1 U135 ( .A(n12), .Z(n590) );
  BUF_X1 U136 ( .A(n12), .Z(n591) );
  BUF_X1 U137 ( .A(n12), .Z(n592) );
  BUF_X1 U138 ( .A(n12), .Z(n593) );
  BUF_X1 U139 ( .A(n13), .Z(n579) );
  BUF_X1 U140 ( .A(n13), .Z(n580) );
  BUF_X1 U141 ( .A(n13), .Z(n581) );
  BUF_X1 U142 ( .A(n13), .Z(n582) );
  BUF_X1 U143 ( .A(n13), .Z(n583) );
  BUF_X1 U144 ( .A(n13), .Z(n584) );
  BUF_X1 U145 ( .A(n14), .Z(n552) );
  BUF_X1 U146 ( .A(n14), .Z(n553) );
  BUF_X1 U147 ( .A(n14), .Z(n554) );
  BUF_X1 U148 ( .A(n14), .Z(n555) );
  BUF_X1 U149 ( .A(n14), .Z(n556) );
  BUF_X1 U150 ( .A(n14), .Z(n557) );
  BUF_X1 U151 ( .A(n15), .Z(n415) );
  BUF_X1 U152 ( .A(n15), .Z(n416) );
  BUF_X1 U153 ( .A(n15), .Z(n545) );
  BUF_X1 U154 ( .A(n15), .Z(n546) );
  BUF_X1 U155 ( .A(n15), .Z(n547) );
  BUF_X1 U156 ( .A(n15), .Z(n548) );
  BUF_X1 U157 ( .A(n16), .Z(n597) );
  BUF_X1 U158 ( .A(n16), .Z(n598) );
  BUF_X1 U159 ( .A(n16), .Z(n599) );
  BUF_X1 U160 ( .A(n16), .Z(n600) );
  BUF_X1 U161 ( .A(n16), .Z(n601) );
  BUF_X1 U162 ( .A(n16), .Z(n602) );
  BUF_X1 U163 ( .A(n1068), .Z(n925) );
  BUF_X1 U164 ( .A(n1068), .Z(n926) );
  BUF_X1 U165 ( .A(n1068), .Z(n927) );
  BUF_X1 U166 ( .A(n1068), .Z(n928) );
  BUF_X1 U167 ( .A(n1068), .Z(n923) );
  BUF_X1 U168 ( .A(n1068), .Z(n924) );
  BUF_X1 U169 ( .A(n1078), .Z(n914) );
  BUF_X1 U170 ( .A(n1078), .Z(n915) );
  BUF_X1 U171 ( .A(n1078), .Z(n916) );
  BUF_X1 U172 ( .A(n1078), .Z(n917) );
  BUF_X1 U173 ( .A(n1078), .Z(n918) );
  BUF_X1 U174 ( .A(n1078), .Z(n919) );
  BUF_X1 U175 ( .A(n1121), .Z(n869) );
  BUF_X1 U176 ( .A(n1121), .Z(n870) );
  BUF_X1 U177 ( .A(n1121), .Z(n871) );
  BUF_X1 U178 ( .A(n1121), .Z(n872) );
  BUF_X1 U179 ( .A(n1121), .Z(n873) );
  BUF_X1 U180 ( .A(n1121), .Z(n874) );
  BUF_X1 U181 ( .A(n1160), .Z(n778) );
  BUF_X1 U182 ( .A(n1160), .Z(n779) );
  BUF_X1 U183 ( .A(n1160), .Z(n780) );
  BUF_X1 U184 ( .A(n1160), .Z(n781) );
  BUF_X1 U185 ( .A(n1160), .Z(n782) );
  BUF_X1 U186 ( .A(n1160), .Z(n783) );
  BUF_X1 U187 ( .A(n1193), .Z(n769) );
  BUF_X1 U188 ( .A(n1193), .Z(n770) );
  BUF_X1 U189 ( .A(n1193), .Z(n771) );
  BUF_X1 U190 ( .A(n1193), .Z(n772) );
  BUF_X1 U191 ( .A(n1193), .Z(n773) );
  BUF_X1 U192 ( .A(n1193), .Z(n774) );
  BUF_X1 U193 ( .A(n1228), .Z(n742) );
  BUF_X1 U194 ( .A(n1228), .Z(n743) );
  BUF_X1 U195 ( .A(n1228), .Z(n744) );
  BUF_X1 U196 ( .A(n1228), .Z(n745) );
  BUF_X1 U197 ( .A(n1228), .Z(n746) );
  BUF_X1 U198 ( .A(n1228), .Z(n747) );
  BUF_X1 U199 ( .A(n1261), .Z(n733) );
  BUF_X1 U200 ( .A(n1261), .Z(n734) );
  BUF_X1 U201 ( .A(n1261), .Z(n735) );
  BUF_X1 U202 ( .A(n1261), .Z(n736) );
  BUF_X1 U203 ( .A(n1261), .Z(n737) );
  BUF_X1 U204 ( .A(n1261), .Z(n738) );
  BUF_X1 U205 ( .A(n1295), .Z(n724) );
  BUF_X1 U206 ( .A(n1295), .Z(n725) );
  BUF_X1 U207 ( .A(n1295), .Z(n726) );
  BUF_X1 U208 ( .A(n1295), .Z(n727) );
  BUF_X1 U209 ( .A(n1295), .Z(n728) );
  BUF_X1 U210 ( .A(n1295), .Z(n729) );
  BUF_X1 U211 ( .A(n1329), .Z(n715) );
  BUF_X1 U212 ( .A(n1329), .Z(n716) );
  BUF_X1 U213 ( .A(n1329), .Z(n717) );
  BUF_X1 U214 ( .A(n1329), .Z(n718) );
  BUF_X1 U215 ( .A(n1329), .Z(n719) );
  BUF_X1 U216 ( .A(n1329), .Z(n720) );
  BUF_X1 U217 ( .A(n1364), .Z(n688) );
  BUF_X1 U218 ( .A(n1364), .Z(n689) );
  BUF_X1 U219 ( .A(n1364), .Z(n690) );
  BUF_X1 U220 ( .A(n1364), .Z(n691) );
  BUF_X1 U221 ( .A(n1364), .Z(n692) );
  BUF_X1 U222 ( .A(n1364), .Z(n693) );
  BUF_X1 U223 ( .A(n1397), .Z(n679) );
  BUF_X1 U224 ( .A(n1397), .Z(n680) );
  BUF_X1 U225 ( .A(n1397), .Z(n681) );
  BUF_X1 U226 ( .A(n1397), .Z(n682) );
  BUF_X1 U227 ( .A(n1397), .Z(n683) );
  BUF_X1 U228 ( .A(n1397), .Z(n684) );
  BUF_X1 U229 ( .A(n1435), .Z(n570) );
  BUF_X1 U230 ( .A(n1435), .Z(n571) );
  BUF_X1 U231 ( .A(n1435), .Z(n572) );
  BUF_X1 U232 ( .A(n1435), .Z(n573) );
  BUF_X1 U233 ( .A(n1435), .Z(n574) );
  BUF_X1 U234 ( .A(n1435), .Z(n575) );
  BUF_X1 U235 ( .A(n1468), .Z(n561) );
  BUF_X1 U236 ( .A(n1468), .Z(n562) );
  BUF_X1 U237 ( .A(n1468), .Z(n563) );
  BUF_X1 U238 ( .A(n1468), .Z(n564) );
  BUF_X1 U239 ( .A(n1468), .Z(n565) );
  BUF_X1 U240 ( .A(n1468), .Z(n566) );
  BUF_X1 U241 ( .A(n1503), .Z(n406) );
  BUF_X1 U242 ( .A(n1503), .Z(n407) );
  BUF_X1 U243 ( .A(n1503), .Z(n408) );
  BUF_X1 U244 ( .A(n1503), .Z(n409) );
  BUF_X1 U245 ( .A(n1503), .Z(n410) );
  BUF_X1 U246 ( .A(n1503), .Z(n411) );
  BUF_X1 U247 ( .A(n1536), .Z(n397) );
  BUF_X1 U248 ( .A(n1536), .Z(n398) );
  BUF_X1 U249 ( .A(n1536), .Z(n399) );
  BUF_X1 U250 ( .A(n1536), .Z(n400) );
  BUF_X1 U251 ( .A(n1536), .Z(n401) );
  BUF_X1 U252 ( .A(n1536), .Z(n402) );
  BUF_X1 U253 ( .A(n1), .Z(n911) );
  BUF_X1 U254 ( .A(n2), .Z(n902) );
  BUF_X1 U255 ( .A(n3), .Z(n893) );
  BUF_X1 U256 ( .A(n4), .Z(n884) );
  BUF_X1 U257 ( .A(n5), .Z(n866) );
  BUF_X1 U258 ( .A(n6), .Z(n793) );
  BUF_X1 U259 ( .A(n7), .Z(n766) );
  BUF_X1 U260 ( .A(n8), .Z(n757) );
  BUF_X1 U261 ( .A(n9), .Z(n712) );
  BUF_X1 U262 ( .A(n10), .Z(n703) );
  BUF_X1 U263 ( .A(n11), .Z(n676) );
  BUF_X1 U264 ( .A(n12), .Z(n594) );
  BUF_X1 U265 ( .A(n13), .Z(n585) );
  BUF_X1 U266 ( .A(n14), .Z(n558) );
  BUF_X1 U267 ( .A(n15), .Z(n549) );
  BUF_X1 U268 ( .A(n16), .Z(n603) );
  BUF_X1 U269 ( .A(n1078), .Z(n920) );
  BUF_X1 U270 ( .A(n1121), .Z(n875) );
  BUF_X1 U271 ( .A(n1160), .Z(n784) );
  BUF_X1 U272 ( .A(n1193), .Z(n775) );
  BUF_X1 U273 ( .A(n1228), .Z(n748) );
  BUF_X1 U274 ( .A(n1261), .Z(n739) );
  BUF_X1 U275 ( .A(n1295), .Z(n730) );
  BUF_X1 U276 ( .A(n1329), .Z(n721) );
  BUF_X1 U277 ( .A(n1364), .Z(n694) );
  BUF_X1 U278 ( .A(n1397), .Z(n685) );
  BUF_X1 U279 ( .A(n1435), .Z(n576) );
  BUF_X1 U280 ( .A(n1468), .Z(n567) );
  BUF_X1 U281 ( .A(n1503), .Z(n412) );
  BUF_X1 U282 ( .A(n1536), .Z(n403) );
  BUF_X1 U283 ( .A(n1009), .Z(n3321) );
  BUF_X1 U284 ( .A(n1009), .Z(n3320) );
  BUF_X1 U285 ( .A(n1008), .Z(n3319) );
  BUF_X1 U286 ( .A(n1008), .Z(n3318) );
  BUF_X1 U287 ( .A(n1007), .Z(n3317) );
  BUF_X1 U288 ( .A(n1007), .Z(n3316) );
  BUF_X1 U289 ( .A(n1006), .Z(n3315) );
  BUF_X1 U290 ( .A(n1006), .Z(n3314) );
  BUF_X1 U291 ( .A(n1005), .Z(n3313) );
  BUF_X1 U292 ( .A(n1005), .Z(n3312) );
  BUF_X1 U293 ( .A(n1004), .Z(n3311) );
  BUF_X1 U294 ( .A(n1004), .Z(n3310) );
  BUF_X1 U295 ( .A(n1003), .Z(n3309) );
  BUF_X1 U296 ( .A(n1003), .Z(n3308) );
  BUF_X1 U297 ( .A(n1002), .Z(n3307) );
  BUF_X1 U298 ( .A(n1002), .Z(n3306) );
  NOR3_X1 U299 ( .A1(n3805), .A2(n3806), .A3(n3804), .ZN(n1157) );
  BUF_X1 U300 ( .A(n1629), .Z(n259) );
  BUF_X1 U301 ( .A(n1634), .Z(n247) );
  BUF_X1 U302 ( .A(n1629), .Z(n260) );
  BUF_X1 U303 ( .A(n1634), .Z(n248) );
  BUF_X1 U304 ( .A(n2225), .Z(n26) );
  BUF_X1 U305 ( .A(n2220), .Z(n166) );
  BUF_X1 U306 ( .A(n2225), .Z(n27) );
  BUF_X1 U307 ( .A(n2220), .Z(n167) );
  BUF_X1 U308 ( .A(n1619), .Z(n280) );
  BUF_X1 U309 ( .A(n1619), .Z(n281) );
  BUF_X1 U310 ( .A(n2210), .Z(n187) );
  BUF_X1 U311 ( .A(n2210), .Z(n188) );
  BUF_X1 U312 ( .A(n1602), .Z(n386) );
  BUF_X1 U313 ( .A(n1607), .Z(n374) );
  BUF_X1 U314 ( .A(n1612), .Z(n362) );
  BUF_X1 U315 ( .A(n1617), .Z(n286) );
  BUF_X1 U316 ( .A(n1627), .Z(n265) );
  BUF_X1 U317 ( .A(n1602), .Z(n387) );
  BUF_X1 U318 ( .A(n1607), .Z(n375) );
  BUF_X1 U319 ( .A(n1612), .Z(n363) );
  BUF_X1 U320 ( .A(n1617), .Z(n287) );
  BUF_X1 U321 ( .A(n1627), .Z(n266) );
  BUF_X1 U322 ( .A(n2193), .Z(n229) );
  BUF_X1 U323 ( .A(n2198), .Z(n217) );
  BUF_X1 U324 ( .A(n2203), .Z(n205) );
  BUF_X1 U325 ( .A(n2208), .Z(n193) );
  BUF_X1 U326 ( .A(n2218), .Z(n172) );
  BUF_X1 U327 ( .A(n2193), .Z(n230) );
  BUF_X1 U328 ( .A(n2198), .Z(n218) );
  BUF_X1 U329 ( .A(n2203), .Z(n206) );
  BUF_X1 U330 ( .A(n2208), .Z(n194) );
  BUF_X1 U331 ( .A(n2218), .Z(n173) );
  BUF_X1 U332 ( .A(n1630), .Z(n256) );
  BUF_X1 U333 ( .A(n1635), .Z(n244) );
  BUF_X1 U334 ( .A(n1630), .Z(n257) );
  BUF_X1 U335 ( .A(n1635), .Z(n245) );
  BUF_X1 U336 ( .A(n2226), .Z(n23) );
  BUF_X1 U337 ( .A(n2221), .Z(n163) );
  BUF_X1 U338 ( .A(n2226), .Z(n24) );
  BUF_X1 U339 ( .A(n2221), .Z(n164) );
  BUF_X1 U340 ( .A(n1599), .Z(n392) );
  BUF_X1 U341 ( .A(n1604), .Z(n380) );
  BUF_X1 U342 ( .A(n1609), .Z(n368) );
  BUF_X1 U343 ( .A(n1614), .Z(n356) );
  BUF_X1 U344 ( .A(n1624), .Z(n271) );
  BUF_X1 U345 ( .A(n2190), .Z(n235) );
  BUF_X1 U346 ( .A(n2195), .Z(n223) );
  BUF_X1 U347 ( .A(n2200), .Z(n211) );
  BUF_X1 U348 ( .A(n2205), .Z(n199) );
  BUF_X1 U349 ( .A(n2215), .Z(n178) );
  BUF_X1 U350 ( .A(n1603), .Z(n383) );
  BUF_X1 U351 ( .A(n1608), .Z(n371) );
  BUF_X1 U352 ( .A(n1613), .Z(n359) );
  BUF_X1 U353 ( .A(n1618), .Z(n283) );
  BUF_X1 U354 ( .A(n1628), .Z(n262) );
  BUF_X1 U355 ( .A(n1603), .Z(n384) );
  BUF_X1 U356 ( .A(n1608), .Z(n372) );
  BUF_X1 U357 ( .A(n1613), .Z(n360) );
  BUF_X1 U358 ( .A(n1618), .Z(n284) );
  BUF_X1 U359 ( .A(n1628), .Z(n263) );
  BUF_X1 U360 ( .A(n2194), .Z(n226) );
  BUF_X1 U361 ( .A(n2199), .Z(n214) );
  BUF_X1 U362 ( .A(n2204), .Z(n202) );
  BUF_X1 U363 ( .A(n2209), .Z(n190) );
  BUF_X1 U364 ( .A(n2219), .Z(n169) );
  BUF_X1 U365 ( .A(n2194), .Z(n227) );
  BUF_X1 U366 ( .A(n2199), .Z(n215) );
  BUF_X1 U367 ( .A(n2204), .Z(n203) );
  BUF_X1 U368 ( .A(n2209), .Z(n191) );
  BUF_X1 U369 ( .A(n2219), .Z(n170) );
  BUF_X1 U370 ( .A(n1600), .Z(n391) );
  BUF_X1 U371 ( .A(n1605), .Z(n379) );
  BUF_X1 U372 ( .A(n1610), .Z(n367) );
  BUF_X1 U373 ( .A(n1615), .Z(n355) );
  BUF_X1 U374 ( .A(n1625), .Z(n270) );
  BUF_X1 U375 ( .A(n2191), .Z(n234) );
  BUF_X1 U376 ( .A(n2196), .Z(n222) );
  BUF_X1 U377 ( .A(n2201), .Z(n210) );
  BUF_X1 U378 ( .A(n2206), .Z(n198) );
  BUF_X1 U379 ( .A(n2216), .Z(n177) );
  BUF_X1 U380 ( .A(n1634), .Z(n249) );
  BUF_X1 U381 ( .A(n1629), .Z(n261) );
  BUF_X1 U382 ( .A(n2225), .Z(n28) );
  BUF_X1 U383 ( .A(n2220), .Z(n168) );
  BUF_X1 U384 ( .A(n1619), .Z(n282) );
  BUF_X1 U385 ( .A(n2210), .Z(n189) );
  BUF_X1 U386 ( .A(n1602), .Z(n388) );
  BUF_X1 U387 ( .A(n1607), .Z(n376) );
  BUF_X1 U388 ( .A(n1612), .Z(n364) );
  BUF_X1 U389 ( .A(n1617), .Z(n288) );
  BUF_X1 U390 ( .A(n1627), .Z(n267) );
  BUF_X1 U391 ( .A(n2193), .Z(n231) );
  BUF_X1 U392 ( .A(n2198), .Z(n219) );
  BUF_X1 U393 ( .A(n2203), .Z(n207) );
  BUF_X1 U394 ( .A(n2208), .Z(n195) );
  BUF_X1 U395 ( .A(n2218), .Z(n174) );
  BUF_X1 U396 ( .A(n1635), .Z(n246) );
  BUF_X1 U397 ( .A(n1630), .Z(n258) );
  BUF_X1 U398 ( .A(n2226), .Z(n25) );
  BUF_X1 U399 ( .A(n2221), .Z(n165) );
  BUF_X1 U400 ( .A(n1599), .Z(n394) );
  BUF_X1 U401 ( .A(n1604), .Z(n382) );
  BUF_X1 U402 ( .A(n1609), .Z(n370) );
  BUF_X1 U403 ( .A(n1614), .Z(n358) );
  BUF_X1 U404 ( .A(n1624), .Z(n273) );
  BUF_X1 U405 ( .A(n2190), .Z(n237) );
  BUF_X1 U406 ( .A(n2195), .Z(n225) );
  BUF_X1 U407 ( .A(n2200), .Z(n213) );
  BUF_X1 U408 ( .A(n2205), .Z(n201) );
  BUF_X1 U409 ( .A(n2215), .Z(n180) );
  BUF_X1 U410 ( .A(n1603), .Z(n385) );
  BUF_X1 U411 ( .A(n1608), .Z(n373) );
  BUF_X1 U412 ( .A(n1613), .Z(n361) );
  BUF_X1 U413 ( .A(n1618), .Z(n285) );
  BUF_X1 U414 ( .A(n1628), .Z(n264) );
  BUF_X1 U415 ( .A(n2194), .Z(n228) );
  BUF_X1 U416 ( .A(n2199), .Z(n216) );
  BUF_X1 U417 ( .A(n2204), .Z(n204) );
  BUF_X1 U418 ( .A(n2209), .Z(n192) );
  BUF_X1 U419 ( .A(n2219), .Z(n171) );
  BUF_X1 U420 ( .A(n1622), .Z(n277) );
  BUF_X1 U421 ( .A(n1637), .Z(n241) );
  BUF_X1 U422 ( .A(n1622), .Z(n278) );
  BUF_X1 U423 ( .A(n1637), .Z(n242) );
  BUF_X1 U424 ( .A(n2213), .Z(n184) );
  BUF_X1 U425 ( .A(n2228), .Z(n20) );
  BUF_X1 U426 ( .A(n2213), .Z(n185) );
  BUF_X1 U427 ( .A(n2228), .Z(n21) );
  BUF_X1 U428 ( .A(n1632), .Z(n253) );
  BUF_X1 U429 ( .A(n1632), .Z(n254) );
  BUF_X1 U430 ( .A(n2223), .Z(n32) );
  BUF_X1 U431 ( .A(n2223), .Z(n161) );
  BUF_X1 U432 ( .A(n1623), .Z(n274) );
  BUF_X1 U433 ( .A(n1638), .Z(n238) );
  BUF_X1 U434 ( .A(n1623), .Z(n275) );
  BUF_X1 U435 ( .A(n1638), .Z(n239) );
  BUF_X1 U436 ( .A(n2214), .Z(n181) );
  BUF_X1 U437 ( .A(n2229), .Z(n17) );
  BUF_X1 U438 ( .A(n2214), .Z(n182) );
  BUF_X1 U439 ( .A(n2229), .Z(n18) );
  BUF_X1 U440 ( .A(n1633), .Z(n250) );
  BUF_X1 U441 ( .A(n1633), .Z(n251) );
  BUF_X1 U442 ( .A(n2224), .Z(n29) );
  BUF_X1 U443 ( .A(n2224), .Z(n30) );
  BUF_X1 U444 ( .A(n1622), .Z(n279) );
  BUF_X1 U445 ( .A(n1637), .Z(n243) );
  BUF_X1 U446 ( .A(n2213), .Z(n186) );
  BUF_X1 U447 ( .A(n2228), .Z(n22) );
  BUF_X1 U448 ( .A(n1632), .Z(n255) );
  BUF_X1 U449 ( .A(n2223), .Z(n162) );
  NAND2_X1 U450 ( .A1(n1157), .A2(n1111), .ZN(n1068) );
  NAND2_X1 U451 ( .A1(n1110), .A2(n1111), .ZN(n1078) );
  NAND2_X1 U452 ( .A1(n1153), .A2(n1111), .ZN(n1121) );
  BUF_X1 U453 ( .A(n1623), .Z(n276) );
  BUF_X1 U454 ( .A(n1638), .Z(n240) );
  BUF_X1 U455 ( .A(n2214), .Z(n183) );
  BUF_X1 U456 ( .A(n2229), .Z(n19) );
  BUF_X1 U457 ( .A(n1633), .Z(n252) );
  BUF_X1 U458 ( .A(n2224), .Z(n31) );
  BUF_X1 U459 ( .A(n1600), .Z(n389) );
  BUF_X1 U460 ( .A(n1605), .Z(n377) );
  BUF_X1 U461 ( .A(n1610), .Z(n365) );
  BUF_X1 U462 ( .A(n1615), .Z(n353) );
  BUF_X1 U463 ( .A(n1625), .Z(n268) );
  BUF_X1 U464 ( .A(n1600), .Z(n390) );
  BUF_X1 U465 ( .A(n1605), .Z(n378) );
  BUF_X1 U466 ( .A(n1610), .Z(n366) );
  BUF_X1 U467 ( .A(n1615), .Z(n354) );
  BUF_X1 U468 ( .A(n1625), .Z(n269) );
  BUF_X1 U469 ( .A(n2191), .Z(n232) );
  BUF_X1 U470 ( .A(n2196), .Z(n220) );
  BUF_X1 U471 ( .A(n2201), .Z(n208) );
  BUF_X1 U472 ( .A(n2206), .Z(n196) );
  BUF_X1 U473 ( .A(n2216), .Z(n175) );
  BUF_X1 U474 ( .A(n2191), .Z(n233) );
  BUF_X1 U475 ( .A(n2196), .Z(n221) );
  BUF_X1 U476 ( .A(n2201), .Z(n209) );
  BUF_X1 U477 ( .A(n2206), .Z(n197) );
  BUF_X1 U478 ( .A(n2216), .Z(n176) );
  BUF_X1 U479 ( .A(n1599), .Z(n393) );
  BUF_X1 U480 ( .A(n1604), .Z(n381) );
  BUF_X1 U481 ( .A(n1609), .Z(n369) );
  BUF_X1 U482 ( .A(n1614), .Z(n357) );
  BUF_X1 U483 ( .A(n1624), .Z(n272) );
  BUF_X1 U484 ( .A(n2190), .Z(n236) );
  BUF_X1 U485 ( .A(n2195), .Z(n224) );
  BUF_X1 U486 ( .A(n2200), .Z(n212) );
  BUF_X1 U487 ( .A(n2205), .Z(n200) );
  BUF_X1 U488 ( .A(n2215), .Z(n179) );
  NAND2_X1 U489 ( .A1(n1156), .A2(n1113), .ZN(n1160) );
  NAND2_X1 U490 ( .A1(n1156), .A2(n1115), .ZN(n1193) );
  NAND2_X1 U491 ( .A1(n1156), .A2(n1153), .ZN(n1228) );
  NAND2_X1 U492 ( .A1(n1327), .A2(n1157), .ZN(n1295) );
  NAND2_X1 U493 ( .A1(n1327), .A2(n1110), .ZN(n1329) );
  NAND2_X1 U494 ( .A1(n1327), .A2(n1117), .ZN(n1364) );
  NAND2_X1 U495 ( .A1(n1327), .A2(n1119), .ZN(n1397) );
  NAND2_X1 U496 ( .A1(n1432), .A2(n1113), .ZN(n1435) );
  NAND2_X1 U497 ( .A1(n1432), .A2(n1115), .ZN(n1468) );
  NAND2_X1 U498 ( .A1(n1432), .A2(n1153), .ZN(n1503) );
  NAND2_X1 U499 ( .A1(n1156), .A2(n1154), .ZN(n1261) );
  NAND2_X1 U500 ( .A1(n1432), .A2(n1154), .ZN(n1536) );
  AND2_X1 U501 ( .A1(n1113), .A2(n1111), .ZN(n1) );
  AND2_X1 U502 ( .A1(n1115), .A2(n1111), .ZN(n2) );
  AND2_X1 U503 ( .A1(n1117), .A2(n1111), .ZN(n3) );
  AND2_X1 U504 ( .A1(n1119), .A2(n1111), .ZN(n4) );
  AND2_X1 U505 ( .A1(n1156), .A2(n1157), .ZN(n5) );
  AND2_X1 U506 ( .A1(n1156), .A2(n1110), .ZN(n6) );
  AND2_X1 U507 ( .A1(n1156), .A2(n1117), .ZN(n7) );
  AND2_X1 U508 ( .A1(n1156), .A2(n1119), .ZN(n8) );
  AND2_X1 U509 ( .A1(n1327), .A2(n1113), .ZN(n9) );
  AND2_X1 U510 ( .A1(n1327), .A2(n1115), .ZN(n10) );
  AND2_X1 U511 ( .A1(n1327), .A2(n1153), .ZN(n11) );
  AND2_X1 U512 ( .A1(n1432), .A2(n1157), .ZN(n12) );
  AND2_X1 U513 ( .A1(n1432), .A2(n1110), .ZN(n13) );
  AND2_X1 U514 ( .A1(n1432), .A2(n1117), .ZN(n14) );
  AND2_X1 U515 ( .A1(n1432), .A2(n1119), .ZN(n15) );
  AND2_X1 U516 ( .A1(n1327), .A2(n1154), .ZN(n16) );
  BUF_X1 U517 ( .A(n1010), .Z(n1009) );
  BUF_X1 U518 ( .A(n1010), .Z(n1008) );
  BUF_X1 U519 ( .A(n1010), .Z(n1007) );
  BUF_X1 U520 ( .A(n1011), .Z(n1006) );
  BUF_X1 U521 ( .A(n1011), .Z(n1005) );
  BUF_X1 U522 ( .A(n1011), .Z(n1004) );
  BUF_X1 U523 ( .A(n1012), .Z(n1003) );
  BUF_X1 U524 ( .A(n1012), .Z(n1002) );
  INV_X1 U525 ( .A(DATAIN[0]), .ZN(n3844) );
  INV_X1 U526 ( .A(DATAIN[1]), .ZN(n3843) );
  INV_X1 U527 ( .A(DATAIN[2]), .ZN(n3842) );
  INV_X1 U528 ( .A(DATAIN[3]), .ZN(n3841) );
  INV_X1 U529 ( .A(DATAIN[4]), .ZN(n3840) );
  INV_X1 U530 ( .A(DATAIN[5]), .ZN(n3839) );
  INV_X1 U531 ( .A(DATAIN[6]), .ZN(n3838) );
  INV_X1 U532 ( .A(DATAIN[7]), .ZN(n3837) );
  INV_X1 U533 ( .A(DATAIN[8]), .ZN(n3836) );
  INV_X1 U534 ( .A(DATAIN[9]), .ZN(n3835) );
  INV_X1 U535 ( .A(DATAIN[10]), .ZN(n3834) );
  INV_X1 U536 ( .A(DATAIN[11]), .ZN(n3833) );
  INV_X1 U537 ( .A(DATAIN[12]), .ZN(n3832) );
  INV_X1 U538 ( .A(DATAIN[13]), .ZN(n3831) );
  INV_X1 U539 ( .A(DATAIN[14]), .ZN(n3830) );
  INV_X1 U540 ( .A(DATAIN[15]), .ZN(n3829) );
  INV_X1 U541 ( .A(DATAIN[16]), .ZN(n3828) );
  INV_X1 U542 ( .A(DATAIN[17]), .ZN(n3827) );
  INV_X1 U543 ( .A(DATAIN[18]), .ZN(n3826) );
  INV_X1 U544 ( .A(DATAIN[19]), .ZN(n3825) );
  INV_X1 U545 ( .A(DATAIN[20]), .ZN(n3824) );
  INV_X1 U546 ( .A(DATAIN[21]), .ZN(n3823) );
  INV_X1 U547 ( .A(DATAIN[22]), .ZN(n3822) );
  INV_X1 U548 ( .A(DATAIN[23]), .ZN(n3821) );
  INV_X1 U549 ( .A(DATAIN[24]), .ZN(n3820) );
  INV_X1 U550 ( .A(DATAIN[25]), .ZN(n3819) );
  INV_X1 U551 ( .A(DATAIN[26]), .ZN(n3818) );
  INV_X1 U552 ( .A(DATAIN[27]), .ZN(n3817) );
  INV_X1 U553 ( .A(DATAIN[28]), .ZN(n3816) );
  INV_X1 U554 ( .A(DATAIN[29]), .ZN(n3815) );
  INV_X1 U555 ( .A(DATAIN[30]), .ZN(n3814) );
  INV_X1 U556 ( .A(DATAIN[31]), .ZN(n3813) );
  NOR3_X1 U557 ( .A1(n3806), .A2(ADD_WR[1]), .A3(n3804), .ZN(n1113) );
  NOR3_X1 U558 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n3804), .ZN(n1115) );
  NOR3_X1 U559 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n3806), .ZN(n1153) );
  NOR3_X1 U560 ( .A1(n3805), .A2(ADD_WR[0]), .A3(n3804), .ZN(n1110) );
  NOR3_X1 U561 ( .A1(n3806), .A2(ADD_WR[2]), .A3(n3805), .ZN(n1117) );
  NOR3_X1 U562 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n3805), .ZN(n1119) );
  NOR3_X1 U563 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n1154) );
  AND3_X1 U564 ( .A1(ADD_WR[3]), .A2(n1293), .A3(ADD_WR[4]), .ZN(n1156) );
  AND3_X1 U565 ( .A1(n1293), .A2(n3546), .A3(ADD_WR[3]), .ZN(n1432) );
  AND3_X1 U566 ( .A1(n1293), .A2(n3803), .A3(ADD_WR[4]), .ZN(n1327) );
  AND3_X1 U567 ( .A1(n3803), .A2(n3546), .A3(n1293), .ZN(n1111) );
  NAND2_X1 U568 ( .A1(n2159), .A2(n2167), .ZN(n1610) );
  NAND2_X1 U569 ( .A1(n2750), .A2(n2758), .ZN(n2201) );
  NAND2_X1 U570 ( .A1(n2159), .A2(n2168), .ZN(n1609) );
  NAND2_X1 U571 ( .A1(n2750), .A2(n2759), .ZN(n2200) );
  INV_X1 U572 ( .A(ADD_WR[2]), .ZN(n3804) );
  INV_X1 U573 ( .A(ADD_WR[1]), .ZN(n3805) );
  INV_X1 U574 ( .A(ADD_WR[0]), .ZN(n3806) );
  NAND2_X1 U575 ( .A1(n2173), .A2(n2159), .ZN(n1623) );
  NAND2_X1 U576 ( .A1(n2174), .A2(n2159), .ZN(n1622) );
  NAND2_X1 U577 ( .A1(n2178), .A2(n2159), .ZN(n1638) );
  NAND2_X1 U578 ( .A1(n2179), .A2(n2159), .ZN(n1637) );
  NAND2_X1 U579 ( .A1(n2764), .A2(n2750), .ZN(n2214) );
  NAND2_X1 U580 ( .A1(n2765), .A2(n2750), .ZN(n2213) );
  NAND2_X1 U581 ( .A1(n2769), .A2(n2750), .ZN(n2229) );
  NAND2_X1 U582 ( .A1(n2770), .A2(n2750), .ZN(n2228) );
  AND2_X1 U583 ( .A1(n2170), .A2(n3812), .ZN(n2167) );
  AND2_X1 U584 ( .A1(n2761), .A2(n3809), .ZN(n2758) );
  NAND2_X1 U585 ( .A1(n2158), .A2(n2161), .ZN(n1600) );
  AND2_X1 U586 ( .A1(n2181), .A2(n3812), .ZN(n2179) );
  AND2_X1 U587 ( .A1(n2772), .A2(n3809), .ZN(n2770) );
  AND2_X1 U588 ( .A1(n2165), .A2(n3812), .ZN(n2158) );
  AND2_X1 U589 ( .A1(n2756), .A2(n3809), .ZN(n2749) );
  NAND2_X1 U590 ( .A1(n2749), .A2(n2752), .ZN(n2191) );
  NAND2_X1 U591 ( .A1(n2158), .A2(n2164), .ZN(n1605) );
  NAND2_X1 U592 ( .A1(n2174), .A2(n2164), .ZN(n1625) );
  NAND2_X1 U593 ( .A1(n2749), .A2(n2755), .ZN(n2196) );
  NAND2_X1 U594 ( .A1(n2765), .A2(n2755), .ZN(n2216) );
  NAND2_X1 U595 ( .A1(n2167), .A2(n2163), .ZN(n1615) );
  NAND2_X1 U596 ( .A1(n2179), .A2(n2163), .ZN(n1632) );
  NAND2_X1 U597 ( .A1(n2178), .A2(n2163), .ZN(n1633) );
  NAND2_X1 U598 ( .A1(n2758), .A2(n2754), .ZN(n2206) );
  NAND2_X1 U599 ( .A1(n2770), .A2(n2754), .ZN(n2223) );
  NAND2_X1 U600 ( .A1(n2769), .A2(n2754), .ZN(n2224) );
  NAND2_X1 U601 ( .A1(n2160), .A2(n2161), .ZN(n1599) );
  NAND2_X1 U602 ( .A1(n2751), .A2(n2752), .ZN(n2190) );
  NAND2_X1 U603 ( .A1(n2163), .A2(n2168), .ZN(n1614) );
  NAND2_X1 U604 ( .A1(n2754), .A2(n2759), .ZN(n2205) );
  AND2_X1 U605 ( .A1(n2176), .A2(n3812), .ZN(n2174) );
  AND2_X1 U606 ( .A1(n2767), .A2(n3809), .ZN(n2765) );
  NAND2_X1 U607 ( .A1(n2160), .A2(n2164), .ZN(n1604) );
  NAND2_X1 U608 ( .A1(n2173), .A2(n2164), .ZN(n1624) );
  NAND2_X1 U609 ( .A1(n2751), .A2(n2755), .ZN(n2195) );
  NAND2_X1 U610 ( .A1(n2764), .A2(n2755), .ZN(n2215) );
  AND2_X1 U611 ( .A1(n2158), .A2(n2159), .ZN(n1603) );
  AND2_X1 U612 ( .A1(n2160), .A2(n2159), .ZN(n1602) );
  AND2_X1 U613 ( .A1(n2749), .A2(n2750), .ZN(n2194) );
  AND2_X1 U614 ( .A1(n2751), .A2(n2750), .ZN(n2193) );
  AND2_X1 U615 ( .A1(n2161), .A2(n2167), .ZN(n1613) );
  AND2_X1 U616 ( .A1(n2161), .A2(n2168), .ZN(n1612) );
  AND2_X1 U617 ( .A1(n2752), .A2(n2758), .ZN(n2204) );
  AND2_X1 U618 ( .A1(n2752), .A2(n2759), .ZN(n2203) );
  AND2_X1 U619 ( .A1(n2173), .A2(n2161), .ZN(n1619) );
  AND2_X1 U620 ( .A1(n2178), .A2(n2161), .ZN(n1634) );
  AND2_X1 U621 ( .A1(n2179), .A2(n2161), .ZN(n1635) );
  AND2_X1 U622 ( .A1(n2764), .A2(n2752), .ZN(n2210) );
  AND2_X1 U623 ( .A1(n2769), .A2(n2752), .ZN(n2225) );
  AND2_X1 U624 ( .A1(n2770), .A2(n2752), .ZN(n2226) );
  AND2_X1 U625 ( .A1(n2164), .A2(n2167), .ZN(n1618) );
  AND2_X1 U626 ( .A1(n2164), .A2(n2168), .ZN(n1617) );
  AND2_X1 U627 ( .A1(n2755), .A2(n2758), .ZN(n2209) );
  AND2_X1 U628 ( .A1(n2755), .A2(n2759), .ZN(n2208) );
  AND2_X1 U629 ( .A1(n2178), .A2(n2164), .ZN(n1629) );
  AND2_X1 U630 ( .A1(n2179), .A2(n2164), .ZN(n1630) );
  AND2_X1 U631 ( .A1(n2769), .A2(n2755), .ZN(n2220) );
  AND2_X1 U632 ( .A1(n2770), .A2(n2755), .ZN(n2221) );
  AND2_X1 U633 ( .A1(n2158), .A2(n2163), .ZN(n1608) );
  AND2_X1 U634 ( .A1(n2160), .A2(n2163), .ZN(n1607) );
  AND2_X1 U635 ( .A1(n2174), .A2(n2163), .ZN(n1628) );
  AND2_X1 U636 ( .A1(n2173), .A2(n2163), .ZN(n1627) );
  AND2_X1 U637 ( .A1(n2749), .A2(n2754), .ZN(n2199) );
  AND2_X1 U638 ( .A1(n2751), .A2(n2754), .ZN(n2198) );
  AND2_X1 U639 ( .A1(n2765), .A2(n2754), .ZN(n2219) );
  AND2_X1 U640 ( .A1(n2764), .A2(n2754), .ZN(n2218) );
  INV_X1 U641 ( .A(ADD_WR[4]), .ZN(n3546) );
  INV_X1 U642 ( .A(ADD_WR[3]), .ZN(n3803) );
  BUF_X1 U643 ( .A(RST_AN), .Z(n1010) );
  BUF_X1 U644 ( .A(RST_AN), .Z(n1011) );
  BUF_X1 U645 ( .A(RST_AN), .Z(n1012) );
  NOR2_X1 U646 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n2161) );
  NOR2_X1 U647 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2752) );
  NOR4_X1 U648 ( .A1(n1779), .A2(n1780), .A3(n1781), .A4(n1782), .ZN(n1778) );
  OAI221_X1 U649 ( .B1(n970), .B2(n358), .C1(n938), .C2(n355), .A(n1786), .ZN(
        n1779) );
  OAI221_X1 U650 ( .B1(n842), .B2(n370), .C1(n810), .C2(n367), .A(n1785), .ZN(
        n1780) );
  OAI221_X1 U651 ( .B1(n650), .B2(n382), .C1(n618), .C2(n379), .A(n1784), .ZN(
        n1781) );
  NOR4_X1 U652 ( .A1(n1762), .A2(n1763), .A3(n1764), .A4(n1765), .ZN(n1761) );
  OAI221_X1 U653 ( .B1(n969), .B2(n358), .C1(n937), .C2(n355), .A(n1769), .ZN(
        n1762) );
  OAI221_X1 U654 ( .B1(n841), .B2(n370), .C1(n809), .C2(n367), .A(n1768), .ZN(
        n1763) );
  OAI221_X1 U655 ( .B1(n649), .B2(n382), .C1(n617), .C2(n379), .A(n1767), .ZN(
        n1764) );
  NOR4_X1 U656 ( .A1(n1745), .A2(n1746), .A3(n1747), .A4(n1748), .ZN(n1744) );
  OAI221_X1 U657 ( .B1(n968), .B2(n358), .C1(n936), .C2(n355), .A(n1752), .ZN(
        n1745) );
  OAI221_X1 U658 ( .B1(n840), .B2(n370), .C1(n808), .C2(n367), .A(n1751), .ZN(
        n1746) );
  OAI221_X1 U659 ( .B1(n648), .B2(n382), .C1(n616), .C2(n379), .A(n1750), .ZN(
        n1747) );
  NOR4_X1 U660 ( .A1(n1728), .A2(n1729), .A3(n1730), .A4(n1731), .ZN(n1727) );
  OAI221_X1 U661 ( .B1(n967), .B2(n358), .C1(n935), .C2(n355), .A(n1735), .ZN(
        n1728) );
  OAI221_X1 U662 ( .B1(n839), .B2(n370), .C1(n807), .C2(n367), .A(n1734), .ZN(
        n1729) );
  OAI221_X1 U663 ( .B1(n647), .B2(n382), .C1(n615), .C2(n379), .A(n1733), .ZN(
        n1730) );
  NOR4_X1 U664 ( .A1(n1711), .A2(n1712), .A3(n1713), .A4(n1714), .ZN(n1710) );
  OAI221_X1 U665 ( .B1(n966), .B2(n358), .C1(n934), .C2(n355), .A(n1718), .ZN(
        n1711) );
  OAI221_X1 U666 ( .B1(n838), .B2(n370), .C1(n806), .C2(n367), .A(n1717), .ZN(
        n1712) );
  OAI221_X1 U667 ( .B1(n646), .B2(n382), .C1(n614), .C2(n379), .A(n1716), .ZN(
        n1713) );
  NOR4_X1 U668 ( .A1(n1694), .A2(n1695), .A3(n1696), .A4(n1697), .ZN(n1693) );
  OAI221_X1 U669 ( .B1(n965), .B2(n358), .C1(n933), .C2(n355), .A(n1701), .ZN(
        n1694) );
  OAI221_X1 U670 ( .B1(n837), .B2(n370), .C1(n805), .C2(n367), .A(n1700), .ZN(
        n1695) );
  OAI221_X1 U671 ( .B1(n645), .B2(n382), .C1(n613), .C2(n379), .A(n1699), .ZN(
        n1696) );
  NOR4_X1 U672 ( .A1(n1677), .A2(n1678), .A3(n1679), .A4(n1680), .ZN(n1676) );
  OAI221_X1 U673 ( .B1(n964), .B2(n358), .C1(n932), .C2(n355), .A(n1684), .ZN(
        n1677) );
  OAI221_X1 U674 ( .B1(n836), .B2(n370), .C1(n804), .C2(n367), .A(n1683), .ZN(
        n1678) );
  OAI221_X1 U675 ( .B1(n644), .B2(n382), .C1(n612), .C2(n379), .A(n1682), .ZN(
        n1679) );
  NOR4_X1 U676 ( .A1(n1660), .A2(n1661), .A3(n1662), .A4(n1663), .ZN(n1659) );
  OAI221_X1 U677 ( .B1(n963), .B2(n358), .C1(n931), .C2(n355), .A(n1667), .ZN(
        n1660) );
  OAI221_X1 U678 ( .B1(n835), .B2(n370), .C1(n803), .C2(n367), .A(n1666), .ZN(
        n1661) );
  OAI221_X1 U679 ( .B1(n643), .B2(n382), .C1(n611), .C2(n379), .A(n1665), .ZN(
        n1662) );
  NOR4_X1 U680 ( .A1(n1643), .A2(n1644), .A3(n1645), .A4(n1646), .ZN(n1642) );
  OAI221_X1 U681 ( .B1(n962), .B2(n358), .C1(n930), .C2(n355), .A(n1650), .ZN(
        n1643) );
  OAI221_X1 U682 ( .B1(n834), .B2(n370), .C1(n802), .C2(n367), .A(n1649), .ZN(
        n1644) );
  OAI221_X1 U683 ( .B1(n642), .B2(n382), .C1(n610), .C2(n379), .A(n1648), .ZN(
        n1645) );
  NOR4_X1 U684 ( .A1(n1595), .A2(n1596), .A3(n1597), .A4(n1598), .ZN(n1594) );
  OAI221_X1 U685 ( .B1(n961), .B2(n358), .C1(n929), .C2(n355), .A(n1616), .ZN(
        n1595) );
  OAI221_X1 U686 ( .B1(n833), .B2(n370), .C1(n801), .C2(n367), .A(n1611), .ZN(
        n1596) );
  OAI221_X1 U687 ( .B1(n641), .B2(n382), .C1(n609), .C2(n379), .A(n1606), .ZN(
        n1597) );
  NOR4_X1 U688 ( .A1(n2370), .A2(n2371), .A3(n2372), .A4(n2373), .ZN(n2369) );
  OAI221_X1 U689 ( .B1(n970), .B2(n201), .C1(n938), .C2(n198), .A(n2377), .ZN(
        n2370) );
  OAI221_X1 U690 ( .B1(n842), .B2(n213), .C1(n810), .C2(n210), .A(n2376), .ZN(
        n2371) );
  OAI221_X1 U691 ( .B1(n650), .B2(n225), .C1(n618), .C2(n222), .A(n2375), .ZN(
        n2372) );
  NOR4_X1 U692 ( .A1(n2353), .A2(n2354), .A3(n2355), .A4(n2356), .ZN(n2352) );
  OAI221_X1 U693 ( .B1(n969), .B2(n201), .C1(n937), .C2(n198), .A(n2360), .ZN(
        n2353) );
  OAI221_X1 U694 ( .B1(n841), .B2(n213), .C1(n809), .C2(n210), .A(n2359), .ZN(
        n2354) );
  OAI221_X1 U695 ( .B1(n649), .B2(n225), .C1(n617), .C2(n222), .A(n2358), .ZN(
        n2355) );
  NOR4_X1 U696 ( .A1(n2336), .A2(n2337), .A3(n2338), .A4(n2339), .ZN(n2335) );
  OAI221_X1 U697 ( .B1(n968), .B2(n201), .C1(n936), .C2(n198), .A(n2343), .ZN(
        n2336) );
  OAI221_X1 U698 ( .B1(n840), .B2(n213), .C1(n808), .C2(n210), .A(n2342), .ZN(
        n2337) );
  OAI221_X1 U699 ( .B1(n648), .B2(n225), .C1(n616), .C2(n222), .A(n2341), .ZN(
        n2338) );
  NOR4_X1 U700 ( .A1(n2319), .A2(n2320), .A3(n2321), .A4(n2322), .ZN(n2318) );
  OAI221_X1 U701 ( .B1(n967), .B2(n201), .C1(n935), .C2(n198), .A(n2326), .ZN(
        n2319) );
  OAI221_X1 U702 ( .B1(n839), .B2(n213), .C1(n807), .C2(n210), .A(n2325), .ZN(
        n2320) );
  OAI221_X1 U703 ( .B1(n647), .B2(n225), .C1(n615), .C2(n222), .A(n2324), .ZN(
        n2321) );
  NOR4_X1 U704 ( .A1(n2302), .A2(n2303), .A3(n2304), .A4(n2305), .ZN(n2301) );
  OAI221_X1 U705 ( .B1(n966), .B2(n201), .C1(n934), .C2(n198), .A(n2309), .ZN(
        n2302) );
  OAI221_X1 U706 ( .B1(n838), .B2(n213), .C1(n806), .C2(n210), .A(n2308), .ZN(
        n2303) );
  OAI221_X1 U707 ( .B1(n646), .B2(n225), .C1(n614), .C2(n222), .A(n2307), .ZN(
        n2304) );
  NOR4_X1 U708 ( .A1(n2285), .A2(n2286), .A3(n2287), .A4(n2288), .ZN(n2284) );
  OAI221_X1 U709 ( .B1(n965), .B2(n201), .C1(n933), .C2(n198), .A(n2292), .ZN(
        n2285) );
  OAI221_X1 U710 ( .B1(n837), .B2(n213), .C1(n805), .C2(n210), .A(n2291), .ZN(
        n2286) );
  OAI221_X1 U711 ( .B1(n645), .B2(n225), .C1(n613), .C2(n222), .A(n2290), .ZN(
        n2287) );
  NOR4_X1 U712 ( .A1(n2268), .A2(n2269), .A3(n2270), .A4(n2271), .ZN(n2267) );
  OAI221_X1 U713 ( .B1(n964), .B2(n201), .C1(n932), .C2(n198), .A(n2275), .ZN(
        n2268) );
  OAI221_X1 U714 ( .B1(n836), .B2(n213), .C1(n804), .C2(n210), .A(n2274), .ZN(
        n2269) );
  OAI221_X1 U715 ( .B1(n644), .B2(n225), .C1(n612), .C2(n222), .A(n2273), .ZN(
        n2270) );
  NOR4_X1 U716 ( .A1(n2251), .A2(n2252), .A3(n2253), .A4(n2254), .ZN(n2250) );
  OAI221_X1 U717 ( .B1(n963), .B2(n201), .C1(n931), .C2(n198), .A(n2258), .ZN(
        n2251) );
  OAI221_X1 U718 ( .B1(n835), .B2(n213), .C1(n803), .C2(n210), .A(n2257), .ZN(
        n2252) );
  OAI221_X1 U719 ( .B1(n643), .B2(n225), .C1(n611), .C2(n222), .A(n2256), .ZN(
        n2253) );
  NOR4_X1 U720 ( .A1(n2234), .A2(n2235), .A3(n2236), .A4(n2237), .ZN(n2233) );
  OAI221_X1 U721 ( .B1(n962), .B2(n201), .C1(n930), .C2(n198), .A(n2241), .ZN(
        n2234) );
  OAI221_X1 U722 ( .B1(n834), .B2(n213), .C1(n802), .C2(n210), .A(n2240), .ZN(
        n2235) );
  OAI221_X1 U723 ( .B1(n642), .B2(n225), .C1(n610), .C2(n222), .A(n2239), .ZN(
        n2236) );
  NOR4_X1 U724 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(n2185) );
  OAI221_X1 U725 ( .B1(n961), .B2(n201), .C1(n929), .C2(n198), .A(n2207), .ZN(
        n2186) );
  OAI221_X1 U726 ( .B1(n833), .B2(n213), .C1(n801), .C2(n210), .A(n2202), .ZN(
        n2187) );
  OAI221_X1 U727 ( .B1(n641), .B2(n225), .C1(n609), .C2(n222), .A(n2197), .ZN(
        n2188) );
  NOR4_X1 U728 ( .A1(n2153), .A2(n2154), .A3(n2155), .A4(n2156), .ZN(n2152) );
  OAI221_X1 U729 ( .B1(n992), .B2(n356), .C1(n960), .C2(n353), .A(n2169), .ZN(
        n2153) );
  OAI221_X1 U730 ( .B1(n864), .B2(n368), .C1(n832), .C2(n365), .A(n2166), .ZN(
        n2154) );
  OAI221_X1 U731 ( .B1(n672), .B2(n380), .C1(n640), .C2(n377), .A(n2162), .ZN(
        n2155) );
  NOR4_X1 U732 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2135) );
  OAI221_X1 U733 ( .B1(n991), .B2(n356), .C1(n959), .C2(n353), .A(n2143), .ZN(
        n2136) );
  OAI221_X1 U734 ( .B1(n863), .B2(n368), .C1(n831), .C2(n365), .A(n2142), .ZN(
        n2137) );
  OAI221_X1 U735 ( .B1(n671), .B2(n380), .C1(n639), .C2(n377), .A(n2141), .ZN(
        n2138) );
  NOR4_X1 U736 ( .A1(n2119), .A2(n2120), .A3(n2121), .A4(n2122), .ZN(n2118) );
  OAI221_X1 U737 ( .B1(n990), .B2(n356), .C1(n958), .C2(n353), .A(n2126), .ZN(
        n2119) );
  OAI221_X1 U738 ( .B1(n862), .B2(n368), .C1(n830), .C2(n365), .A(n2125), .ZN(
        n2120) );
  OAI221_X1 U739 ( .B1(n670), .B2(n380), .C1(n638), .C2(n377), .A(n2124), .ZN(
        n2121) );
  NOR4_X1 U740 ( .A1(n2102), .A2(n2103), .A3(n2104), .A4(n2105), .ZN(n2101) );
  OAI221_X1 U741 ( .B1(n989), .B2(n356), .C1(n957), .C2(n353), .A(n2109), .ZN(
        n2102) );
  OAI221_X1 U742 ( .B1(n861), .B2(n368), .C1(n829), .C2(n365), .A(n2108), .ZN(
        n2103) );
  OAI221_X1 U743 ( .B1(n669), .B2(n380), .C1(n637), .C2(n377), .A(n2107), .ZN(
        n2104) );
  NOR4_X1 U744 ( .A1(n2085), .A2(n2086), .A3(n2087), .A4(n2088), .ZN(n2084) );
  OAI221_X1 U745 ( .B1(n988), .B2(n356), .C1(n956), .C2(n353), .A(n2092), .ZN(
        n2085) );
  OAI221_X1 U746 ( .B1(n860), .B2(n368), .C1(n828), .C2(n365), .A(n2091), .ZN(
        n2086) );
  OAI221_X1 U747 ( .B1(n668), .B2(n380), .C1(n636), .C2(n377), .A(n2090), .ZN(
        n2087) );
  NOR4_X1 U748 ( .A1(n2068), .A2(n2069), .A3(n2070), .A4(n2071), .ZN(n2067) );
  OAI221_X1 U749 ( .B1(n987), .B2(n356), .C1(n955), .C2(n353), .A(n2075), .ZN(
        n2068) );
  OAI221_X1 U750 ( .B1(n859), .B2(n368), .C1(n827), .C2(n365), .A(n2074), .ZN(
        n2069) );
  OAI221_X1 U751 ( .B1(n667), .B2(n380), .C1(n635), .C2(n377), .A(n2073), .ZN(
        n2070) );
  NOR4_X1 U752 ( .A1(n2051), .A2(n2052), .A3(n2053), .A4(n2054), .ZN(n2050) );
  OAI221_X1 U753 ( .B1(n986), .B2(n356), .C1(n954), .C2(n353), .A(n2058), .ZN(
        n2051) );
  OAI221_X1 U754 ( .B1(n858), .B2(n368), .C1(n826), .C2(n365), .A(n2057), .ZN(
        n2052) );
  OAI221_X1 U755 ( .B1(n666), .B2(n380), .C1(n634), .C2(n377), .A(n2056), .ZN(
        n2053) );
  NOR4_X1 U756 ( .A1(n2034), .A2(n2035), .A3(n2036), .A4(n2037), .ZN(n2033) );
  OAI221_X1 U757 ( .B1(n985), .B2(n356), .C1(n953), .C2(n353), .A(n2041), .ZN(
        n2034) );
  OAI221_X1 U758 ( .B1(n857), .B2(n368), .C1(n825), .C2(n365), .A(n2040), .ZN(
        n2035) );
  OAI221_X1 U759 ( .B1(n665), .B2(n380), .C1(n633), .C2(n377), .A(n2039), .ZN(
        n2036) );
  NOR4_X1 U760 ( .A1(n2017), .A2(n2018), .A3(n2019), .A4(n2020), .ZN(n2016) );
  OAI221_X1 U761 ( .B1(n984), .B2(n356), .C1(n952), .C2(n353), .A(n2024), .ZN(
        n2017) );
  OAI221_X1 U762 ( .B1(n856), .B2(n368), .C1(n824), .C2(n365), .A(n2023), .ZN(
        n2018) );
  OAI221_X1 U763 ( .B1(n664), .B2(n380), .C1(n632), .C2(n377), .A(n2022), .ZN(
        n2019) );
  NOR4_X1 U764 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(n1999) );
  OAI221_X1 U765 ( .B1(n983), .B2(n356), .C1(n951), .C2(n353), .A(n2007), .ZN(
        n2000) );
  OAI221_X1 U766 ( .B1(n855), .B2(n368), .C1(n823), .C2(n365), .A(n2006), .ZN(
        n2001) );
  OAI221_X1 U767 ( .B1(n663), .B2(n380), .C1(n631), .C2(n377), .A(n2005), .ZN(
        n2002) );
  NOR4_X1 U768 ( .A1(n1983), .A2(n1984), .A3(n1985), .A4(n1986), .ZN(n1982) );
  OAI221_X1 U769 ( .B1(n982), .B2(n356), .C1(n950), .C2(n353), .A(n1990), .ZN(
        n1983) );
  OAI221_X1 U770 ( .B1(n854), .B2(n368), .C1(n822), .C2(n365), .A(n1989), .ZN(
        n1984) );
  OAI221_X1 U771 ( .B1(n662), .B2(n380), .C1(n630), .C2(n377), .A(n1988), .ZN(
        n1985) );
  NOR4_X1 U772 ( .A1(n1966), .A2(n1967), .A3(n1968), .A4(n1969), .ZN(n1965) );
  OAI221_X1 U773 ( .B1(n981), .B2(n357), .C1(n949), .C2(n354), .A(n1973), .ZN(
        n1966) );
  OAI221_X1 U774 ( .B1(n853), .B2(n369), .C1(n821), .C2(n366), .A(n1972), .ZN(
        n1967) );
  OAI221_X1 U775 ( .B1(n661), .B2(n381), .C1(n629), .C2(n378), .A(n1971), .ZN(
        n1968) );
  NOR4_X1 U776 ( .A1(n1949), .A2(n1950), .A3(n1951), .A4(n1952), .ZN(n1948) );
  OAI221_X1 U777 ( .B1(n980), .B2(n357), .C1(n948), .C2(n354), .A(n1956), .ZN(
        n1949) );
  OAI221_X1 U778 ( .B1(n852), .B2(n369), .C1(n820), .C2(n366), .A(n1955), .ZN(
        n1950) );
  OAI221_X1 U779 ( .B1(n660), .B2(n381), .C1(n628), .C2(n378), .A(n1954), .ZN(
        n1951) );
  NOR4_X1 U780 ( .A1(n1932), .A2(n1933), .A3(n1934), .A4(n1935), .ZN(n1931) );
  OAI221_X1 U781 ( .B1(n979), .B2(n357), .C1(n947), .C2(n354), .A(n1939), .ZN(
        n1932) );
  OAI221_X1 U782 ( .B1(n851), .B2(n369), .C1(n819), .C2(n366), .A(n1938), .ZN(
        n1933) );
  OAI221_X1 U783 ( .B1(n659), .B2(n381), .C1(n627), .C2(n378), .A(n1937), .ZN(
        n1934) );
  NOR4_X1 U784 ( .A1(n1915), .A2(n1916), .A3(n1917), .A4(n1918), .ZN(n1914) );
  OAI221_X1 U785 ( .B1(n978), .B2(n357), .C1(n946), .C2(n354), .A(n1922), .ZN(
        n1915) );
  OAI221_X1 U786 ( .B1(n850), .B2(n369), .C1(n818), .C2(n366), .A(n1921), .ZN(
        n1916) );
  OAI221_X1 U787 ( .B1(n658), .B2(n381), .C1(n626), .C2(n378), .A(n1920), .ZN(
        n1917) );
  NOR4_X1 U788 ( .A1(n1898), .A2(n1899), .A3(n1900), .A4(n1901), .ZN(n1897) );
  OAI221_X1 U789 ( .B1(n977), .B2(n357), .C1(n945), .C2(n354), .A(n1905), .ZN(
        n1898) );
  OAI221_X1 U790 ( .B1(n849), .B2(n369), .C1(n817), .C2(n366), .A(n1904), .ZN(
        n1899) );
  OAI221_X1 U791 ( .B1(n657), .B2(n381), .C1(n625), .C2(n378), .A(n1903), .ZN(
        n1900) );
  NOR4_X1 U792 ( .A1(n1881), .A2(n1882), .A3(n1883), .A4(n1884), .ZN(n1880) );
  OAI221_X1 U793 ( .B1(n976), .B2(n357), .C1(n944), .C2(n354), .A(n1888), .ZN(
        n1881) );
  OAI221_X1 U794 ( .B1(n848), .B2(n369), .C1(n816), .C2(n366), .A(n1887), .ZN(
        n1882) );
  OAI221_X1 U795 ( .B1(n656), .B2(n381), .C1(n624), .C2(n378), .A(n1886), .ZN(
        n1883) );
  NOR4_X1 U796 ( .A1(n1864), .A2(n1865), .A3(n1866), .A4(n1867), .ZN(n1863) );
  OAI221_X1 U797 ( .B1(n975), .B2(n357), .C1(n943), .C2(n354), .A(n1871), .ZN(
        n1864) );
  OAI221_X1 U798 ( .B1(n847), .B2(n369), .C1(n815), .C2(n366), .A(n1870), .ZN(
        n1865) );
  OAI221_X1 U799 ( .B1(n655), .B2(n381), .C1(n623), .C2(n378), .A(n1869), .ZN(
        n1866) );
  NOR4_X1 U800 ( .A1(n1847), .A2(n1848), .A3(n1849), .A4(n1850), .ZN(n1846) );
  OAI221_X1 U801 ( .B1(n974), .B2(n357), .C1(n942), .C2(n354), .A(n1854), .ZN(
        n1847) );
  OAI221_X1 U802 ( .B1(n846), .B2(n369), .C1(n814), .C2(n366), .A(n1853), .ZN(
        n1848) );
  OAI221_X1 U803 ( .B1(n654), .B2(n381), .C1(n622), .C2(n378), .A(n1852), .ZN(
        n1849) );
  NOR4_X1 U804 ( .A1(n1830), .A2(n1831), .A3(n1832), .A4(n1833), .ZN(n1829) );
  OAI221_X1 U805 ( .B1(n973), .B2(n357), .C1(n941), .C2(n354), .A(n1837), .ZN(
        n1830) );
  OAI221_X1 U806 ( .B1(n845), .B2(n369), .C1(n813), .C2(n366), .A(n1836), .ZN(
        n1831) );
  OAI221_X1 U807 ( .B1(n653), .B2(n381), .C1(n621), .C2(n378), .A(n1835), .ZN(
        n1832) );
  NOR4_X1 U808 ( .A1(n1813), .A2(n1814), .A3(n1815), .A4(n1816), .ZN(n1812) );
  OAI221_X1 U809 ( .B1(n972), .B2(n357), .C1(n940), .C2(n354), .A(n1820), .ZN(
        n1813) );
  OAI221_X1 U810 ( .B1(n844), .B2(n369), .C1(n812), .C2(n366), .A(n1819), .ZN(
        n1814) );
  OAI221_X1 U811 ( .B1(n652), .B2(n381), .C1(n620), .C2(n378), .A(n1818), .ZN(
        n1815) );
  NOR4_X1 U812 ( .A1(n1796), .A2(n1797), .A3(n1798), .A4(n1799), .ZN(n1795) );
  OAI221_X1 U813 ( .B1(n971), .B2(n357), .C1(n939), .C2(n354), .A(n1803), .ZN(
        n1796) );
  OAI221_X1 U814 ( .B1(n843), .B2(n369), .C1(n811), .C2(n366), .A(n1802), .ZN(
        n1797) );
  OAI221_X1 U815 ( .B1(n651), .B2(n381), .C1(n619), .C2(n378), .A(n1801), .ZN(
        n1798) );
  NOR4_X1 U816 ( .A1(n2744), .A2(n2745), .A3(n2746), .A4(n2747), .ZN(n2743) );
  OAI221_X1 U817 ( .B1(n992), .B2(n199), .C1(n960), .C2(n196), .A(n2760), .ZN(
        n2744) );
  OAI221_X1 U818 ( .B1(n864), .B2(n211), .C1(n832), .C2(n208), .A(n2757), .ZN(
        n2745) );
  OAI221_X1 U819 ( .B1(n672), .B2(n223), .C1(n640), .C2(n220), .A(n2753), .ZN(
        n2746) );
  NOR4_X1 U820 ( .A1(n2727), .A2(n2728), .A3(n2729), .A4(n2730), .ZN(n2726) );
  OAI221_X1 U821 ( .B1(n991), .B2(n199), .C1(n959), .C2(n196), .A(n2734), .ZN(
        n2727) );
  OAI221_X1 U822 ( .B1(n863), .B2(n211), .C1(n831), .C2(n208), .A(n2733), .ZN(
        n2728) );
  OAI221_X1 U823 ( .B1(n671), .B2(n223), .C1(n639), .C2(n220), .A(n2732), .ZN(
        n2729) );
  NOR4_X1 U824 ( .A1(n2710), .A2(n2711), .A3(n2712), .A4(n2713), .ZN(n2709) );
  OAI221_X1 U825 ( .B1(n990), .B2(n199), .C1(n958), .C2(n196), .A(n2717), .ZN(
        n2710) );
  OAI221_X1 U826 ( .B1(n862), .B2(n211), .C1(n830), .C2(n208), .A(n2716), .ZN(
        n2711) );
  OAI221_X1 U827 ( .B1(n670), .B2(n223), .C1(n638), .C2(n220), .A(n2715), .ZN(
        n2712) );
  NOR4_X1 U828 ( .A1(n2693), .A2(n2694), .A3(n2695), .A4(n2696), .ZN(n2692) );
  OAI221_X1 U829 ( .B1(n989), .B2(n199), .C1(n957), .C2(n196), .A(n2700), .ZN(
        n2693) );
  OAI221_X1 U830 ( .B1(n861), .B2(n211), .C1(n829), .C2(n208), .A(n2699), .ZN(
        n2694) );
  OAI221_X1 U831 ( .B1(n669), .B2(n223), .C1(n637), .C2(n220), .A(n2698), .ZN(
        n2695) );
  NOR4_X1 U832 ( .A1(n2676), .A2(n2677), .A3(n2678), .A4(n2679), .ZN(n2675) );
  OAI221_X1 U833 ( .B1(n988), .B2(n199), .C1(n956), .C2(n196), .A(n2683), .ZN(
        n2676) );
  OAI221_X1 U834 ( .B1(n860), .B2(n211), .C1(n828), .C2(n208), .A(n2682), .ZN(
        n2677) );
  OAI221_X1 U835 ( .B1(n668), .B2(n223), .C1(n636), .C2(n220), .A(n2681), .ZN(
        n2678) );
  NOR4_X1 U836 ( .A1(n2659), .A2(n2660), .A3(n2661), .A4(n2662), .ZN(n2658) );
  OAI221_X1 U837 ( .B1(n987), .B2(n199), .C1(n955), .C2(n196), .A(n2666), .ZN(
        n2659) );
  OAI221_X1 U838 ( .B1(n859), .B2(n211), .C1(n827), .C2(n208), .A(n2665), .ZN(
        n2660) );
  OAI221_X1 U839 ( .B1(n667), .B2(n223), .C1(n635), .C2(n220), .A(n2664), .ZN(
        n2661) );
  NOR4_X1 U840 ( .A1(n2642), .A2(n2643), .A3(n2644), .A4(n2645), .ZN(n2641) );
  OAI221_X1 U841 ( .B1(n986), .B2(n199), .C1(n954), .C2(n196), .A(n2649), .ZN(
        n2642) );
  OAI221_X1 U842 ( .B1(n858), .B2(n211), .C1(n826), .C2(n208), .A(n2648), .ZN(
        n2643) );
  OAI221_X1 U843 ( .B1(n666), .B2(n223), .C1(n634), .C2(n220), .A(n2647), .ZN(
        n2644) );
  NOR4_X1 U844 ( .A1(n2625), .A2(n2626), .A3(n2627), .A4(n2628), .ZN(n2624) );
  OAI221_X1 U845 ( .B1(n985), .B2(n199), .C1(n953), .C2(n196), .A(n2632), .ZN(
        n2625) );
  OAI221_X1 U846 ( .B1(n857), .B2(n211), .C1(n825), .C2(n208), .A(n2631), .ZN(
        n2626) );
  OAI221_X1 U847 ( .B1(n665), .B2(n223), .C1(n633), .C2(n220), .A(n2630), .ZN(
        n2627) );
  NOR4_X1 U848 ( .A1(n2608), .A2(n2609), .A3(n2610), .A4(n2611), .ZN(n2607) );
  OAI221_X1 U849 ( .B1(n984), .B2(n199), .C1(n952), .C2(n196), .A(n2615), .ZN(
        n2608) );
  OAI221_X1 U850 ( .B1(n856), .B2(n211), .C1(n824), .C2(n208), .A(n2614), .ZN(
        n2609) );
  OAI221_X1 U851 ( .B1(n664), .B2(n223), .C1(n632), .C2(n220), .A(n2613), .ZN(
        n2610) );
  NOR4_X1 U852 ( .A1(n2591), .A2(n2592), .A3(n2593), .A4(n2594), .ZN(n2590) );
  OAI221_X1 U853 ( .B1(n983), .B2(n199), .C1(n951), .C2(n196), .A(n2598), .ZN(
        n2591) );
  OAI221_X1 U854 ( .B1(n855), .B2(n211), .C1(n823), .C2(n208), .A(n2597), .ZN(
        n2592) );
  OAI221_X1 U855 ( .B1(n663), .B2(n223), .C1(n631), .C2(n220), .A(n2596), .ZN(
        n2593) );
  NOR4_X1 U856 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2577), .ZN(n2573) );
  OAI221_X1 U857 ( .B1(n982), .B2(n199), .C1(n950), .C2(n196), .A(n2581), .ZN(
        n2574) );
  OAI221_X1 U858 ( .B1(n854), .B2(n211), .C1(n822), .C2(n208), .A(n2580), .ZN(
        n2575) );
  OAI221_X1 U859 ( .B1(n662), .B2(n223), .C1(n630), .C2(n220), .A(n2579), .ZN(
        n2576) );
  NOR4_X1 U860 ( .A1(n2557), .A2(n2558), .A3(n2559), .A4(n2560), .ZN(n2556) );
  OAI221_X1 U861 ( .B1(n981), .B2(n200), .C1(n949), .C2(n197), .A(n2564), .ZN(
        n2557) );
  OAI221_X1 U862 ( .B1(n853), .B2(n212), .C1(n821), .C2(n209), .A(n2563), .ZN(
        n2558) );
  OAI221_X1 U863 ( .B1(n661), .B2(n224), .C1(n629), .C2(n221), .A(n2562), .ZN(
        n2559) );
  NOR4_X1 U864 ( .A1(n2540), .A2(n2541), .A3(n2542), .A4(n2543), .ZN(n2539) );
  OAI221_X1 U865 ( .B1(n980), .B2(n200), .C1(n948), .C2(n197), .A(n2547), .ZN(
        n2540) );
  OAI221_X1 U866 ( .B1(n852), .B2(n212), .C1(n820), .C2(n209), .A(n2546), .ZN(
        n2541) );
  OAI221_X1 U867 ( .B1(n660), .B2(n224), .C1(n628), .C2(n221), .A(n2545), .ZN(
        n2542) );
  NOR4_X1 U868 ( .A1(n2523), .A2(n2524), .A3(n2525), .A4(n2526), .ZN(n2522) );
  OAI221_X1 U869 ( .B1(n979), .B2(n200), .C1(n947), .C2(n197), .A(n2530), .ZN(
        n2523) );
  OAI221_X1 U870 ( .B1(n851), .B2(n212), .C1(n819), .C2(n209), .A(n2529), .ZN(
        n2524) );
  OAI221_X1 U871 ( .B1(n659), .B2(n224), .C1(n627), .C2(n221), .A(n2528), .ZN(
        n2525) );
  NOR4_X1 U872 ( .A1(n2506), .A2(n2507), .A3(n2508), .A4(n2509), .ZN(n2505) );
  OAI221_X1 U873 ( .B1(n978), .B2(n200), .C1(n946), .C2(n197), .A(n2513), .ZN(
        n2506) );
  OAI221_X1 U874 ( .B1(n850), .B2(n212), .C1(n818), .C2(n209), .A(n2512), .ZN(
        n2507) );
  OAI221_X1 U875 ( .B1(n658), .B2(n224), .C1(n626), .C2(n221), .A(n2511), .ZN(
        n2508) );
  NOR4_X1 U876 ( .A1(n2489), .A2(n2490), .A3(n2491), .A4(n2492), .ZN(n2488) );
  OAI221_X1 U877 ( .B1(n977), .B2(n200), .C1(n945), .C2(n197), .A(n2496), .ZN(
        n2489) );
  OAI221_X1 U878 ( .B1(n849), .B2(n212), .C1(n817), .C2(n209), .A(n2495), .ZN(
        n2490) );
  OAI221_X1 U879 ( .B1(n657), .B2(n224), .C1(n625), .C2(n221), .A(n2494), .ZN(
        n2491) );
  NOR4_X1 U880 ( .A1(n2472), .A2(n2473), .A3(n2474), .A4(n2475), .ZN(n2471) );
  OAI221_X1 U881 ( .B1(n976), .B2(n200), .C1(n944), .C2(n197), .A(n2479), .ZN(
        n2472) );
  OAI221_X1 U882 ( .B1(n848), .B2(n212), .C1(n816), .C2(n209), .A(n2478), .ZN(
        n2473) );
  OAI221_X1 U883 ( .B1(n656), .B2(n224), .C1(n624), .C2(n221), .A(n2477), .ZN(
        n2474) );
  NOR4_X1 U884 ( .A1(n2455), .A2(n2456), .A3(n2457), .A4(n2458), .ZN(n2454) );
  OAI221_X1 U885 ( .B1(n975), .B2(n200), .C1(n943), .C2(n197), .A(n2462), .ZN(
        n2455) );
  OAI221_X1 U886 ( .B1(n847), .B2(n212), .C1(n815), .C2(n209), .A(n2461), .ZN(
        n2456) );
  OAI221_X1 U887 ( .B1(n655), .B2(n224), .C1(n623), .C2(n221), .A(n2460), .ZN(
        n2457) );
  NOR4_X1 U888 ( .A1(n2438), .A2(n2439), .A3(n2440), .A4(n2441), .ZN(n2437) );
  OAI221_X1 U889 ( .B1(n974), .B2(n200), .C1(n942), .C2(n197), .A(n2445), .ZN(
        n2438) );
  OAI221_X1 U890 ( .B1(n846), .B2(n212), .C1(n814), .C2(n209), .A(n2444), .ZN(
        n2439) );
  OAI221_X1 U891 ( .B1(n654), .B2(n224), .C1(n622), .C2(n221), .A(n2443), .ZN(
        n2440) );
  NOR4_X1 U892 ( .A1(n2421), .A2(n2422), .A3(n2423), .A4(n2424), .ZN(n2420) );
  OAI221_X1 U893 ( .B1(n973), .B2(n200), .C1(n941), .C2(n197), .A(n2428), .ZN(
        n2421) );
  OAI221_X1 U894 ( .B1(n845), .B2(n212), .C1(n813), .C2(n209), .A(n2427), .ZN(
        n2422) );
  OAI221_X1 U895 ( .B1(n653), .B2(n224), .C1(n621), .C2(n221), .A(n2426), .ZN(
        n2423) );
  NOR4_X1 U896 ( .A1(n2404), .A2(n2405), .A3(n2406), .A4(n2407), .ZN(n2403) );
  OAI221_X1 U897 ( .B1(n972), .B2(n200), .C1(n940), .C2(n197), .A(n2411), .ZN(
        n2404) );
  OAI221_X1 U898 ( .B1(n844), .B2(n212), .C1(n812), .C2(n209), .A(n2410), .ZN(
        n2405) );
  OAI221_X1 U899 ( .B1(n652), .B2(n224), .C1(n620), .C2(n221), .A(n2409), .ZN(
        n2406) );
  NOR4_X1 U900 ( .A1(n2387), .A2(n2388), .A3(n2389), .A4(n2390), .ZN(n2386) );
  OAI221_X1 U901 ( .B1(n971), .B2(n200), .C1(n939), .C2(n197), .A(n2394), .ZN(
        n2387) );
  OAI221_X1 U902 ( .B1(n843), .B2(n212), .C1(n811), .C2(n209), .A(n2393), .ZN(
        n2388) );
  OAI221_X1 U903 ( .B1(n651), .B2(n224), .C1(n619), .C2(n221), .A(n2392), .ZN(
        n2389) );
  OAI221_X1 U904 ( .B1(n544), .B2(n392), .C1(n512), .C2(n389), .A(n2157), .ZN(
        n2156) );
  AOI22_X1 U905 ( .A1(n386), .A2(\registers[19][0] ), .B1(n383), .B2(
        \registers[18][0] ), .ZN(n2157) );
  OAI221_X1 U906 ( .B1(n543), .B2(n392), .C1(n511), .C2(n389), .A(n2140), .ZN(
        n2139) );
  AOI22_X1 U907 ( .A1(n386), .A2(\registers[19][1] ), .B1(n383), .B2(
        \registers[18][1] ), .ZN(n2140) );
  OAI221_X1 U908 ( .B1(n542), .B2(n392), .C1(n510), .C2(n389), .A(n2123), .ZN(
        n2122) );
  AOI22_X1 U909 ( .A1(n386), .A2(\registers[19][2] ), .B1(n383), .B2(
        \registers[18][2] ), .ZN(n2123) );
  OAI221_X1 U910 ( .B1(n541), .B2(n392), .C1(n509), .C2(n389), .A(n2106), .ZN(
        n2105) );
  AOI22_X1 U911 ( .A1(n386), .A2(\registers[19][3] ), .B1(n383), .B2(
        \registers[18][3] ), .ZN(n2106) );
  OAI221_X1 U912 ( .B1(n540), .B2(n392), .C1(n508), .C2(n389), .A(n2089), .ZN(
        n2088) );
  AOI22_X1 U913 ( .A1(n386), .A2(\registers[19][4] ), .B1(n383), .B2(
        \registers[18][4] ), .ZN(n2089) );
  OAI221_X1 U914 ( .B1(n539), .B2(n392), .C1(n507), .C2(n389), .A(n2072), .ZN(
        n2071) );
  AOI22_X1 U915 ( .A1(n386), .A2(\registers[19][5] ), .B1(n383), .B2(
        \registers[18][5] ), .ZN(n2072) );
  OAI221_X1 U916 ( .B1(n538), .B2(n392), .C1(n506), .C2(n389), .A(n2055), .ZN(
        n2054) );
  AOI22_X1 U917 ( .A1(n386), .A2(\registers[19][6] ), .B1(n383), .B2(
        \registers[18][6] ), .ZN(n2055) );
  OAI221_X1 U918 ( .B1(n537), .B2(n392), .C1(n505), .C2(n389), .A(n2038), .ZN(
        n2037) );
  AOI22_X1 U919 ( .A1(n386), .A2(\registers[19][7] ), .B1(n383), .B2(
        \registers[18][7] ), .ZN(n2038) );
  OAI221_X1 U920 ( .B1(n536), .B2(n392), .C1(n504), .C2(n389), .A(n2021), .ZN(
        n2020) );
  AOI22_X1 U921 ( .A1(n386), .A2(\registers[19][8] ), .B1(n383), .B2(
        \registers[18][8] ), .ZN(n2021) );
  OAI221_X1 U922 ( .B1(n535), .B2(n392), .C1(n503), .C2(n389), .A(n2004), .ZN(
        n2003) );
  AOI22_X1 U923 ( .A1(n386), .A2(\registers[19][9] ), .B1(n383), .B2(
        \registers[18][9] ), .ZN(n2004) );
  OAI221_X1 U924 ( .B1(n534), .B2(n392), .C1(n502), .C2(n389), .A(n1987), .ZN(
        n1986) );
  AOI22_X1 U925 ( .A1(n386), .A2(\registers[19][10] ), .B1(n383), .B2(
        \registers[18][10] ), .ZN(n1987) );
  OAI221_X1 U926 ( .B1(n544), .B2(n235), .C1(n512), .C2(n232), .A(n2748), .ZN(
        n2747) );
  AOI22_X1 U927 ( .A1(n229), .A2(\registers[19][0] ), .B1(n226), .B2(
        \registers[18][0] ), .ZN(n2748) );
  OAI221_X1 U928 ( .B1(n543), .B2(n235), .C1(n511), .C2(n232), .A(n2731), .ZN(
        n2730) );
  AOI22_X1 U929 ( .A1(n229), .A2(\registers[19][1] ), .B1(n226), .B2(
        \registers[18][1] ), .ZN(n2731) );
  OAI221_X1 U930 ( .B1(n542), .B2(n235), .C1(n510), .C2(n232), .A(n2714), .ZN(
        n2713) );
  AOI22_X1 U931 ( .A1(n229), .A2(\registers[19][2] ), .B1(n226), .B2(
        \registers[18][2] ), .ZN(n2714) );
  OAI221_X1 U932 ( .B1(n541), .B2(n235), .C1(n509), .C2(n232), .A(n2697), .ZN(
        n2696) );
  AOI22_X1 U933 ( .A1(n229), .A2(\registers[19][3] ), .B1(n226), .B2(
        \registers[18][3] ), .ZN(n2697) );
  OAI221_X1 U934 ( .B1(n540), .B2(n235), .C1(n508), .C2(n232), .A(n2680), .ZN(
        n2679) );
  AOI22_X1 U935 ( .A1(n229), .A2(\registers[19][4] ), .B1(n226), .B2(
        \registers[18][4] ), .ZN(n2680) );
  OAI221_X1 U936 ( .B1(n539), .B2(n235), .C1(n507), .C2(n232), .A(n2663), .ZN(
        n2662) );
  AOI22_X1 U937 ( .A1(n229), .A2(\registers[19][5] ), .B1(n226), .B2(
        \registers[18][5] ), .ZN(n2663) );
  OAI221_X1 U938 ( .B1(n538), .B2(n235), .C1(n506), .C2(n232), .A(n2646), .ZN(
        n2645) );
  AOI22_X1 U939 ( .A1(n229), .A2(\registers[19][6] ), .B1(n226), .B2(
        \registers[18][6] ), .ZN(n2646) );
  OAI221_X1 U940 ( .B1(n537), .B2(n235), .C1(n505), .C2(n232), .A(n2629), .ZN(
        n2628) );
  AOI22_X1 U941 ( .A1(n229), .A2(\registers[19][7] ), .B1(n226), .B2(
        \registers[18][7] ), .ZN(n2629) );
  OAI221_X1 U942 ( .B1(n536), .B2(n235), .C1(n504), .C2(n232), .A(n2612), .ZN(
        n2611) );
  AOI22_X1 U943 ( .A1(n229), .A2(\registers[19][8] ), .B1(n226), .B2(
        \registers[18][8] ), .ZN(n2612) );
  OAI221_X1 U944 ( .B1(n535), .B2(n235), .C1(n503), .C2(n232), .A(n2595), .ZN(
        n2594) );
  AOI22_X1 U945 ( .A1(n229), .A2(\registers[19][9] ), .B1(n226), .B2(
        \registers[18][9] ), .ZN(n2595) );
  OAI221_X1 U946 ( .B1(n534), .B2(n235), .C1(n502), .C2(n232), .A(n2578), .ZN(
        n2577) );
  AOI22_X1 U947 ( .A1(n229), .A2(\registers[19][10] ), .B1(n226), .B2(
        \registers[18][10] ), .ZN(n2578) );
  OAI221_X1 U948 ( .B1(n522), .B2(n394), .C1(n490), .C2(n391), .A(n1783), .ZN(
        n1782) );
  AOI22_X1 U949 ( .A1(n388), .A2(\registers[19][22] ), .B1(n385), .B2(
        \registers[18][22] ), .ZN(n1783) );
  OAI221_X1 U950 ( .B1(n521), .B2(n394), .C1(n489), .C2(n391), .A(n1766), .ZN(
        n1765) );
  AOI22_X1 U951 ( .A1(n388), .A2(\registers[19][23] ), .B1(n385), .B2(
        \registers[18][23] ), .ZN(n1766) );
  OAI221_X1 U952 ( .B1(n520), .B2(n394), .C1(n488), .C2(n391), .A(n1749), .ZN(
        n1748) );
  AOI22_X1 U953 ( .A1(n388), .A2(\registers[19][24] ), .B1(n385), .B2(
        \registers[18][24] ), .ZN(n1749) );
  OAI221_X1 U954 ( .B1(n519), .B2(n394), .C1(n487), .C2(n391), .A(n1732), .ZN(
        n1731) );
  AOI22_X1 U955 ( .A1(n388), .A2(\registers[19][25] ), .B1(n385), .B2(
        \registers[18][25] ), .ZN(n1732) );
  OAI221_X1 U956 ( .B1(n518), .B2(n394), .C1(n486), .C2(n391), .A(n1715), .ZN(
        n1714) );
  AOI22_X1 U957 ( .A1(n388), .A2(\registers[19][26] ), .B1(n385), .B2(
        \registers[18][26] ), .ZN(n1715) );
  OAI221_X1 U958 ( .B1(n517), .B2(n394), .C1(n485), .C2(n391), .A(n1698), .ZN(
        n1697) );
  AOI22_X1 U959 ( .A1(n388), .A2(\registers[19][27] ), .B1(n385), .B2(
        \registers[18][27] ), .ZN(n1698) );
  OAI221_X1 U960 ( .B1(n516), .B2(n394), .C1(n484), .C2(n391), .A(n1681), .ZN(
        n1680) );
  AOI22_X1 U961 ( .A1(n388), .A2(\registers[19][28] ), .B1(n385), .B2(
        \registers[18][28] ), .ZN(n1681) );
  OAI221_X1 U962 ( .B1(n515), .B2(n394), .C1(n483), .C2(n391), .A(n1664), .ZN(
        n1663) );
  AOI22_X1 U963 ( .A1(n388), .A2(\registers[19][29] ), .B1(n385), .B2(
        \registers[18][29] ), .ZN(n1664) );
  OAI221_X1 U964 ( .B1(n514), .B2(n394), .C1(n482), .C2(n391), .A(n1647), .ZN(
        n1646) );
  AOI22_X1 U965 ( .A1(n388), .A2(\registers[19][30] ), .B1(n385), .B2(
        \registers[18][30] ), .ZN(n1647) );
  OAI221_X1 U966 ( .B1(n513), .B2(n394), .C1(n481), .C2(n391), .A(n1601), .ZN(
        n1598) );
  AOI22_X1 U967 ( .A1(n388), .A2(\registers[19][31] ), .B1(n385), .B2(
        \registers[18][31] ), .ZN(n1601) );
  OAI221_X1 U968 ( .B1(n522), .B2(n237), .C1(n490), .C2(n234), .A(n2374), .ZN(
        n2373) );
  AOI22_X1 U969 ( .A1(n231), .A2(\registers[19][22] ), .B1(n228), .B2(
        \registers[18][22] ), .ZN(n2374) );
  OAI221_X1 U970 ( .B1(n521), .B2(n237), .C1(n489), .C2(n234), .A(n2357), .ZN(
        n2356) );
  AOI22_X1 U971 ( .A1(n231), .A2(\registers[19][23] ), .B1(n228), .B2(
        \registers[18][23] ), .ZN(n2357) );
  OAI221_X1 U972 ( .B1(n520), .B2(n237), .C1(n488), .C2(n234), .A(n2340), .ZN(
        n2339) );
  AOI22_X1 U973 ( .A1(n231), .A2(\registers[19][24] ), .B1(n228), .B2(
        \registers[18][24] ), .ZN(n2340) );
  OAI221_X1 U974 ( .B1(n519), .B2(n237), .C1(n487), .C2(n234), .A(n2323), .ZN(
        n2322) );
  AOI22_X1 U975 ( .A1(n231), .A2(\registers[19][25] ), .B1(n228), .B2(
        \registers[18][25] ), .ZN(n2323) );
  OAI221_X1 U976 ( .B1(n518), .B2(n237), .C1(n486), .C2(n234), .A(n2306), .ZN(
        n2305) );
  AOI22_X1 U977 ( .A1(n231), .A2(\registers[19][26] ), .B1(n228), .B2(
        \registers[18][26] ), .ZN(n2306) );
  OAI221_X1 U978 ( .B1(n517), .B2(n237), .C1(n485), .C2(n234), .A(n2289), .ZN(
        n2288) );
  AOI22_X1 U979 ( .A1(n231), .A2(\registers[19][27] ), .B1(n228), .B2(
        \registers[18][27] ), .ZN(n2289) );
  OAI221_X1 U980 ( .B1(n516), .B2(n237), .C1(n484), .C2(n234), .A(n2272), .ZN(
        n2271) );
  AOI22_X1 U981 ( .A1(n231), .A2(\registers[19][28] ), .B1(n228), .B2(
        \registers[18][28] ), .ZN(n2272) );
  OAI221_X1 U982 ( .B1(n515), .B2(n237), .C1(n483), .C2(n234), .A(n2255), .ZN(
        n2254) );
  AOI22_X1 U983 ( .A1(n231), .A2(\registers[19][29] ), .B1(n228), .B2(
        \registers[18][29] ), .ZN(n2255) );
  OAI221_X1 U984 ( .B1(n514), .B2(n237), .C1(n482), .C2(n234), .A(n2238), .ZN(
        n2237) );
  AOI22_X1 U985 ( .A1(n231), .A2(\registers[19][30] ), .B1(n228), .B2(
        \registers[18][30] ), .ZN(n2238) );
  OAI221_X1 U986 ( .B1(n513), .B2(n237), .C1(n481), .C2(n234), .A(n2192), .ZN(
        n2189) );
  AOI22_X1 U987 ( .A1(n231), .A2(\registers[19][31] ), .B1(n228), .B2(
        \registers[18][31] ), .ZN(n2192) );
  OAI221_X1 U988 ( .B1(n533), .B2(n393), .C1(n501), .C2(n390), .A(n1970), .ZN(
        n1969) );
  AOI22_X1 U989 ( .A1(n387), .A2(\registers[19][11] ), .B1(n384), .B2(
        \registers[18][11] ), .ZN(n1970) );
  OAI221_X1 U990 ( .B1(n532), .B2(n393), .C1(n500), .C2(n390), .A(n1953), .ZN(
        n1952) );
  AOI22_X1 U991 ( .A1(n387), .A2(\registers[19][12] ), .B1(n384), .B2(
        \registers[18][12] ), .ZN(n1953) );
  OAI221_X1 U992 ( .B1(n531), .B2(n393), .C1(n499), .C2(n390), .A(n1936), .ZN(
        n1935) );
  AOI22_X1 U993 ( .A1(n387), .A2(\registers[19][13] ), .B1(n384), .B2(
        \registers[18][13] ), .ZN(n1936) );
  OAI221_X1 U994 ( .B1(n530), .B2(n393), .C1(n498), .C2(n390), .A(n1919), .ZN(
        n1918) );
  AOI22_X1 U995 ( .A1(n387), .A2(\registers[19][14] ), .B1(n384), .B2(
        \registers[18][14] ), .ZN(n1919) );
  OAI221_X1 U996 ( .B1(n529), .B2(n393), .C1(n497), .C2(n390), .A(n1902), .ZN(
        n1901) );
  AOI22_X1 U997 ( .A1(n387), .A2(\registers[19][15] ), .B1(n384), .B2(
        \registers[18][15] ), .ZN(n1902) );
  OAI221_X1 U998 ( .B1(n528), .B2(n393), .C1(n496), .C2(n390), .A(n1885), .ZN(
        n1884) );
  AOI22_X1 U999 ( .A1(n387), .A2(\registers[19][16] ), .B1(n384), .B2(
        \registers[18][16] ), .ZN(n1885) );
  OAI221_X1 U1000 ( .B1(n527), .B2(n393), .C1(n495), .C2(n390), .A(n1868), 
        .ZN(n1867) );
  AOI22_X1 U1001 ( .A1(n387), .A2(\registers[19][17] ), .B1(n384), .B2(
        \registers[18][17] ), .ZN(n1868) );
  OAI221_X1 U1002 ( .B1(n526), .B2(n393), .C1(n494), .C2(n390), .A(n1851), 
        .ZN(n1850) );
  AOI22_X1 U1003 ( .A1(n387), .A2(\registers[19][18] ), .B1(n384), .B2(
        \registers[18][18] ), .ZN(n1851) );
  OAI221_X1 U1004 ( .B1(n525), .B2(n393), .C1(n493), .C2(n390), .A(n1834), 
        .ZN(n1833) );
  AOI22_X1 U1005 ( .A1(n387), .A2(\registers[19][19] ), .B1(n384), .B2(
        \registers[18][19] ), .ZN(n1834) );
  OAI221_X1 U1006 ( .B1(n524), .B2(n393), .C1(n492), .C2(n390), .A(n1817), 
        .ZN(n1816) );
  AOI22_X1 U1007 ( .A1(n387), .A2(\registers[19][20] ), .B1(n384), .B2(
        \registers[18][20] ), .ZN(n1817) );
  OAI221_X1 U1008 ( .B1(n523), .B2(n393), .C1(n491), .C2(n390), .A(n1800), 
        .ZN(n1799) );
  AOI22_X1 U1009 ( .A1(n387), .A2(\registers[19][21] ), .B1(n384), .B2(
        \registers[18][21] ), .ZN(n1800) );
  OAI221_X1 U1010 ( .B1(n533), .B2(n236), .C1(n501), .C2(n233), .A(n2561), 
        .ZN(n2560) );
  AOI22_X1 U1011 ( .A1(n230), .A2(\registers[19][11] ), .B1(n227), .B2(
        \registers[18][11] ), .ZN(n2561) );
  OAI221_X1 U1012 ( .B1(n532), .B2(n236), .C1(n500), .C2(n233), .A(n2544), 
        .ZN(n2543) );
  AOI22_X1 U1013 ( .A1(n230), .A2(\registers[19][12] ), .B1(n227), .B2(
        \registers[18][12] ), .ZN(n2544) );
  OAI221_X1 U1014 ( .B1(n531), .B2(n236), .C1(n499), .C2(n233), .A(n2527), 
        .ZN(n2526) );
  AOI22_X1 U1015 ( .A1(n230), .A2(\registers[19][13] ), .B1(n227), .B2(
        \registers[18][13] ), .ZN(n2527) );
  OAI221_X1 U1016 ( .B1(n530), .B2(n236), .C1(n498), .C2(n233), .A(n2510), 
        .ZN(n2509) );
  AOI22_X1 U1017 ( .A1(n230), .A2(\registers[19][14] ), .B1(n227), .B2(
        \registers[18][14] ), .ZN(n2510) );
  OAI221_X1 U1018 ( .B1(n529), .B2(n236), .C1(n497), .C2(n233), .A(n2493), 
        .ZN(n2492) );
  AOI22_X1 U1019 ( .A1(n230), .A2(\registers[19][15] ), .B1(n227), .B2(
        \registers[18][15] ), .ZN(n2493) );
  OAI221_X1 U1020 ( .B1(n528), .B2(n236), .C1(n496), .C2(n233), .A(n2476), 
        .ZN(n2475) );
  AOI22_X1 U1021 ( .A1(n230), .A2(\registers[19][16] ), .B1(n227), .B2(
        \registers[18][16] ), .ZN(n2476) );
  OAI221_X1 U1022 ( .B1(n527), .B2(n236), .C1(n495), .C2(n233), .A(n2459), 
        .ZN(n2458) );
  AOI22_X1 U1023 ( .A1(n230), .A2(\registers[19][17] ), .B1(n227), .B2(
        \registers[18][17] ), .ZN(n2459) );
  OAI221_X1 U1024 ( .B1(n526), .B2(n236), .C1(n494), .C2(n233), .A(n2442), 
        .ZN(n2441) );
  AOI22_X1 U1025 ( .A1(n230), .A2(\registers[19][18] ), .B1(n227), .B2(
        \registers[18][18] ), .ZN(n2442) );
  OAI221_X1 U1026 ( .B1(n525), .B2(n236), .C1(n493), .C2(n233), .A(n2425), 
        .ZN(n2424) );
  AOI22_X1 U1027 ( .A1(n230), .A2(\registers[19][19] ), .B1(n227), .B2(
        \registers[18][19] ), .ZN(n2425) );
  OAI221_X1 U1028 ( .B1(n524), .B2(n236), .C1(n492), .C2(n233), .A(n2408), 
        .ZN(n2407) );
  AOI22_X1 U1029 ( .A1(n230), .A2(\registers[19][20] ), .B1(n227), .B2(
        \registers[18][20] ), .ZN(n2408) );
  OAI221_X1 U1030 ( .B1(n523), .B2(n236), .C1(n491), .C2(n233), .A(n2391), 
        .ZN(n2390) );
  AOI22_X1 U1031 ( .A1(n230), .A2(\registers[19][21] ), .B1(n227), .B2(
        \registers[18][21] ), .ZN(n2391) );
  OAI221_X1 U1032 ( .B1(n160), .B2(n271), .C1(n128), .C2(n268), .A(n2175), 
        .ZN(n2171) );
  AOI22_X1 U1033 ( .A1(n265), .A2(\registers[7][0] ), .B1(n262), .B2(
        \registers[6][0] ), .ZN(n2175) );
  OAI221_X1 U1034 ( .B1(n159), .B2(n271), .C1(n127), .C2(n268), .A(n2146), 
        .ZN(n2144) );
  AOI22_X1 U1035 ( .A1(n265), .A2(\registers[7][1] ), .B1(n262), .B2(
        \registers[6][1] ), .ZN(n2146) );
  OAI221_X1 U1036 ( .B1(n158), .B2(n271), .C1(n126), .C2(n268), .A(n2129), 
        .ZN(n2127) );
  AOI22_X1 U1037 ( .A1(n265), .A2(\registers[7][2] ), .B1(n262), .B2(
        \registers[6][2] ), .ZN(n2129) );
  OAI221_X1 U1038 ( .B1(n157), .B2(n271), .C1(n125), .C2(n268), .A(n2112), 
        .ZN(n2110) );
  AOI22_X1 U1039 ( .A1(n265), .A2(\registers[7][3] ), .B1(n262), .B2(
        \registers[6][3] ), .ZN(n2112) );
  OAI221_X1 U1040 ( .B1(n156), .B2(n271), .C1(n124), .C2(n268), .A(n2095), 
        .ZN(n2093) );
  AOI22_X1 U1041 ( .A1(n265), .A2(\registers[7][4] ), .B1(n262), .B2(
        \registers[6][4] ), .ZN(n2095) );
  OAI221_X1 U1042 ( .B1(n155), .B2(n271), .C1(n123), .C2(n268), .A(n2078), 
        .ZN(n2076) );
  AOI22_X1 U1043 ( .A1(n265), .A2(\registers[7][5] ), .B1(n262), .B2(
        \registers[6][5] ), .ZN(n2078) );
  OAI221_X1 U1044 ( .B1(n154), .B2(n271), .C1(n122), .C2(n268), .A(n2061), 
        .ZN(n2059) );
  AOI22_X1 U1045 ( .A1(n265), .A2(\registers[7][6] ), .B1(n262), .B2(
        \registers[6][6] ), .ZN(n2061) );
  OAI221_X1 U1046 ( .B1(n153), .B2(n271), .C1(n121), .C2(n268), .A(n2044), 
        .ZN(n2042) );
  AOI22_X1 U1047 ( .A1(n265), .A2(\registers[7][7] ), .B1(n262), .B2(
        \registers[6][7] ), .ZN(n2044) );
  OAI221_X1 U1048 ( .B1(n152), .B2(n271), .C1(n120), .C2(n268), .A(n2027), 
        .ZN(n2025) );
  AOI22_X1 U1049 ( .A1(n265), .A2(\registers[7][8] ), .B1(n262), .B2(
        \registers[6][8] ), .ZN(n2027) );
  OAI221_X1 U1050 ( .B1(n151), .B2(n271), .C1(n119), .C2(n268), .A(n2010), 
        .ZN(n2008) );
  AOI22_X1 U1051 ( .A1(n265), .A2(\registers[7][9] ), .B1(n262), .B2(
        \registers[6][9] ), .ZN(n2010) );
  OAI221_X1 U1052 ( .B1(n150), .B2(n271), .C1(n118), .C2(n268), .A(n1993), 
        .ZN(n1991) );
  AOI22_X1 U1053 ( .A1(n265), .A2(\registers[7][10] ), .B1(n262), .B2(
        \registers[6][10] ), .ZN(n1993) );
  OAI221_X1 U1054 ( .B1(n138), .B2(n273), .C1(n106), .C2(n270), .A(n1789), 
        .ZN(n1787) );
  AOI22_X1 U1055 ( .A1(n267), .A2(\registers[7][22] ), .B1(n264), .B2(
        \registers[6][22] ), .ZN(n1789) );
  OAI221_X1 U1056 ( .B1(n137), .B2(n273), .C1(n105), .C2(n270), .A(n1772), 
        .ZN(n1770) );
  AOI22_X1 U1057 ( .A1(n267), .A2(\registers[7][23] ), .B1(n264), .B2(
        \registers[6][23] ), .ZN(n1772) );
  OAI221_X1 U1058 ( .B1(n136), .B2(n273), .C1(n104), .C2(n270), .A(n1755), 
        .ZN(n1753) );
  AOI22_X1 U1059 ( .A1(n267), .A2(\registers[7][24] ), .B1(n264), .B2(
        \registers[6][24] ), .ZN(n1755) );
  OAI221_X1 U1060 ( .B1(n135), .B2(n273), .C1(n103), .C2(n270), .A(n1738), 
        .ZN(n1736) );
  AOI22_X1 U1061 ( .A1(n267), .A2(\registers[7][25] ), .B1(n264), .B2(
        \registers[6][25] ), .ZN(n1738) );
  OAI221_X1 U1062 ( .B1(n134), .B2(n273), .C1(n102), .C2(n270), .A(n1721), 
        .ZN(n1719) );
  AOI22_X1 U1063 ( .A1(n267), .A2(\registers[7][26] ), .B1(n264), .B2(
        \registers[6][26] ), .ZN(n1721) );
  OAI221_X1 U1064 ( .B1(n133), .B2(n273), .C1(n101), .C2(n270), .A(n1704), 
        .ZN(n1702) );
  AOI22_X1 U1065 ( .A1(n267), .A2(\registers[7][27] ), .B1(n264), .B2(
        \registers[6][27] ), .ZN(n1704) );
  OAI221_X1 U1066 ( .B1(n132), .B2(n273), .C1(n100), .C2(n270), .A(n1687), 
        .ZN(n1685) );
  AOI22_X1 U1067 ( .A1(n267), .A2(\registers[7][28] ), .B1(n264), .B2(
        \registers[6][28] ), .ZN(n1687) );
  OAI221_X1 U1068 ( .B1(n131), .B2(n273), .C1(n99), .C2(n270), .A(n1670), .ZN(
        n1668) );
  AOI22_X1 U1069 ( .A1(n267), .A2(\registers[7][29] ), .B1(n264), .B2(
        \registers[6][29] ), .ZN(n1670) );
  OAI221_X1 U1070 ( .B1(n130), .B2(n273), .C1(n98), .C2(n270), .A(n1653), .ZN(
        n1651) );
  AOI22_X1 U1071 ( .A1(n267), .A2(\registers[7][30] ), .B1(n264), .B2(
        \registers[6][30] ), .ZN(n1653) );
  OAI221_X1 U1072 ( .B1(n129), .B2(n273), .C1(n97), .C2(n270), .A(n1626), .ZN(
        n1620) );
  AOI22_X1 U1073 ( .A1(n267), .A2(\registers[7][31] ), .B1(n264), .B2(
        \registers[6][31] ), .ZN(n1626) );
  OAI221_X1 U1074 ( .B1(n138), .B2(n180), .C1(n106), .C2(n177), .A(n2380), 
        .ZN(n2378) );
  AOI22_X1 U1075 ( .A1(n174), .A2(\registers[7][22] ), .B1(n171), .B2(
        \registers[6][22] ), .ZN(n2380) );
  OAI221_X1 U1076 ( .B1(n137), .B2(n180), .C1(n105), .C2(n177), .A(n2363), 
        .ZN(n2361) );
  AOI22_X1 U1077 ( .A1(n174), .A2(\registers[7][23] ), .B1(n171), .B2(
        \registers[6][23] ), .ZN(n2363) );
  OAI221_X1 U1078 ( .B1(n136), .B2(n180), .C1(n104), .C2(n177), .A(n2346), 
        .ZN(n2344) );
  AOI22_X1 U1079 ( .A1(n174), .A2(\registers[7][24] ), .B1(n171), .B2(
        \registers[6][24] ), .ZN(n2346) );
  OAI221_X1 U1080 ( .B1(n135), .B2(n180), .C1(n103), .C2(n177), .A(n2329), 
        .ZN(n2327) );
  AOI22_X1 U1081 ( .A1(n174), .A2(\registers[7][25] ), .B1(n171), .B2(
        \registers[6][25] ), .ZN(n2329) );
  OAI221_X1 U1082 ( .B1(n134), .B2(n180), .C1(n102), .C2(n177), .A(n2312), 
        .ZN(n2310) );
  AOI22_X1 U1083 ( .A1(n174), .A2(\registers[7][26] ), .B1(n171), .B2(
        \registers[6][26] ), .ZN(n2312) );
  OAI221_X1 U1084 ( .B1(n133), .B2(n180), .C1(n101), .C2(n177), .A(n2295), 
        .ZN(n2293) );
  AOI22_X1 U1085 ( .A1(n174), .A2(\registers[7][27] ), .B1(n171), .B2(
        \registers[6][27] ), .ZN(n2295) );
  OAI221_X1 U1086 ( .B1(n132), .B2(n180), .C1(n100), .C2(n177), .A(n2278), 
        .ZN(n2276) );
  AOI22_X1 U1087 ( .A1(n174), .A2(\registers[7][28] ), .B1(n171), .B2(
        \registers[6][28] ), .ZN(n2278) );
  OAI221_X1 U1088 ( .B1(n131), .B2(n180), .C1(n99), .C2(n177), .A(n2261), .ZN(
        n2259) );
  AOI22_X1 U1089 ( .A1(n174), .A2(\registers[7][29] ), .B1(n171), .B2(
        \registers[6][29] ), .ZN(n2261) );
  OAI221_X1 U1090 ( .B1(n130), .B2(n180), .C1(n98), .C2(n177), .A(n2244), .ZN(
        n2242) );
  AOI22_X1 U1091 ( .A1(n174), .A2(\registers[7][30] ), .B1(n171), .B2(
        \registers[6][30] ), .ZN(n2244) );
  OAI221_X1 U1092 ( .B1(n129), .B2(n180), .C1(n97), .C2(n177), .A(n2217), .ZN(
        n2211) );
  AOI22_X1 U1093 ( .A1(n174), .A2(\registers[7][31] ), .B1(n171), .B2(
        \registers[6][31] ), .ZN(n2217) );
  OAI221_X1 U1094 ( .B1(n149), .B2(n272), .C1(n117), .C2(n269), .A(n1976), 
        .ZN(n1974) );
  AOI22_X1 U1095 ( .A1(n266), .A2(\registers[7][11] ), .B1(n263), .B2(
        \registers[6][11] ), .ZN(n1976) );
  OAI221_X1 U1096 ( .B1(n148), .B2(n272), .C1(n116), .C2(n269), .A(n1959), 
        .ZN(n1957) );
  AOI22_X1 U1097 ( .A1(n266), .A2(\registers[7][12] ), .B1(n263), .B2(
        \registers[6][12] ), .ZN(n1959) );
  OAI221_X1 U1098 ( .B1(n147), .B2(n272), .C1(n115), .C2(n269), .A(n1942), 
        .ZN(n1940) );
  AOI22_X1 U1099 ( .A1(n266), .A2(\registers[7][13] ), .B1(n263), .B2(
        \registers[6][13] ), .ZN(n1942) );
  OAI221_X1 U1100 ( .B1(n146), .B2(n272), .C1(n114), .C2(n269), .A(n1925), 
        .ZN(n1923) );
  AOI22_X1 U1101 ( .A1(n266), .A2(\registers[7][14] ), .B1(n263), .B2(
        \registers[6][14] ), .ZN(n1925) );
  OAI221_X1 U1102 ( .B1(n145), .B2(n272), .C1(n113), .C2(n269), .A(n1908), 
        .ZN(n1906) );
  AOI22_X1 U1103 ( .A1(n266), .A2(\registers[7][15] ), .B1(n263), .B2(
        \registers[6][15] ), .ZN(n1908) );
  OAI221_X1 U1104 ( .B1(n144), .B2(n272), .C1(n112), .C2(n269), .A(n1891), 
        .ZN(n1889) );
  AOI22_X1 U1105 ( .A1(n266), .A2(\registers[7][16] ), .B1(n263), .B2(
        \registers[6][16] ), .ZN(n1891) );
  OAI221_X1 U1106 ( .B1(n143), .B2(n272), .C1(n111), .C2(n269), .A(n1874), 
        .ZN(n1872) );
  AOI22_X1 U1107 ( .A1(n266), .A2(\registers[7][17] ), .B1(n263), .B2(
        \registers[6][17] ), .ZN(n1874) );
  OAI221_X1 U1108 ( .B1(n142), .B2(n272), .C1(n110), .C2(n269), .A(n1857), 
        .ZN(n1855) );
  AOI22_X1 U1109 ( .A1(n266), .A2(\registers[7][18] ), .B1(n263), .B2(
        \registers[6][18] ), .ZN(n1857) );
  OAI221_X1 U1110 ( .B1(n141), .B2(n272), .C1(n109), .C2(n269), .A(n1840), 
        .ZN(n1838) );
  AOI22_X1 U1111 ( .A1(n266), .A2(\registers[7][19] ), .B1(n263), .B2(
        \registers[6][19] ), .ZN(n1840) );
  OAI221_X1 U1112 ( .B1(n140), .B2(n272), .C1(n108), .C2(n269), .A(n1823), 
        .ZN(n1821) );
  AOI22_X1 U1113 ( .A1(n266), .A2(\registers[7][20] ), .B1(n263), .B2(
        \registers[6][20] ), .ZN(n1823) );
  OAI221_X1 U1114 ( .B1(n139), .B2(n272), .C1(n107), .C2(n269), .A(n1806), 
        .ZN(n1804) );
  AOI22_X1 U1115 ( .A1(n266), .A2(\registers[7][21] ), .B1(n263), .B2(
        \registers[6][21] ), .ZN(n1806) );
  AND2_X1 U1116 ( .A1(ADD_RD2[2]), .A2(n3811), .ZN(n2164) );
  AND2_X1 U1117 ( .A1(ADD_RD1[2]), .A2(n3808), .ZN(n2755) );
  AND2_X1 U1118 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n2163) );
  AND2_X1 U1119 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n2754) );
  OAI22_X1 U1120 ( .A1(n296), .A2(n243), .B1(n328), .B2(n240), .ZN(n1757) );
  OAI22_X1 U1121 ( .A1(n295), .A2(n243), .B1(n327), .B2(n240), .ZN(n1740) );
  OAI22_X1 U1122 ( .A1(n294), .A2(n243), .B1(n326), .B2(n240), .ZN(n1723) );
  OAI22_X1 U1123 ( .A1(n293), .A2(n243), .B1(n325), .B2(n240), .ZN(n1706) );
  OAI22_X1 U1124 ( .A1(n292), .A2(n243), .B1(n324), .B2(n240), .ZN(n1689) );
  OAI22_X1 U1125 ( .A1(n291), .A2(n243), .B1(n323), .B2(n240), .ZN(n1672) );
  OAI22_X1 U1126 ( .A1(n290), .A2(n243), .B1(n322), .B2(n240), .ZN(n1655) );
  OAI22_X1 U1127 ( .A1(n289), .A2(n243), .B1(n321), .B2(n240), .ZN(n1636) );
  OAI22_X1 U1128 ( .A1(n296), .A2(n22), .B1(n328), .B2(n19), .ZN(n2348) );
  OAI22_X1 U1129 ( .A1(n295), .A2(n22), .B1(n327), .B2(n19), .ZN(n2331) );
  OAI22_X1 U1130 ( .A1(n294), .A2(n22), .B1(n326), .B2(n19), .ZN(n2314) );
  OAI22_X1 U1131 ( .A1(n293), .A2(n22), .B1(n325), .B2(n19), .ZN(n2297) );
  OAI22_X1 U1132 ( .A1(n292), .A2(n22), .B1(n324), .B2(n19), .ZN(n2280) );
  OAI22_X1 U1133 ( .A1(n291), .A2(n22), .B1(n323), .B2(n19), .ZN(n2263) );
  OAI22_X1 U1134 ( .A1(n290), .A2(n22), .B1(n322), .B2(n19), .ZN(n2246) );
  OAI22_X1 U1135 ( .A1(n289), .A2(n22), .B1(n321), .B2(n19), .ZN(n2227) );
  OAI22_X1 U1136 ( .A1(n424), .A2(n255), .B1(n456), .B2(n252), .ZN(n1756) );
  OAI22_X1 U1137 ( .A1(n423), .A2(n255), .B1(n455), .B2(n252), .ZN(n1739) );
  OAI22_X1 U1138 ( .A1(n422), .A2(n255), .B1(n454), .B2(n252), .ZN(n1722) );
  OAI22_X1 U1139 ( .A1(n421), .A2(n255), .B1(n453), .B2(n252), .ZN(n1705) );
  OAI22_X1 U1140 ( .A1(n420), .A2(n255), .B1(n452), .B2(n252), .ZN(n1688) );
  OAI22_X1 U1141 ( .A1(n419), .A2(n255), .B1(n451), .B2(n252), .ZN(n1671) );
  OAI22_X1 U1142 ( .A1(n418), .A2(n255), .B1(n450), .B2(n252), .ZN(n1654) );
  OAI22_X1 U1143 ( .A1(n417), .A2(n255), .B1(n449), .B2(n252), .ZN(n1631) );
  OAI22_X1 U1144 ( .A1(n424), .A2(n162), .B1(n456), .B2(n31), .ZN(n2347) );
  OAI22_X1 U1145 ( .A1(n423), .A2(n162), .B1(n455), .B2(n31), .ZN(n2330) );
  OAI22_X1 U1146 ( .A1(n422), .A2(n162), .B1(n454), .B2(n31), .ZN(n2313) );
  OAI22_X1 U1147 ( .A1(n421), .A2(n162), .B1(n453), .B2(n31), .ZN(n2296) );
  OAI22_X1 U1148 ( .A1(n420), .A2(n162), .B1(n452), .B2(n31), .ZN(n2279) );
  OAI22_X1 U1149 ( .A1(n419), .A2(n162), .B1(n451), .B2(n31), .ZN(n2262) );
  OAI22_X1 U1150 ( .A1(n418), .A2(n162), .B1(n450), .B2(n31), .ZN(n2245) );
  OAI22_X1 U1151 ( .A1(n417), .A2(n162), .B1(n449), .B2(n31), .ZN(n2222) );
  OAI22_X1 U1152 ( .A1(n448), .A2(n253), .B1(n480), .B2(n250), .ZN(n2177) );
  OAI22_X1 U1153 ( .A1(n320), .A2(n241), .B1(n352), .B2(n238), .ZN(n2180) );
  OAI22_X1 U1154 ( .A1(n447), .A2(n253), .B1(n479), .B2(n250), .ZN(n2147) );
  OAI22_X1 U1155 ( .A1(n319), .A2(n241), .B1(n351), .B2(n238), .ZN(n2148) );
  OAI22_X1 U1156 ( .A1(n446), .A2(n253), .B1(n478), .B2(n250), .ZN(n2130) );
  OAI22_X1 U1157 ( .A1(n318), .A2(n241), .B1(n350), .B2(n238), .ZN(n2131) );
  OAI22_X1 U1158 ( .A1(n445), .A2(n253), .B1(n477), .B2(n250), .ZN(n2113) );
  OAI22_X1 U1159 ( .A1(n317), .A2(n241), .B1(n349), .B2(n238), .ZN(n2114) );
  OAI22_X1 U1160 ( .A1(n444), .A2(n253), .B1(n476), .B2(n250), .ZN(n2096) );
  OAI22_X1 U1161 ( .A1(n316), .A2(n241), .B1(n348), .B2(n238), .ZN(n2097) );
  OAI22_X1 U1162 ( .A1(n443), .A2(n253), .B1(n475), .B2(n250), .ZN(n2079) );
  OAI22_X1 U1163 ( .A1(n315), .A2(n241), .B1(n347), .B2(n238), .ZN(n2080) );
  OAI22_X1 U1164 ( .A1(n442), .A2(n253), .B1(n474), .B2(n250), .ZN(n2062) );
  OAI22_X1 U1165 ( .A1(n314), .A2(n241), .B1(n346), .B2(n238), .ZN(n2063) );
  OAI22_X1 U1166 ( .A1(n441), .A2(n253), .B1(n473), .B2(n250), .ZN(n2045) );
  OAI22_X1 U1167 ( .A1(n313), .A2(n241), .B1(n345), .B2(n238), .ZN(n2046) );
  OAI22_X1 U1168 ( .A1(n440), .A2(n253), .B1(n472), .B2(n250), .ZN(n2028) );
  OAI22_X1 U1169 ( .A1(n312), .A2(n241), .B1(n344), .B2(n238), .ZN(n2029) );
  OAI22_X1 U1170 ( .A1(n439), .A2(n253), .B1(n471), .B2(n250), .ZN(n2011) );
  OAI22_X1 U1171 ( .A1(n311), .A2(n241), .B1(n343), .B2(n238), .ZN(n2012) );
  OAI22_X1 U1172 ( .A1(n438), .A2(n253), .B1(n470), .B2(n250), .ZN(n1994) );
  OAI22_X1 U1173 ( .A1(n310), .A2(n241), .B1(n342), .B2(n238), .ZN(n1995) );
  OAI22_X1 U1174 ( .A1(n437), .A2(n253), .B1(n469), .B2(n250), .ZN(n1977) );
  OAI22_X1 U1175 ( .A1(n309), .A2(n241), .B1(n341), .B2(n238), .ZN(n1978) );
  OAI22_X1 U1176 ( .A1(n436), .A2(n254), .B1(n468), .B2(n251), .ZN(n1960) );
  OAI22_X1 U1177 ( .A1(n308), .A2(n242), .B1(n340), .B2(n239), .ZN(n1961) );
  OAI22_X1 U1178 ( .A1(n435), .A2(n254), .B1(n467), .B2(n251), .ZN(n1943) );
  OAI22_X1 U1179 ( .A1(n307), .A2(n242), .B1(n339), .B2(n239), .ZN(n1944) );
  OAI22_X1 U1180 ( .A1(n434), .A2(n254), .B1(n466), .B2(n251), .ZN(n1926) );
  OAI22_X1 U1181 ( .A1(n306), .A2(n242), .B1(n338), .B2(n239), .ZN(n1927) );
  OAI22_X1 U1182 ( .A1(n433), .A2(n254), .B1(n465), .B2(n251), .ZN(n1909) );
  OAI22_X1 U1183 ( .A1(n305), .A2(n242), .B1(n337), .B2(n239), .ZN(n1910) );
  OAI22_X1 U1184 ( .A1(n432), .A2(n254), .B1(n464), .B2(n251), .ZN(n1892) );
  OAI22_X1 U1185 ( .A1(n304), .A2(n242), .B1(n336), .B2(n239), .ZN(n1893) );
  OAI22_X1 U1186 ( .A1(n431), .A2(n254), .B1(n463), .B2(n251), .ZN(n1875) );
  OAI22_X1 U1187 ( .A1(n303), .A2(n242), .B1(n335), .B2(n239), .ZN(n1876) );
  OAI22_X1 U1188 ( .A1(n430), .A2(n254), .B1(n462), .B2(n251), .ZN(n1858) );
  OAI22_X1 U1189 ( .A1(n302), .A2(n242), .B1(n334), .B2(n239), .ZN(n1859) );
  OAI22_X1 U1190 ( .A1(n429), .A2(n254), .B1(n461), .B2(n251), .ZN(n1841) );
  OAI22_X1 U1191 ( .A1(n301), .A2(n242), .B1(n333), .B2(n239), .ZN(n1842) );
  OAI22_X1 U1192 ( .A1(n428), .A2(n254), .B1(n460), .B2(n251), .ZN(n1824) );
  OAI22_X1 U1193 ( .A1(n300), .A2(n242), .B1(n332), .B2(n239), .ZN(n1825) );
  OAI22_X1 U1194 ( .A1(n427), .A2(n254), .B1(n459), .B2(n251), .ZN(n1807) );
  OAI22_X1 U1195 ( .A1(n299), .A2(n242), .B1(n331), .B2(n239), .ZN(n1808) );
  OAI22_X1 U1196 ( .A1(n426), .A2(n254), .B1(n458), .B2(n251), .ZN(n1790) );
  OAI22_X1 U1197 ( .A1(n298), .A2(n242), .B1(n330), .B2(n239), .ZN(n1791) );
  OAI22_X1 U1198 ( .A1(n425), .A2(n254), .B1(n457), .B2(n251), .ZN(n1773) );
  OAI22_X1 U1199 ( .A1(n297), .A2(n242), .B1(n329), .B2(n239), .ZN(n1774) );
  OAI22_X1 U1200 ( .A1(n320), .A2(n20), .B1(n352), .B2(n17), .ZN(n2771) );
  OAI22_X1 U1201 ( .A1(n448), .A2(n32), .B1(n480), .B2(n29), .ZN(n2768) );
  OAI22_X1 U1202 ( .A1(n319), .A2(n20), .B1(n351), .B2(n17), .ZN(n2739) );
  OAI22_X1 U1203 ( .A1(n447), .A2(n32), .B1(n479), .B2(n29), .ZN(n2738) );
  OAI22_X1 U1204 ( .A1(n318), .A2(n20), .B1(n350), .B2(n17), .ZN(n2722) );
  OAI22_X1 U1205 ( .A1(n446), .A2(n32), .B1(n478), .B2(n29), .ZN(n2721) );
  OAI22_X1 U1206 ( .A1(n317), .A2(n20), .B1(n349), .B2(n17), .ZN(n2705) );
  OAI22_X1 U1207 ( .A1(n445), .A2(n32), .B1(n477), .B2(n29), .ZN(n2704) );
  OAI22_X1 U1208 ( .A1(n316), .A2(n20), .B1(n348), .B2(n17), .ZN(n2688) );
  OAI22_X1 U1209 ( .A1(n444), .A2(n32), .B1(n476), .B2(n29), .ZN(n2687) );
  OAI22_X1 U1210 ( .A1(n315), .A2(n20), .B1(n347), .B2(n17), .ZN(n2671) );
  OAI22_X1 U1211 ( .A1(n443), .A2(n32), .B1(n475), .B2(n29), .ZN(n2670) );
  OAI22_X1 U1212 ( .A1(n314), .A2(n20), .B1(n346), .B2(n17), .ZN(n2654) );
  OAI22_X1 U1213 ( .A1(n442), .A2(n32), .B1(n474), .B2(n29), .ZN(n2653) );
  OAI22_X1 U1214 ( .A1(n313), .A2(n20), .B1(n345), .B2(n17), .ZN(n2637) );
  OAI22_X1 U1215 ( .A1(n441), .A2(n32), .B1(n473), .B2(n29), .ZN(n2636) );
  OAI22_X1 U1216 ( .A1(n312), .A2(n20), .B1(n344), .B2(n17), .ZN(n2620) );
  OAI22_X1 U1217 ( .A1(n440), .A2(n32), .B1(n472), .B2(n29), .ZN(n2619) );
  OAI22_X1 U1218 ( .A1(n311), .A2(n20), .B1(n343), .B2(n17), .ZN(n2603) );
  OAI22_X1 U1219 ( .A1(n439), .A2(n32), .B1(n471), .B2(n29), .ZN(n2602) );
  OAI22_X1 U1220 ( .A1(n310), .A2(n20), .B1(n342), .B2(n17), .ZN(n2586) );
  OAI22_X1 U1221 ( .A1(n438), .A2(n32), .B1(n470), .B2(n29), .ZN(n2585) );
  OAI22_X1 U1222 ( .A1(n309), .A2(n20), .B1(n341), .B2(n17), .ZN(n2569) );
  OAI22_X1 U1223 ( .A1(n437), .A2(n32), .B1(n469), .B2(n29), .ZN(n2568) );
  OAI22_X1 U1224 ( .A1(n308), .A2(n21), .B1(n340), .B2(n18), .ZN(n2552) );
  OAI22_X1 U1225 ( .A1(n436), .A2(n161), .B1(n468), .B2(n30), .ZN(n2551) );
  OAI22_X1 U1226 ( .A1(n307), .A2(n21), .B1(n339), .B2(n18), .ZN(n2535) );
  OAI22_X1 U1227 ( .A1(n435), .A2(n161), .B1(n467), .B2(n30), .ZN(n2534) );
  OAI22_X1 U1228 ( .A1(n306), .A2(n21), .B1(n338), .B2(n18), .ZN(n2518) );
  OAI22_X1 U1229 ( .A1(n434), .A2(n161), .B1(n466), .B2(n30), .ZN(n2517) );
  OAI22_X1 U1230 ( .A1(n305), .A2(n21), .B1(n337), .B2(n18), .ZN(n2501) );
  OAI22_X1 U1231 ( .A1(n433), .A2(n161), .B1(n465), .B2(n30), .ZN(n2500) );
  OAI22_X1 U1232 ( .A1(n304), .A2(n21), .B1(n336), .B2(n18), .ZN(n2484) );
  OAI22_X1 U1233 ( .A1(n432), .A2(n161), .B1(n464), .B2(n30), .ZN(n2483) );
  OAI22_X1 U1234 ( .A1(n303), .A2(n21), .B1(n335), .B2(n18), .ZN(n2467) );
  OAI22_X1 U1235 ( .A1(n431), .A2(n161), .B1(n463), .B2(n30), .ZN(n2466) );
  OAI22_X1 U1236 ( .A1(n302), .A2(n21), .B1(n334), .B2(n18), .ZN(n2450) );
  OAI22_X1 U1237 ( .A1(n430), .A2(n161), .B1(n462), .B2(n30), .ZN(n2449) );
  OAI22_X1 U1238 ( .A1(n301), .A2(n21), .B1(n333), .B2(n18), .ZN(n2433) );
  OAI22_X1 U1239 ( .A1(n429), .A2(n161), .B1(n461), .B2(n30), .ZN(n2432) );
  OAI22_X1 U1240 ( .A1(n300), .A2(n21), .B1(n332), .B2(n18), .ZN(n2416) );
  OAI22_X1 U1241 ( .A1(n428), .A2(n161), .B1(n460), .B2(n30), .ZN(n2415) );
  OAI22_X1 U1242 ( .A1(n299), .A2(n21), .B1(n331), .B2(n18), .ZN(n2399) );
  OAI22_X1 U1243 ( .A1(n427), .A2(n161), .B1(n459), .B2(n30), .ZN(n2398) );
  OAI22_X1 U1244 ( .A1(n298), .A2(n21), .B1(n330), .B2(n18), .ZN(n2382) );
  OAI22_X1 U1245 ( .A1(n426), .A2(n161), .B1(n458), .B2(n30), .ZN(n2381) );
  OAI22_X1 U1246 ( .A1(n297), .A2(n21), .B1(n329), .B2(n18), .ZN(n2365) );
  OAI22_X1 U1247 ( .A1(n425), .A2(n161), .B1(n457), .B2(n30), .ZN(n2364) );
  OAI22_X1 U1248 ( .A1(n40), .A2(n279), .B1(n72), .B2(n276), .ZN(n1754) );
  OAI22_X1 U1249 ( .A1(n39), .A2(n279), .B1(n71), .B2(n276), .ZN(n1737) );
  OAI22_X1 U1250 ( .A1(n38), .A2(n279), .B1(n70), .B2(n276), .ZN(n1720) );
  OAI22_X1 U1251 ( .A1(n37), .A2(n279), .B1(n69), .B2(n276), .ZN(n1703) );
  OAI22_X1 U1252 ( .A1(n36), .A2(n279), .B1(n68), .B2(n276), .ZN(n1686) );
  OAI22_X1 U1253 ( .A1(n35), .A2(n279), .B1(n67), .B2(n276), .ZN(n1669) );
  OAI22_X1 U1254 ( .A1(n34), .A2(n279), .B1(n66), .B2(n276), .ZN(n1652) );
  OAI22_X1 U1255 ( .A1(n33), .A2(n279), .B1(n65), .B2(n276), .ZN(n1621) );
  OAI22_X1 U1256 ( .A1(n40), .A2(n186), .B1(n72), .B2(n183), .ZN(n2345) );
  OAI22_X1 U1257 ( .A1(n39), .A2(n186), .B1(n71), .B2(n183), .ZN(n2328) );
  OAI22_X1 U1258 ( .A1(n38), .A2(n186), .B1(n70), .B2(n183), .ZN(n2311) );
  OAI22_X1 U1259 ( .A1(n37), .A2(n186), .B1(n69), .B2(n183), .ZN(n2294) );
  OAI22_X1 U1260 ( .A1(n36), .A2(n186), .B1(n68), .B2(n183), .ZN(n2277) );
  OAI22_X1 U1261 ( .A1(n35), .A2(n186), .B1(n67), .B2(n183), .ZN(n2260) );
  OAI22_X1 U1262 ( .A1(n34), .A2(n186), .B1(n66), .B2(n183), .ZN(n2243) );
  OAI22_X1 U1263 ( .A1(n33), .A2(n186), .B1(n65), .B2(n183), .ZN(n2212) );
  OAI22_X1 U1264 ( .A1(n64), .A2(n277), .B1(n96), .B2(n274), .ZN(n2172) );
  OAI22_X1 U1265 ( .A1(n63), .A2(n277), .B1(n95), .B2(n274), .ZN(n2145) );
  OAI22_X1 U1266 ( .A1(n62), .A2(n277), .B1(n94), .B2(n274), .ZN(n2128) );
  OAI22_X1 U1267 ( .A1(n61), .A2(n277), .B1(n93), .B2(n274), .ZN(n2111) );
  OAI22_X1 U1268 ( .A1(n60), .A2(n277), .B1(n92), .B2(n274), .ZN(n2094) );
  OAI22_X1 U1269 ( .A1(n59), .A2(n277), .B1(n91), .B2(n274), .ZN(n2077) );
  OAI22_X1 U1270 ( .A1(n58), .A2(n277), .B1(n90), .B2(n274), .ZN(n2060) );
  OAI22_X1 U1271 ( .A1(n57), .A2(n277), .B1(n89), .B2(n274), .ZN(n2043) );
  OAI22_X1 U1272 ( .A1(n56), .A2(n277), .B1(n88), .B2(n274), .ZN(n2026) );
  OAI22_X1 U1273 ( .A1(n55), .A2(n277), .B1(n87), .B2(n274), .ZN(n2009) );
  OAI22_X1 U1274 ( .A1(n54), .A2(n277), .B1(n86), .B2(n274), .ZN(n1992) );
  OAI22_X1 U1275 ( .A1(n53), .A2(n277), .B1(n85), .B2(n274), .ZN(n1975) );
  OAI22_X1 U1276 ( .A1(n52), .A2(n278), .B1(n84), .B2(n275), .ZN(n1958) );
  OAI22_X1 U1277 ( .A1(n51), .A2(n278), .B1(n83), .B2(n275), .ZN(n1941) );
  OAI22_X1 U1278 ( .A1(n50), .A2(n278), .B1(n82), .B2(n275), .ZN(n1924) );
  OAI22_X1 U1279 ( .A1(n49), .A2(n278), .B1(n81), .B2(n275), .ZN(n1907) );
  OAI22_X1 U1280 ( .A1(n48), .A2(n278), .B1(n80), .B2(n275), .ZN(n1890) );
  OAI22_X1 U1281 ( .A1(n47), .A2(n278), .B1(n79), .B2(n275), .ZN(n1873) );
  OAI22_X1 U1282 ( .A1(n46), .A2(n278), .B1(n78), .B2(n275), .ZN(n1856) );
  OAI22_X1 U1283 ( .A1(n45), .A2(n278), .B1(n77), .B2(n275), .ZN(n1839) );
  OAI22_X1 U1284 ( .A1(n44), .A2(n278), .B1(n76), .B2(n275), .ZN(n1822) );
  OAI22_X1 U1285 ( .A1(n43), .A2(n278), .B1(n75), .B2(n275), .ZN(n1805) );
  OAI22_X1 U1286 ( .A1(n42), .A2(n278), .B1(n74), .B2(n275), .ZN(n1788) );
  OAI22_X1 U1287 ( .A1(n41), .A2(n278), .B1(n73), .B2(n275), .ZN(n1771) );
  OAI22_X1 U1288 ( .A1(n64), .A2(n184), .B1(n96), .B2(n181), .ZN(n2763) );
  OAI22_X1 U1289 ( .A1(n63), .A2(n184), .B1(n95), .B2(n181), .ZN(n2736) );
  OAI22_X1 U1290 ( .A1(n62), .A2(n184), .B1(n94), .B2(n181), .ZN(n2719) );
  OAI22_X1 U1291 ( .A1(n61), .A2(n184), .B1(n93), .B2(n181), .ZN(n2702) );
  OAI22_X1 U1292 ( .A1(n60), .A2(n184), .B1(n92), .B2(n181), .ZN(n2685) );
  OAI22_X1 U1293 ( .A1(n59), .A2(n184), .B1(n91), .B2(n181), .ZN(n2668) );
  OAI22_X1 U1294 ( .A1(n58), .A2(n184), .B1(n90), .B2(n181), .ZN(n2651) );
  OAI22_X1 U1295 ( .A1(n57), .A2(n184), .B1(n89), .B2(n181), .ZN(n2634) );
  OAI22_X1 U1296 ( .A1(n56), .A2(n184), .B1(n88), .B2(n181), .ZN(n2617) );
  OAI22_X1 U1297 ( .A1(n55), .A2(n184), .B1(n87), .B2(n181), .ZN(n2600) );
  OAI22_X1 U1298 ( .A1(n54), .A2(n184), .B1(n86), .B2(n181), .ZN(n2583) );
  OAI22_X1 U1299 ( .A1(n53), .A2(n184), .B1(n85), .B2(n181), .ZN(n2566) );
  OAI22_X1 U1300 ( .A1(n52), .A2(n185), .B1(n84), .B2(n182), .ZN(n2549) );
  OAI22_X1 U1301 ( .A1(n51), .A2(n185), .B1(n83), .B2(n182), .ZN(n2532) );
  OAI22_X1 U1302 ( .A1(n50), .A2(n185), .B1(n82), .B2(n182), .ZN(n2515) );
  OAI22_X1 U1303 ( .A1(n49), .A2(n185), .B1(n81), .B2(n182), .ZN(n2498) );
  OAI22_X1 U1304 ( .A1(n48), .A2(n185), .B1(n80), .B2(n182), .ZN(n2481) );
  OAI22_X1 U1305 ( .A1(n47), .A2(n185), .B1(n79), .B2(n182), .ZN(n2464) );
  OAI22_X1 U1306 ( .A1(n46), .A2(n185), .B1(n78), .B2(n182), .ZN(n2447) );
  OAI22_X1 U1307 ( .A1(n45), .A2(n185), .B1(n77), .B2(n182), .ZN(n2430) );
  OAI22_X1 U1308 ( .A1(n44), .A2(n185), .B1(n76), .B2(n182), .ZN(n2413) );
  OAI22_X1 U1309 ( .A1(n43), .A2(n185), .B1(n75), .B2(n182), .ZN(n2396) );
  OAI22_X1 U1310 ( .A1(n42), .A2(n185), .B1(n74), .B2(n182), .ZN(n2379) );
  OAI22_X1 U1311 ( .A1(n41), .A2(n185), .B1(n73), .B2(n182), .ZN(n2362) );
  OAI22_X1 U1312 ( .A1(n3844), .A2(n795), .B1(n796), .B2(n992), .ZN(n2773) );
  OAI22_X1 U1313 ( .A1(n3843), .A2(n794), .B1(n796), .B2(n991), .ZN(n2774) );
  OAI22_X1 U1314 ( .A1(n3842), .A2(n795), .B1(n796), .B2(n990), .ZN(n2775) );
  OAI22_X1 U1315 ( .A1(n3841), .A2(n794), .B1(n796), .B2(n989), .ZN(n2776) );
  OAI22_X1 U1316 ( .A1(n3840), .A2(n795), .B1(n796), .B2(n988), .ZN(n2777) );
  OAI22_X1 U1317 ( .A1(n3839), .A2(n794), .B1(n797), .B2(n987), .ZN(n2778) );
  OAI22_X1 U1318 ( .A1(n3838), .A2(n795), .B1(n797), .B2(n986), .ZN(n2779) );
  OAI22_X1 U1319 ( .A1(n3837), .A2(n794), .B1(n797), .B2(n985), .ZN(n2780) );
  OAI22_X1 U1320 ( .A1(n3836), .A2(n795), .B1(n797), .B2(n984), .ZN(n2781) );
  OAI22_X1 U1321 ( .A1(n3835), .A2(n795), .B1(n797), .B2(n983), .ZN(n2782) );
  OAI22_X1 U1322 ( .A1(n3834), .A2(n795), .B1(n798), .B2(n982), .ZN(n2783) );
  OAI22_X1 U1323 ( .A1(n3833), .A2(n795), .B1(n798), .B2(n981), .ZN(n2784) );
  OAI22_X1 U1324 ( .A1(n3832), .A2(n795), .B1(n798), .B2(n980), .ZN(n2785) );
  OAI22_X1 U1325 ( .A1(n3831), .A2(n795), .B1(n798), .B2(n979), .ZN(n2786) );
  OAI22_X1 U1326 ( .A1(n3830), .A2(n795), .B1(n798), .B2(n978), .ZN(n2787) );
  OAI22_X1 U1327 ( .A1(n3829), .A2(n795), .B1(n799), .B2(n977), .ZN(n2788) );
  OAI22_X1 U1328 ( .A1(n3828), .A2(n795), .B1(n799), .B2(n976), .ZN(n2789) );
  OAI22_X1 U1329 ( .A1(n3827), .A2(n795), .B1(n799), .B2(n975), .ZN(n2790) );
  OAI22_X1 U1330 ( .A1(n3826), .A2(n795), .B1(n799), .B2(n974), .ZN(n2791) );
  OAI22_X1 U1331 ( .A1(n3825), .A2(n795), .B1(n799), .B2(n973), .ZN(n2792) );
  OAI22_X1 U1332 ( .A1(n3824), .A2(n794), .B1(n800), .B2(n972), .ZN(n2793) );
  OAI22_X1 U1333 ( .A1(n3823), .A2(n794), .B1(n800), .B2(n971), .ZN(n2794) );
  OAI22_X1 U1334 ( .A1(n3822), .A2(n794), .B1(n800), .B2(n970), .ZN(n2795) );
  OAI22_X1 U1335 ( .A1(n3844), .A2(n786), .B1(n787), .B2(n960), .ZN(n2805) );
  OAI22_X1 U1336 ( .A1(n3843), .A2(n785), .B1(n787), .B2(n959), .ZN(n2806) );
  OAI22_X1 U1337 ( .A1(n3842), .A2(n786), .B1(n787), .B2(n958), .ZN(n2807) );
  OAI22_X1 U1338 ( .A1(n3841), .A2(n785), .B1(n787), .B2(n957), .ZN(n2808) );
  OAI22_X1 U1339 ( .A1(n3840), .A2(n786), .B1(n787), .B2(n956), .ZN(n2809) );
  OAI22_X1 U1340 ( .A1(n3839), .A2(n785), .B1(n788), .B2(n955), .ZN(n2810) );
  OAI22_X1 U1341 ( .A1(n3838), .A2(n786), .B1(n788), .B2(n954), .ZN(n2811) );
  OAI22_X1 U1342 ( .A1(n3837), .A2(n785), .B1(n788), .B2(n953), .ZN(n2812) );
  OAI22_X1 U1343 ( .A1(n3836), .A2(n786), .B1(n788), .B2(n952), .ZN(n2813) );
  OAI22_X1 U1344 ( .A1(n3835), .A2(n786), .B1(n788), .B2(n951), .ZN(n2814) );
  OAI22_X1 U1345 ( .A1(n3834), .A2(n786), .B1(n789), .B2(n950), .ZN(n2815) );
  OAI22_X1 U1346 ( .A1(n3833), .A2(n786), .B1(n789), .B2(n949), .ZN(n2816) );
  OAI22_X1 U1347 ( .A1(n3832), .A2(n786), .B1(n789), .B2(n948), .ZN(n2817) );
  OAI22_X1 U1348 ( .A1(n3831), .A2(n786), .B1(n789), .B2(n947), .ZN(n2818) );
  OAI22_X1 U1349 ( .A1(n3830), .A2(n786), .B1(n789), .B2(n946), .ZN(n2819) );
  OAI22_X1 U1350 ( .A1(n3829), .A2(n786), .B1(n790), .B2(n945), .ZN(n2820) );
  OAI22_X1 U1351 ( .A1(n3828), .A2(n786), .B1(n790), .B2(n944), .ZN(n2821) );
  OAI22_X1 U1352 ( .A1(n3827), .A2(n786), .B1(n790), .B2(n943), .ZN(n2822) );
  OAI22_X1 U1353 ( .A1(n3826), .A2(n786), .B1(n790), .B2(n942), .ZN(n2823) );
  OAI22_X1 U1354 ( .A1(n3825), .A2(n786), .B1(n790), .B2(n941), .ZN(n2824) );
  OAI22_X1 U1355 ( .A1(n3824), .A2(n785), .B1(n791), .B2(n940), .ZN(n2825) );
  OAI22_X1 U1356 ( .A1(n3823), .A2(n785), .B1(n791), .B2(n939), .ZN(n2826) );
  OAI22_X1 U1357 ( .A1(n3822), .A2(n785), .B1(n791), .B2(n938), .ZN(n2827) );
  OAI22_X1 U1358 ( .A1(n3844), .A2(n759), .B1(n760), .B2(n864), .ZN(n2837) );
  OAI22_X1 U1359 ( .A1(n3843), .A2(n758), .B1(n760), .B2(n863), .ZN(n2838) );
  OAI22_X1 U1360 ( .A1(n3842), .A2(n759), .B1(n760), .B2(n862), .ZN(n2839) );
  OAI22_X1 U1361 ( .A1(n3841), .A2(n758), .B1(n760), .B2(n861), .ZN(n2840) );
  OAI22_X1 U1362 ( .A1(n3840), .A2(n759), .B1(n760), .B2(n860), .ZN(n2841) );
  OAI22_X1 U1363 ( .A1(n3839), .A2(n758), .B1(n761), .B2(n859), .ZN(n2842) );
  OAI22_X1 U1364 ( .A1(n3838), .A2(n759), .B1(n761), .B2(n858), .ZN(n2843) );
  OAI22_X1 U1365 ( .A1(n3837), .A2(n758), .B1(n761), .B2(n857), .ZN(n2844) );
  OAI22_X1 U1366 ( .A1(n3836), .A2(n759), .B1(n761), .B2(n856), .ZN(n2845) );
  OAI22_X1 U1367 ( .A1(n3835), .A2(n759), .B1(n761), .B2(n855), .ZN(n2846) );
  OAI22_X1 U1368 ( .A1(n3834), .A2(n759), .B1(n762), .B2(n854), .ZN(n2847) );
  OAI22_X1 U1369 ( .A1(n3833), .A2(n759), .B1(n762), .B2(n853), .ZN(n2848) );
  OAI22_X1 U1370 ( .A1(n3832), .A2(n759), .B1(n762), .B2(n852), .ZN(n2849) );
  OAI22_X1 U1371 ( .A1(n3831), .A2(n759), .B1(n762), .B2(n851), .ZN(n2850) );
  OAI22_X1 U1372 ( .A1(n3830), .A2(n759), .B1(n762), .B2(n850), .ZN(n2851) );
  OAI22_X1 U1373 ( .A1(n3829), .A2(n759), .B1(n763), .B2(n849), .ZN(n2852) );
  OAI22_X1 U1374 ( .A1(n3828), .A2(n759), .B1(n763), .B2(n848), .ZN(n2853) );
  OAI22_X1 U1375 ( .A1(n3827), .A2(n759), .B1(n763), .B2(n847), .ZN(n2854) );
  OAI22_X1 U1376 ( .A1(n3826), .A2(n759), .B1(n763), .B2(n846), .ZN(n2855) );
  OAI22_X1 U1377 ( .A1(n3825), .A2(n759), .B1(n763), .B2(n845), .ZN(n2856) );
  OAI22_X1 U1378 ( .A1(n3824), .A2(n758), .B1(n764), .B2(n844), .ZN(n2857) );
  OAI22_X1 U1379 ( .A1(n3823), .A2(n758), .B1(n764), .B2(n843), .ZN(n2858) );
  OAI22_X1 U1380 ( .A1(n3822), .A2(n758), .B1(n764), .B2(n842), .ZN(n2859) );
  OAI22_X1 U1381 ( .A1(n3844), .A2(n750), .B1(n751), .B2(n832), .ZN(n2869) );
  OAI22_X1 U1382 ( .A1(n3843), .A2(n749), .B1(n751), .B2(n831), .ZN(n2870) );
  OAI22_X1 U1383 ( .A1(n3842), .A2(n750), .B1(n751), .B2(n830), .ZN(n2871) );
  OAI22_X1 U1384 ( .A1(n3841), .A2(n749), .B1(n751), .B2(n829), .ZN(n2872) );
  OAI22_X1 U1385 ( .A1(n3840), .A2(n750), .B1(n751), .B2(n828), .ZN(n2873) );
  OAI22_X1 U1386 ( .A1(n3839), .A2(n749), .B1(n752), .B2(n827), .ZN(n2874) );
  OAI22_X1 U1387 ( .A1(n3838), .A2(n750), .B1(n752), .B2(n826), .ZN(n2875) );
  OAI22_X1 U1388 ( .A1(n3837), .A2(n749), .B1(n752), .B2(n825), .ZN(n2876) );
  OAI22_X1 U1389 ( .A1(n3836), .A2(n750), .B1(n752), .B2(n824), .ZN(n2877) );
  OAI22_X1 U1390 ( .A1(n3835), .A2(n750), .B1(n752), .B2(n823), .ZN(n2878) );
  OAI22_X1 U1391 ( .A1(n3834), .A2(n750), .B1(n753), .B2(n822), .ZN(n2879) );
  OAI22_X1 U1392 ( .A1(n3833), .A2(n750), .B1(n753), .B2(n821), .ZN(n2880) );
  OAI22_X1 U1393 ( .A1(n3832), .A2(n750), .B1(n753), .B2(n820), .ZN(n2881) );
  OAI22_X1 U1394 ( .A1(n3831), .A2(n750), .B1(n753), .B2(n819), .ZN(n2882) );
  OAI22_X1 U1395 ( .A1(n3830), .A2(n750), .B1(n753), .B2(n818), .ZN(n2883) );
  OAI22_X1 U1396 ( .A1(n3829), .A2(n750), .B1(n754), .B2(n817), .ZN(n2884) );
  OAI22_X1 U1397 ( .A1(n3828), .A2(n750), .B1(n754), .B2(n816), .ZN(n2885) );
  OAI22_X1 U1398 ( .A1(n3827), .A2(n750), .B1(n754), .B2(n815), .ZN(n2886) );
  OAI22_X1 U1399 ( .A1(n3826), .A2(n750), .B1(n754), .B2(n814), .ZN(n2887) );
  OAI22_X1 U1400 ( .A1(n3825), .A2(n750), .B1(n754), .B2(n813), .ZN(n2888) );
  OAI22_X1 U1401 ( .A1(n3824), .A2(n749), .B1(n755), .B2(n812), .ZN(n2889) );
  OAI22_X1 U1402 ( .A1(n3823), .A2(n749), .B1(n755), .B2(n811), .ZN(n2890) );
  OAI22_X1 U1403 ( .A1(n3822), .A2(n749), .B1(n755), .B2(n810), .ZN(n2891) );
  OAI22_X1 U1404 ( .A1(n3844), .A2(n705), .B1(n706), .B2(n672), .ZN(n2901) );
  OAI22_X1 U1405 ( .A1(n3843), .A2(n704), .B1(n706), .B2(n671), .ZN(n2902) );
  OAI22_X1 U1406 ( .A1(n3842), .A2(n705), .B1(n706), .B2(n670), .ZN(n2903) );
  OAI22_X1 U1407 ( .A1(n3841), .A2(n704), .B1(n706), .B2(n669), .ZN(n2904) );
  OAI22_X1 U1408 ( .A1(n3840), .A2(n705), .B1(n706), .B2(n668), .ZN(n2905) );
  OAI22_X1 U1409 ( .A1(n3839), .A2(n704), .B1(n707), .B2(n667), .ZN(n2906) );
  OAI22_X1 U1410 ( .A1(n3838), .A2(n705), .B1(n707), .B2(n666), .ZN(n2907) );
  OAI22_X1 U1411 ( .A1(n3837), .A2(n704), .B1(n707), .B2(n665), .ZN(n2908) );
  OAI22_X1 U1412 ( .A1(n3836), .A2(n705), .B1(n707), .B2(n664), .ZN(n2909) );
  OAI22_X1 U1413 ( .A1(n3835), .A2(n705), .B1(n707), .B2(n663), .ZN(n2910) );
  OAI22_X1 U1414 ( .A1(n3834), .A2(n705), .B1(n708), .B2(n662), .ZN(n2911) );
  OAI22_X1 U1415 ( .A1(n3833), .A2(n705), .B1(n708), .B2(n661), .ZN(n2912) );
  OAI22_X1 U1416 ( .A1(n3832), .A2(n705), .B1(n708), .B2(n660), .ZN(n2913) );
  OAI22_X1 U1417 ( .A1(n3831), .A2(n705), .B1(n708), .B2(n659), .ZN(n2914) );
  OAI22_X1 U1418 ( .A1(n3830), .A2(n705), .B1(n708), .B2(n658), .ZN(n2915) );
  OAI22_X1 U1419 ( .A1(n3829), .A2(n705), .B1(n709), .B2(n657), .ZN(n2916) );
  OAI22_X1 U1420 ( .A1(n3828), .A2(n705), .B1(n709), .B2(n656), .ZN(n2917) );
  OAI22_X1 U1421 ( .A1(n3827), .A2(n705), .B1(n709), .B2(n655), .ZN(n2918) );
  OAI22_X1 U1422 ( .A1(n3826), .A2(n705), .B1(n709), .B2(n654), .ZN(n2919) );
  OAI22_X1 U1423 ( .A1(n3825), .A2(n705), .B1(n709), .B2(n653), .ZN(n2920) );
  OAI22_X1 U1424 ( .A1(n3824), .A2(n704), .B1(n710), .B2(n652), .ZN(n2921) );
  OAI22_X1 U1425 ( .A1(n3823), .A2(n704), .B1(n710), .B2(n651), .ZN(n2922) );
  OAI22_X1 U1426 ( .A1(n3822), .A2(n704), .B1(n710), .B2(n650), .ZN(n2923) );
  OAI22_X1 U1427 ( .A1(n3844), .A2(n696), .B1(n697), .B2(n640), .ZN(n2933) );
  OAI22_X1 U1428 ( .A1(n3843), .A2(n695), .B1(n697), .B2(n639), .ZN(n2934) );
  OAI22_X1 U1429 ( .A1(n3842), .A2(n696), .B1(n697), .B2(n638), .ZN(n2935) );
  OAI22_X1 U1430 ( .A1(n3841), .A2(n695), .B1(n697), .B2(n637), .ZN(n2936) );
  OAI22_X1 U1431 ( .A1(n3840), .A2(n696), .B1(n697), .B2(n636), .ZN(n2937) );
  OAI22_X1 U1432 ( .A1(n3839), .A2(n695), .B1(n698), .B2(n635), .ZN(n2938) );
  OAI22_X1 U1433 ( .A1(n3838), .A2(n696), .B1(n698), .B2(n634), .ZN(n2939) );
  OAI22_X1 U1434 ( .A1(n3837), .A2(n695), .B1(n698), .B2(n633), .ZN(n2940) );
  OAI22_X1 U1435 ( .A1(n3836), .A2(n696), .B1(n698), .B2(n632), .ZN(n2941) );
  OAI22_X1 U1436 ( .A1(n3835), .A2(n696), .B1(n698), .B2(n631), .ZN(n2942) );
  OAI22_X1 U1437 ( .A1(n3834), .A2(n696), .B1(n699), .B2(n630), .ZN(n2943) );
  OAI22_X1 U1438 ( .A1(n3833), .A2(n696), .B1(n699), .B2(n629), .ZN(n2944) );
  OAI22_X1 U1439 ( .A1(n3832), .A2(n696), .B1(n699), .B2(n628), .ZN(n2945) );
  OAI22_X1 U1440 ( .A1(n3831), .A2(n696), .B1(n699), .B2(n627), .ZN(n2946) );
  OAI22_X1 U1441 ( .A1(n3830), .A2(n696), .B1(n699), .B2(n626), .ZN(n2947) );
  OAI22_X1 U1442 ( .A1(n3829), .A2(n696), .B1(n700), .B2(n625), .ZN(n2948) );
  OAI22_X1 U1443 ( .A1(n3828), .A2(n696), .B1(n700), .B2(n624), .ZN(n2949) );
  OAI22_X1 U1444 ( .A1(n3827), .A2(n696), .B1(n700), .B2(n623), .ZN(n2950) );
  OAI22_X1 U1445 ( .A1(n3826), .A2(n696), .B1(n700), .B2(n622), .ZN(n2951) );
  OAI22_X1 U1446 ( .A1(n3825), .A2(n696), .B1(n700), .B2(n621), .ZN(n2952) );
  OAI22_X1 U1447 ( .A1(n3824), .A2(n695), .B1(n701), .B2(n620), .ZN(n2953) );
  OAI22_X1 U1448 ( .A1(n3823), .A2(n695), .B1(n701), .B2(n619), .ZN(n2954) );
  OAI22_X1 U1449 ( .A1(n3822), .A2(n695), .B1(n701), .B2(n618), .ZN(n2955) );
  OAI22_X1 U1450 ( .A1(n3844), .A2(n605), .B1(n606), .B2(n544), .ZN(n2965) );
  OAI22_X1 U1451 ( .A1(n3843), .A2(n604), .B1(n606), .B2(n543), .ZN(n2966) );
  OAI22_X1 U1452 ( .A1(n3842), .A2(n605), .B1(n606), .B2(n542), .ZN(n2967) );
  OAI22_X1 U1453 ( .A1(n3841), .A2(n604), .B1(n606), .B2(n541), .ZN(n2968) );
  OAI22_X1 U1454 ( .A1(n3840), .A2(n605), .B1(n606), .B2(n540), .ZN(n2969) );
  OAI22_X1 U1455 ( .A1(n3839), .A2(n604), .B1(n607), .B2(n539), .ZN(n2970) );
  OAI22_X1 U1456 ( .A1(n3838), .A2(n605), .B1(n607), .B2(n538), .ZN(n2971) );
  OAI22_X1 U1457 ( .A1(n3837), .A2(n604), .B1(n607), .B2(n537), .ZN(n2972) );
  OAI22_X1 U1458 ( .A1(n3836), .A2(n605), .B1(n607), .B2(n536), .ZN(n2973) );
  OAI22_X1 U1459 ( .A1(n3835), .A2(n605), .B1(n607), .B2(n535), .ZN(n2974) );
  OAI22_X1 U1460 ( .A1(n3834), .A2(n605), .B1(n608), .B2(n534), .ZN(n2975) );
  OAI22_X1 U1461 ( .A1(n3833), .A2(n605), .B1(n608), .B2(n533), .ZN(n2976) );
  OAI22_X1 U1462 ( .A1(n3832), .A2(n605), .B1(n608), .B2(n532), .ZN(n2977) );
  OAI22_X1 U1463 ( .A1(n3831), .A2(n605), .B1(n608), .B2(n531), .ZN(n2978) );
  OAI22_X1 U1464 ( .A1(n3830), .A2(n605), .B1(n608), .B2(n530), .ZN(n2979) );
  OAI22_X1 U1465 ( .A1(n3829), .A2(n605), .B1(n673), .B2(n529), .ZN(n2980) );
  OAI22_X1 U1466 ( .A1(n3828), .A2(n605), .B1(n673), .B2(n528), .ZN(n2981) );
  OAI22_X1 U1467 ( .A1(n3827), .A2(n605), .B1(n673), .B2(n527), .ZN(n2982) );
  OAI22_X1 U1468 ( .A1(n3826), .A2(n605), .B1(n673), .B2(n526), .ZN(n2983) );
  OAI22_X1 U1469 ( .A1(n3825), .A2(n605), .B1(n673), .B2(n525), .ZN(n2984) );
  OAI22_X1 U1470 ( .A1(n3824), .A2(n604), .B1(n674), .B2(n524), .ZN(n2985) );
  OAI22_X1 U1471 ( .A1(n3823), .A2(n604), .B1(n674), .B2(n523), .ZN(n2986) );
  OAI22_X1 U1472 ( .A1(n3822), .A2(n604), .B1(n674), .B2(n522), .ZN(n2987) );
  OAI22_X1 U1473 ( .A1(n3844), .A2(n596), .B1(n597), .B2(n512), .ZN(n2997) );
  OAI22_X1 U1474 ( .A1(n3843), .A2(n595), .B1(n597), .B2(n511), .ZN(n2998) );
  OAI22_X1 U1475 ( .A1(n3842), .A2(n596), .B1(n597), .B2(n510), .ZN(n2999) );
  OAI22_X1 U1476 ( .A1(n3841), .A2(n595), .B1(n597), .B2(n509), .ZN(n3000) );
  OAI22_X1 U1477 ( .A1(n3840), .A2(n596), .B1(n597), .B2(n508), .ZN(n3001) );
  OAI22_X1 U1478 ( .A1(n3839), .A2(n595), .B1(n598), .B2(n507), .ZN(n3002) );
  OAI22_X1 U1479 ( .A1(n3838), .A2(n596), .B1(n598), .B2(n506), .ZN(n3003) );
  OAI22_X1 U1480 ( .A1(n3837), .A2(n595), .B1(n598), .B2(n505), .ZN(n3004) );
  OAI22_X1 U1481 ( .A1(n3836), .A2(n596), .B1(n598), .B2(n504), .ZN(n3005) );
  OAI22_X1 U1482 ( .A1(n3835), .A2(n596), .B1(n598), .B2(n503), .ZN(n3006) );
  OAI22_X1 U1483 ( .A1(n3834), .A2(n596), .B1(n599), .B2(n502), .ZN(n3007) );
  OAI22_X1 U1484 ( .A1(n3833), .A2(n596), .B1(n599), .B2(n501), .ZN(n3008) );
  OAI22_X1 U1485 ( .A1(n3832), .A2(n596), .B1(n599), .B2(n500), .ZN(n3009) );
  OAI22_X1 U1486 ( .A1(n3831), .A2(n596), .B1(n599), .B2(n499), .ZN(n3010) );
  OAI22_X1 U1487 ( .A1(n3830), .A2(n596), .B1(n599), .B2(n498), .ZN(n3011) );
  OAI22_X1 U1488 ( .A1(n3829), .A2(n596), .B1(n600), .B2(n497), .ZN(n3012) );
  OAI22_X1 U1489 ( .A1(n3828), .A2(n596), .B1(n600), .B2(n496), .ZN(n3013) );
  OAI22_X1 U1490 ( .A1(n3827), .A2(n596), .B1(n600), .B2(n495), .ZN(n3014) );
  OAI22_X1 U1491 ( .A1(n3826), .A2(n596), .B1(n600), .B2(n494), .ZN(n3015) );
  OAI22_X1 U1492 ( .A1(n3825), .A2(n596), .B1(n600), .B2(n493), .ZN(n3016) );
  OAI22_X1 U1493 ( .A1(n3824), .A2(n595), .B1(n601), .B2(n492), .ZN(n3017) );
  OAI22_X1 U1494 ( .A1(n3823), .A2(n595), .B1(n601), .B2(n491), .ZN(n3018) );
  OAI22_X1 U1495 ( .A1(n3822), .A2(n595), .B1(n601), .B2(n490), .ZN(n3019) );
  OAI22_X1 U1496 ( .A1(n3844), .A2(n587), .B1(n588), .B2(n480), .ZN(n3029) );
  OAI22_X1 U1497 ( .A1(n3843), .A2(n586), .B1(n588), .B2(n479), .ZN(n3030) );
  OAI22_X1 U1498 ( .A1(n3842), .A2(n587), .B1(n588), .B2(n478), .ZN(n3031) );
  OAI22_X1 U1499 ( .A1(n3841), .A2(n586), .B1(n588), .B2(n477), .ZN(n3032) );
  OAI22_X1 U1500 ( .A1(n3840), .A2(n587), .B1(n588), .B2(n476), .ZN(n3033) );
  OAI22_X1 U1501 ( .A1(n3839), .A2(n586), .B1(n589), .B2(n475), .ZN(n3034) );
  OAI22_X1 U1502 ( .A1(n3838), .A2(n587), .B1(n589), .B2(n474), .ZN(n3035) );
  OAI22_X1 U1503 ( .A1(n3837), .A2(n586), .B1(n589), .B2(n473), .ZN(n3036) );
  OAI22_X1 U1504 ( .A1(n3836), .A2(n587), .B1(n589), .B2(n472), .ZN(n3037) );
  OAI22_X1 U1505 ( .A1(n3835), .A2(n587), .B1(n589), .B2(n471), .ZN(n3038) );
  OAI22_X1 U1506 ( .A1(n3834), .A2(n587), .B1(n590), .B2(n470), .ZN(n3039) );
  OAI22_X1 U1507 ( .A1(n3833), .A2(n587), .B1(n590), .B2(n469), .ZN(n3040) );
  OAI22_X1 U1508 ( .A1(n3832), .A2(n587), .B1(n590), .B2(n468), .ZN(n3041) );
  OAI22_X1 U1509 ( .A1(n3831), .A2(n587), .B1(n590), .B2(n467), .ZN(n3042) );
  OAI22_X1 U1510 ( .A1(n3830), .A2(n587), .B1(n590), .B2(n466), .ZN(n3043) );
  OAI22_X1 U1511 ( .A1(n3829), .A2(n587), .B1(n591), .B2(n465), .ZN(n3044) );
  OAI22_X1 U1512 ( .A1(n3828), .A2(n587), .B1(n591), .B2(n464), .ZN(n3045) );
  OAI22_X1 U1513 ( .A1(n3827), .A2(n587), .B1(n591), .B2(n463), .ZN(n3046) );
  OAI22_X1 U1514 ( .A1(n3826), .A2(n587), .B1(n591), .B2(n462), .ZN(n3047) );
  OAI22_X1 U1515 ( .A1(n3825), .A2(n587), .B1(n591), .B2(n461), .ZN(n3048) );
  OAI22_X1 U1516 ( .A1(n3824), .A2(n586), .B1(n592), .B2(n460), .ZN(n3049) );
  OAI22_X1 U1517 ( .A1(n3823), .A2(n586), .B1(n592), .B2(n459), .ZN(n3050) );
  OAI22_X1 U1518 ( .A1(n3822), .A2(n586), .B1(n592), .B2(n458), .ZN(n3051) );
  OAI22_X1 U1519 ( .A1(n3844), .A2(n578), .B1(n579), .B2(n448), .ZN(n3061) );
  OAI22_X1 U1520 ( .A1(n3843), .A2(n577), .B1(n579), .B2(n447), .ZN(n3062) );
  OAI22_X1 U1521 ( .A1(n3842), .A2(n578), .B1(n579), .B2(n446), .ZN(n3063) );
  OAI22_X1 U1522 ( .A1(n3841), .A2(n577), .B1(n579), .B2(n445), .ZN(n3064) );
  OAI22_X1 U1523 ( .A1(n3840), .A2(n578), .B1(n579), .B2(n444), .ZN(n3065) );
  OAI22_X1 U1524 ( .A1(n3839), .A2(n577), .B1(n580), .B2(n443), .ZN(n3066) );
  OAI22_X1 U1525 ( .A1(n3838), .A2(n578), .B1(n580), .B2(n442), .ZN(n3067) );
  OAI22_X1 U1526 ( .A1(n3837), .A2(n577), .B1(n580), .B2(n441), .ZN(n3068) );
  OAI22_X1 U1527 ( .A1(n3836), .A2(n578), .B1(n580), .B2(n440), .ZN(n3069) );
  OAI22_X1 U1528 ( .A1(n3835), .A2(n578), .B1(n580), .B2(n439), .ZN(n3070) );
  OAI22_X1 U1529 ( .A1(n3834), .A2(n578), .B1(n581), .B2(n438), .ZN(n3071) );
  OAI22_X1 U1530 ( .A1(n3833), .A2(n578), .B1(n581), .B2(n437), .ZN(n3072) );
  OAI22_X1 U1531 ( .A1(n3832), .A2(n578), .B1(n581), .B2(n436), .ZN(n3073) );
  OAI22_X1 U1532 ( .A1(n3831), .A2(n578), .B1(n581), .B2(n435), .ZN(n3074) );
  OAI22_X1 U1533 ( .A1(n3830), .A2(n578), .B1(n581), .B2(n434), .ZN(n3075) );
  OAI22_X1 U1534 ( .A1(n3829), .A2(n578), .B1(n582), .B2(n433), .ZN(n3076) );
  OAI22_X1 U1535 ( .A1(n3828), .A2(n578), .B1(n582), .B2(n432), .ZN(n3077) );
  OAI22_X1 U1536 ( .A1(n3827), .A2(n578), .B1(n582), .B2(n431), .ZN(n3078) );
  OAI22_X1 U1537 ( .A1(n3826), .A2(n578), .B1(n582), .B2(n430), .ZN(n3079) );
  OAI22_X1 U1538 ( .A1(n3825), .A2(n578), .B1(n582), .B2(n429), .ZN(n3080) );
  OAI22_X1 U1539 ( .A1(n3824), .A2(n577), .B1(n583), .B2(n428), .ZN(n3081) );
  OAI22_X1 U1540 ( .A1(n3823), .A2(n577), .B1(n583), .B2(n427), .ZN(n3082) );
  OAI22_X1 U1541 ( .A1(n3822), .A2(n577), .B1(n583), .B2(n426), .ZN(n3083) );
  OAI22_X1 U1542 ( .A1(n3844), .A2(n551), .B1(n552), .B2(n352), .ZN(n3093) );
  OAI22_X1 U1543 ( .A1(n3843), .A2(n550), .B1(n552), .B2(n351), .ZN(n3094) );
  OAI22_X1 U1544 ( .A1(n3842), .A2(n551), .B1(n552), .B2(n350), .ZN(n3095) );
  OAI22_X1 U1545 ( .A1(n3841), .A2(n550), .B1(n552), .B2(n349), .ZN(n3096) );
  OAI22_X1 U1546 ( .A1(n3840), .A2(n551), .B1(n552), .B2(n348), .ZN(n3097) );
  OAI22_X1 U1547 ( .A1(n3839), .A2(n550), .B1(n553), .B2(n347), .ZN(n3098) );
  OAI22_X1 U1548 ( .A1(n3838), .A2(n551), .B1(n553), .B2(n346), .ZN(n3099) );
  OAI22_X1 U1549 ( .A1(n3837), .A2(n550), .B1(n553), .B2(n345), .ZN(n3100) );
  OAI22_X1 U1550 ( .A1(n3836), .A2(n551), .B1(n553), .B2(n344), .ZN(n3101) );
  OAI22_X1 U1551 ( .A1(n3835), .A2(n551), .B1(n553), .B2(n343), .ZN(n3102) );
  OAI22_X1 U1552 ( .A1(n3834), .A2(n551), .B1(n554), .B2(n342), .ZN(n3103) );
  OAI22_X1 U1553 ( .A1(n3833), .A2(n551), .B1(n554), .B2(n341), .ZN(n3104) );
  OAI22_X1 U1554 ( .A1(n3832), .A2(n551), .B1(n554), .B2(n340), .ZN(n3105) );
  OAI22_X1 U1555 ( .A1(n3831), .A2(n551), .B1(n554), .B2(n339), .ZN(n3106) );
  OAI22_X1 U1556 ( .A1(n3830), .A2(n551), .B1(n554), .B2(n338), .ZN(n3107) );
  OAI22_X1 U1557 ( .A1(n3829), .A2(n551), .B1(n555), .B2(n337), .ZN(n3108) );
  OAI22_X1 U1558 ( .A1(n3828), .A2(n551), .B1(n555), .B2(n336), .ZN(n3109) );
  OAI22_X1 U1559 ( .A1(n3827), .A2(n551), .B1(n555), .B2(n335), .ZN(n3110) );
  OAI22_X1 U1560 ( .A1(n3826), .A2(n551), .B1(n555), .B2(n334), .ZN(n3111) );
  OAI22_X1 U1561 ( .A1(n3825), .A2(n551), .B1(n555), .B2(n333), .ZN(n3112) );
  OAI22_X1 U1562 ( .A1(n3824), .A2(n550), .B1(n556), .B2(n332), .ZN(n3113) );
  OAI22_X1 U1563 ( .A1(n3823), .A2(n550), .B1(n556), .B2(n331), .ZN(n3114) );
  OAI22_X1 U1564 ( .A1(n3822), .A2(n550), .B1(n556), .B2(n330), .ZN(n3115) );
  OAI22_X1 U1565 ( .A1(n3844), .A2(n414), .B1(n415), .B2(n320), .ZN(n3125) );
  OAI22_X1 U1566 ( .A1(n3843), .A2(n413), .B1(n415), .B2(n319), .ZN(n3126) );
  OAI22_X1 U1567 ( .A1(n3842), .A2(n414), .B1(n415), .B2(n318), .ZN(n3127) );
  OAI22_X1 U1568 ( .A1(n3841), .A2(n413), .B1(n415), .B2(n317), .ZN(n3128) );
  OAI22_X1 U1569 ( .A1(n3840), .A2(n414), .B1(n415), .B2(n316), .ZN(n3129) );
  OAI22_X1 U1570 ( .A1(n3839), .A2(n413), .B1(n416), .B2(n315), .ZN(n3130) );
  OAI22_X1 U1571 ( .A1(n3838), .A2(n414), .B1(n416), .B2(n314), .ZN(n3131) );
  OAI22_X1 U1572 ( .A1(n3837), .A2(n413), .B1(n416), .B2(n313), .ZN(n3132) );
  OAI22_X1 U1573 ( .A1(n3836), .A2(n414), .B1(n416), .B2(n312), .ZN(n3133) );
  OAI22_X1 U1574 ( .A1(n3835), .A2(n414), .B1(n416), .B2(n311), .ZN(n3134) );
  OAI22_X1 U1575 ( .A1(n3834), .A2(n414), .B1(n545), .B2(n310), .ZN(n3135) );
  OAI22_X1 U1576 ( .A1(n3833), .A2(n414), .B1(n545), .B2(n309), .ZN(n3136) );
  OAI22_X1 U1577 ( .A1(n3832), .A2(n414), .B1(n545), .B2(n308), .ZN(n3137) );
  OAI22_X1 U1578 ( .A1(n3831), .A2(n414), .B1(n545), .B2(n307), .ZN(n3138) );
  OAI22_X1 U1579 ( .A1(n3830), .A2(n414), .B1(n545), .B2(n306), .ZN(n3139) );
  OAI22_X1 U1580 ( .A1(n3829), .A2(n414), .B1(n546), .B2(n305), .ZN(n3140) );
  OAI22_X1 U1581 ( .A1(n3828), .A2(n414), .B1(n546), .B2(n304), .ZN(n3141) );
  OAI22_X1 U1582 ( .A1(n3827), .A2(n414), .B1(n546), .B2(n303), .ZN(n3142) );
  OAI22_X1 U1583 ( .A1(n3826), .A2(n414), .B1(n546), .B2(n302), .ZN(n3143) );
  OAI22_X1 U1584 ( .A1(n3825), .A2(n414), .B1(n546), .B2(n301), .ZN(n3144) );
  OAI22_X1 U1585 ( .A1(n3824), .A2(n413), .B1(n547), .B2(n300), .ZN(n3145) );
  OAI22_X1 U1586 ( .A1(n3823), .A2(n413), .B1(n547), .B2(n299), .ZN(n3146) );
  OAI22_X1 U1587 ( .A1(n3822), .A2(n413), .B1(n547), .B2(n298), .ZN(n3147) );
  OAI22_X1 U1588 ( .A1(n3844), .A2(n904), .B1(n905), .B2(n160), .ZN(n3157) );
  OAI22_X1 U1589 ( .A1(n3843), .A2(n903), .B1(n905), .B2(n159), .ZN(n3158) );
  OAI22_X1 U1590 ( .A1(n3842), .A2(n904), .B1(n905), .B2(n158), .ZN(n3159) );
  OAI22_X1 U1591 ( .A1(n3841), .A2(n903), .B1(n905), .B2(n157), .ZN(n3160) );
  OAI22_X1 U1592 ( .A1(n3840), .A2(n904), .B1(n905), .B2(n156), .ZN(n3161) );
  OAI22_X1 U1593 ( .A1(n3839), .A2(n903), .B1(n906), .B2(n155), .ZN(n3162) );
  OAI22_X1 U1594 ( .A1(n3838), .A2(n904), .B1(n906), .B2(n154), .ZN(n3163) );
  OAI22_X1 U1595 ( .A1(n3837), .A2(n903), .B1(n906), .B2(n153), .ZN(n3164) );
  OAI22_X1 U1596 ( .A1(n3836), .A2(n904), .B1(n906), .B2(n152), .ZN(n3165) );
  OAI22_X1 U1597 ( .A1(n3835), .A2(n904), .B1(n906), .B2(n151), .ZN(n3166) );
  OAI22_X1 U1598 ( .A1(n3834), .A2(n904), .B1(n907), .B2(n150), .ZN(n3167) );
  OAI22_X1 U1599 ( .A1(n3833), .A2(n904), .B1(n907), .B2(n149), .ZN(n3168) );
  OAI22_X1 U1600 ( .A1(n3832), .A2(n904), .B1(n907), .B2(n148), .ZN(n3169) );
  OAI22_X1 U1601 ( .A1(n3831), .A2(n904), .B1(n907), .B2(n147), .ZN(n3170) );
  OAI22_X1 U1602 ( .A1(n3830), .A2(n904), .B1(n907), .B2(n146), .ZN(n3171) );
  OAI22_X1 U1603 ( .A1(n3829), .A2(n904), .B1(n908), .B2(n145), .ZN(n3172) );
  OAI22_X1 U1604 ( .A1(n3828), .A2(n904), .B1(n908), .B2(n144), .ZN(n3173) );
  OAI22_X1 U1605 ( .A1(n3827), .A2(n904), .B1(n908), .B2(n143), .ZN(n3174) );
  OAI22_X1 U1606 ( .A1(n3826), .A2(n904), .B1(n908), .B2(n142), .ZN(n3175) );
  OAI22_X1 U1607 ( .A1(n3825), .A2(n904), .B1(n908), .B2(n141), .ZN(n3176) );
  OAI22_X1 U1608 ( .A1(n3824), .A2(n903), .B1(n909), .B2(n140), .ZN(n3177) );
  OAI22_X1 U1609 ( .A1(n3823), .A2(n903), .B1(n909), .B2(n139), .ZN(n3178) );
  OAI22_X1 U1610 ( .A1(n3822), .A2(n903), .B1(n909), .B2(n138), .ZN(n3179) );
  OAI22_X1 U1611 ( .A1(n3844), .A2(n895), .B1(n896), .B2(n128), .ZN(n3189) );
  OAI22_X1 U1612 ( .A1(n3843), .A2(n894), .B1(n896), .B2(n127), .ZN(n3190) );
  OAI22_X1 U1613 ( .A1(n3842), .A2(n895), .B1(n896), .B2(n126), .ZN(n3191) );
  OAI22_X1 U1614 ( .A1(n3841), .A2(n894), .B1(n896), .B2(n125), .ZN(n3192) );
  OAI22_X1 U1615 ( .A1(n3840), .A2(n895), .B1(n896), .B2(n124), .ZN(n3193) );
  OAI22_X1 U1616 ( .A1(n3839), .A2(n894), .B1(n897), .B2(n123), .ZN(n3194) );
  OAI22_X1 U1617 ( .A1(n3838), .A2(n895), .B1(n897), .B2(n122), .ZN(n3195) );
  OAI22_X1 U1618 ( .A1(n3837), .A2(n894), .B1(n897), .B2(n121), .ZN(n3196) );
  OAI22_X1 U1619 ( .A1(n3836), .A2(n895), .B1(n897), .B2(n120), .ZN(n3197) );
  OAI22_X1 U1620 ( .A1(n3835), .A2(n895), .B1(n897), .B2(n119), .ZN(n3198) );
  OAI22_X1 U1621 ( .A1(n3834), .A2(n895), .B1(n898), .B2(n118), .ZN(n3199) );
  OAI22_X1 U1622 ( .A1(n3833), .A2(n895), .B1(n898), .B2(n117), .ZN(n3200) );
  OAI22_X1 U1623 ( .A1(n3832), .A2(n895), .B1(n898), .B2(n116), .ZN(n3201) );
  OAI22_X1 U1624 ( .A1(n3831), .A2(n895), .B1(n898), .B2(n115), .ZN(n3202) );
  OAI22_X1 U1625 ( .A1(n3830), .A2(n895), .B1(n898), .B2(n114), .ZN(n3203) );
  OAI22_X1 U1626 ( .A1(n3829), .A2(n895), .B1(n899), .B2(n113), .ZN(n3204) );
  OAI22_X1 U1627 ( .A1(n3828), .A2(n895), .B1(n899), .B2(n112), .ZN(n3205) );
  OAI22_X1 U1628 ( .A1(n3827), .A2(n895), .B1(n899), .B2(n111), .ZN(n3206) );
  OAI22_X1 U1629 ( .A1(n3826), .A2(n895), .B1(n899), .B2(n110), .ZN(n3207) );
  OAI22_X1 U1630 ( .A1(n3825), .A2(n895), .B1(n899), .B2(n109), .ZN(n3208) );
  OAI22_X1 U1631 ( .A1(n3824), .A2(n894), .B1(n900), .B2(n108), .ZN(n3209) );
  OAI22_X1 U1632 ( .A1(n3823), .A2(n894), .B1(n900), .B2(n107), .ZN(n3210) );
  OAI22_X1 U1633 ( .A1(n3822), .A2(n894), .B1(n900), .B2(n106), .ZN(n3211) );
  OAI22_X1 U1634 ( .A1(n3844), .A2(n886), .B1(n887), .B2(n96), .ZN(n3221) );
  OAI22_X1 U1635 ( .A1(n3843), .A2(n885), .B1(n887), .B2(n95), .ZN(n3222) );
  OAI22_X1 U1636 ( .A1(n3842), .A2(n886), .B1(n887), .B2(n94), .ZN(n3223) );
  OAI22_X1 U1637 ( .A1(n3841), .A2(n885), .B1(n887), .B2(n93), .ZN(n3224) );
  OAI22_X1 U1638 ( .A1(n3840), .A2(n886), .B1(n887), .B2(n92), .ZN(n3225) );
  OAI22_X1 U1639 ( .A1(n3839), .A2(n885), .B1(n888), .B2(n91), .ZN(n3226) );
  OAI22_X1 U1640 ( .A1(n3838), .A2(n886), .B1(n888), .B2(n90), .ZN(n3227) );
  OAI22_X1 U1641 ( .A1(n3837), .A2(n885), .B1(n888), .B2(n89), .ZN(n3228) );
  OAI22_X1 U1642 ( .A1(n3836), .A2(n886), .B1(n888), .B2(n88), .ZN(n3229) );
  OAI22_X1 U1643 ( .A1(n3835), .A2(n886), .B1(n888), .B2(n87), .ZN(n3230) );
  OAI22_X1 U1644 ( .A1(n3834), .A2(n886), .B1(n889), .B2(n86), .ZN(n3231) );
  OAI22_X1 U1645 ( .A1(n3833), .A2(n886), .B1(n889), .B2(n85), .ZN(n3232) );
  OAI22_X1 U1646 ( .A1(n3832), .A2(n886), .B1(n889), .B2(n84), .ZN(n3233) );
  OAI22_X1 U1647 ( .A1(n3831), .A2(n886), .B1(n889), .B2(n83), .ZN(n3234) );
  OAI22_X1 U1648 ( .A1(n3830), .A2(n886), .B1(n889), .B2(n82), .ZN(n3235) );
  OAI22_X1 U1649 ( .A1(n3829), .A2(n886), .B1(n890), .B2(n81), .ZN(n3236) );
  OAI22_X1 U1650 ( .A1(n3828), .A2(n886), .B1(n890), .B2(n80), .ZN(n3237) );
  OAI22_X1 U1651 ( .A1(n3827), .A2(n886), .B1(n890), .B2(n79), .ZN(n3238) );
  OAI22_X1 U1652 ( .A1(n3826), .A2(n886), .B1(n890), .B2(n78), .ZN(n3239) );
  OAI22_X1 U1653 ( .A1(n3825), .A2(n886), .B1(n890), .B2(n77), .ZN(n3240) );
  OAI22_X1 U1654 ( .A1(n3824), .A2(n885), .B1(n891), .B2(n76), .ZN(n3241) );
  OAI22_X1 U1655 ( .A1(n3823), .A2(n885), .B1(n891), .B2(n75), .ZN(n3242) );
  OAI22_X1 U1656 ( .A1(n3822), .A2(n885), .B1(n891), .B2(n74), .ZN(n3243) );
  OAI22_X1 U1657 ( .A1(n3844), .A2(n877), .B1(n878), .B2(n64), .ZN(n3253) );
  OAI22_X1 U1658 ( .A1(n3843), .A2(n876), .B1(n878), .B2(n63), .ZN(n3254) );
  OAI22_X1 U1659 ( .A1(n3842), .A2(n877), .B1(n878), .B2(n62), .ZN(n3255) );
  OAI22_X1 U1660 ( .A1(n3841), .A2(n876), .B1(n878), .B2(n61), .ZN(n3256) );
  OAI22_X1 U1661 ( .A1(n3840), .A2(n877), .B1(n878), .B2(n60), .ZN(n3257) );
  OAI22_X1 U1662 ( .A1(n3839), .A2(n876), .B1(n879), .B2(n59), .ZN(n3258) );
  OAI22_X1 U1663 ( .A1(n3838), .A2(n877), .B1(n879), .B2(n58), .ZN(n3259) );
  OAI22_X1 U1664 ( .A1(n3837), .A2(n876), .B1(n879), .B2(n57), .ZN(n3260) );
  OAI22_X1 U1665 ( .A1(n3836), .A2(n877), .B1(n879), .B2(n56), .ZN(n3261) );
  OAI22_X1 U1666 ( .A1(n3835), .A2(n877), .B1(n879), .B2(n55), .ZN(n3262) );
  OAI22_X1 U1667 ( .A1(n3834), .A2(n877), .B1(n880), .B2(n54), .ZN(n3263) );
  OAI22_X1 U1668 ( .A1(n3833), .A2(n877), .B1(n880), .B2(n53), .ZN(n3264) );
  OAI22_X1 U1669 ( .A1(n3832), .A2(n877), .B1(n880), .B2(n52), .ZN(n3265) );
  OAI22_X1 U1670 ( .A1(n3831), .A2(n877), .B1(n880), .B2(n51), .ZN(n3266) );
  OAI22_X1 U1671 ( .A1(n3830), .A2(n877), .B1(n880), .B2(n50), .ZN(n3267) );
  OAI22_X1 U1672 ( .A1(n3829), .A2(n877), .B1(n881), .B2(n49), .ZN(n3268) );
  OAI22_X1 U1673 ( .A1(n3828), .A2(n877), .B1(n881), .B2(n48), .ZN(n3269) );
  OAI22_X1 U1674 ( .A1(n3827), .A2(n877), .B1(n881), .B2(n47), .ZN(n3270) );
  OAI22_X1 U1675 ( .A1(n3826), .A2(n877), .B1(n881), .B2(n46), .ZN(n3271) );
  OAI22_X1 U1676 ( .A1(n3825), .A2(n877), .B1(n881), .B2(n45), .ZN(n3272) );
  OAI22_X1 U1677 ( .A1(n3824), .A2(n876), .B1(n882), .B2(n44), .ZN(n3273) );
  OAI22_X1 U1678 ( .A1(n3823), .A2(n876), .B1(n882), .B2(n43), .ZN(n3274) );
  OAI22_X1 U1679 ( .A1(n3822), .A2(n876), .B1(n882), .B2(n42), .ZN(n3275) );
  OAI22_X1 U1680 ( .A1(n3821), .A2(n794), .B1(n800), .B2(n969), .ZN(n2796) );
  OAI22_X1 U1681 ( .A1(n3820), .A2(n794), .B1(n800), .B2(n968), .ZN(n2797) );
  OAI22_X1 U1682 ( .A1(n3819), .A2(n794), .B1(n865), .B2(n967), .ZN(n2798) );
  OAI22_X1 U1683 ( .A1(n3818), .A2(n794), .B1(n865), .B2(n966), .ZN(n2799) );
  OAI22_X1 U1684 ( .A1(n3817), .A2(n794), .B1(n865), .B2(n965), .ZN(n2800) );
  OAI22_X1 U1685 ( .A1(n3816), .A2(n794), .B1(n865), .B2(n964), .ZN(n2801) );
  OAI22_X1 U1686 ( .A1(n3815), .A2(n794), .B1(n865), .B2(n963), .ZN(n2802) );
  OAI22_X1 U1687 ( .A1(n3814), .A2(n794), .B1(n866), .B2(n962), .ZN(n2803) );
  OAI22_X1 U1688 ( .A1(n3813), .A2(n794), .B1(n866), .B2(n961), .ZN(n2804) );
  OAI22_X1 U1689 ( .A1(n3821), .A2(n785), .B1(n791), .B2(n937), .ZN(n2828) );
  OAI22_X1 U1690 ( .A1(n3820), .A2(n785), .B1(n791), .B2(n936), .ZN(n2829) );
  OAI22_X1 U1691 ( .A1(n3819), .A2(n785), .B1(n792), .B2(n935), .ZN(n2830) );
  OAI22_X1 U1692 ( .A1(n3818), .A2(n785), .B1(n792), .B2(n934), .ZN(n2831) );
  OAI22_X1 U1693 ( .A1(n3817), .A2(n785), .B1(n792), .B2(n933), .ZN(n2832) );
  OAI22_X1 U1694 ( .A1(n3816), .A2(n785), .B1(n792), .B2(n932), .ZN(n2833) );
  OAI22_X1 U1695 ( .A1(n3815), .A2(n785), .B1(n792), .B2(n931), .ZN(n2834) );
  OAI22_X1 U1696 ( .A1(n3814), .A2(n785), .B1(n793), .B2(n930), .ZN(n2835) );
  OAI22_X1 U1697 ( .A1(n3813), .A2(n785), .B1(n793), .B2(n929), .ZN(n2836) );
  OAI22_X1 U1698 ( .A1(n3821), .A2(n758), .B1(n764), .B2(n841), .ZN(n2860) );
  OAI22_X1 U1699 ( .A1(n3820), .A2(n758), .B1(n764), .B2(n840), .ZN(n2861) );
  OAI22_X1 U1700 ( .A1(n3819), .A2(n758), .B1(n765), .B2(n839), .ZN(n2862) );
  OAI22_X1 U1701 ( .A1(n3818), .A2(n758), .B1(n765), .B2(n838), .ZN(n2863) );
  OAI22_X1 U1702 ( .A1(n3817), .A2(n758), .B1(n765), .B2(n837), .ZN(n2864) );
  OAI22_X1 U1703 ( .A1(n3816), .A2(n758), .B1(n765), .B2(n836), .ZN(n2865) );
  OAI22_X1 U1704 ( .A1(n3815), .A2(n758), .B1(n765), .B2(n835), .ZN(n2866) );
  OAI22_X1 U1705 ( .A1(n3814), .A2(n758), .B1(n766), .B2(n834), .ZN(n2867) );
  OAI22_X1 U1706 ( .A1(n3813), .A2(n758), .B1(n766), .B2(n833), .ZN(n2868) );
  OAI22_X1 U1707 ( .A1(n3821), .A2(n749), .B1(n755), .B2(n809), .ZN(n2892) );
  OAI22_X1 U1708 ( .A1(n3820), .A2(n749), .B1(n755), .B2(n808), .ZN(n2893) );
  OAI22_X1 U1709 ( .A1(n3819), .A2(n749), .B1(n756), .B2(n807), .ZN(n2894) );
  OAI22_X1 U1710 ( .A1(n3818), .A2(n749), .B1(n756), .B2(n806), .ZN(n2895) );
  OAI22_X1 U1711 ( .A1(n3817), .A2(n749), .B1(n756), .B2(n805), .ZN(n2896) );
  OAI22_X1 U1712 ( .A1(n3816), .A2(n749), .B1(n756), .B2(n804), .ZN(n2897) );
  OAI22_X1 U1713 ( .A1(n3815), .A2(n749), .B1(n756), .B2(n803), .ZN(n2898) );
  OAI22_X1 U1714 ( .A1(n3814), .A2(n749), .B1(n757), .B2(n802), .ZN(n2899) );
  OAI22_X1 U1715 ( .A1(n3813), .A2(n749), .B1(n757), .B2(n801), .ZN(n2900) );
  OAI22_X1 U1716 ( .A1(n3821), .A2(n704), .B1(n710), .B2(n649), .ZN(n2924) );
  OAI22_X1 U1717 ( .A1(n3820), .A2(n704), .B1(n710), .B2(n648), .ZN(n2925) );
  OAI22_X1 U1718 ( .A1(n3819), .A2(n704), .B1(n711), .B2(n647), .ZN(n2926) );
  OAI22_X1 U1719 ( .A1(n3818), .A2(n704), .B1(n711), .B2(n646), .ZN(n2927) );
  OAI22_X1 U1720 ( .A1(n3817), .A2(n704), .B1(n711), .B2(n645), .ZN(n2928) );
  OAI22_X1 U1721 ( .A1(n3816), .A2(n704), .B1(n711), .B2(n644), .ZN(n2929) );
  OAI22_X1 U1722 ( .A1(n3815), .A2(n704), .B1(n711), .B2(n643), .ZN(n2930) );
  OAI22_X1 U1723 ( .A1(n3814), .A2(n704), .B1(n712), .B2(n642), .ZN(n2931) );
  OAI22_X1 U1724 ( .A1(n3813), .A2(n704), .B1(n712), .B2(n641), .ZN(n2932) );
  OAI22_X1 U1725 ( .A1(n3821), .A2(n695), .B1(n701), .B2(n617), .ZN(n2956) );
  OAI22_X1 U1726 ( .A1(n3820), .A2(n695), .B1(n701), .B2(n616), .ZN(n2957) );
  OAI22_X1 U1727 ( .A1(n3819), .A2(n695), .B1(n702), .B2(n615), .ZN(n2958) );
  OAI22_X1 U1728 ( .A1(n3818), .A2(n695), .B1(n702), .B2(n614), .ZN(n2959) );
  OAI22_X1 U1729 ( .A1(n3817), .A2(n695), .B1(n702), .B2(n613), .ZN(n2960) );
  OAI22_X1 U1730 ( .A1(n3816), .A2(n695), .B1(n702), .B2(n612), .ZN(n2961) );
  OAI22_X1 U1731 ( .A1(n3815), .A2(n695), .B1(n702), .B2(n611), .ZN(n2962) );
  OAI22_X1 U1732 ( .A1(n3814), .A2(n695), .B1(n703), .B2(n610), .ZN(n2963) );
  OAI22_X1 U1733 ( .A1(n3813), .A2(n695), .B1(n703), .B2(n609), .ZN(n2964) );
  OAI22_X1 U1734 ( .A1(n3821), .A2(n604), .B1(n674), .B2(n521), .ZN(n2988) );
  OAI22_X1 U1735 ( .A1(n3820), .A2(n604), .B1(n674), .B2(n520), .ZN(n2989) );
  OAI22_X1 U1736 ( .A1(n3819), .A2(n604), .B1(n675), .B2(n519), .ZN(n2990) );
  OAI22_X1 U1737 ( .A1(n3818), .A2(n604), .B1(n675), .B2(n518), .ZN(n2991) );
  OAI22_X1 U1738 ( .A1(n3817), .A2(n604), .B1(n675), .B2(n517), .ZN(n2992) );
  OAI22_X1 U1739 ( .A1(n3816), .A2(n604), .B1(n675), .B2(n516), .ZN(n2993) );
  OAI22_X1 U1740 ( .A1(n3815), .A2(n604), .B1(n675), .B2(n515), .ZN(n2994) );
  OAI22_X1 U1741 ( .A1(n3814), .A2(n604), .B1(n676), .B2(n514), .ZN(n2995) );
  OAI22_X1 U1742 ( .A1(n3813), .A2(n604), .B1(n676), .B2(n513), .ZN(n2996) );
  OAI22_X1 U1743 ( .A1(n3821), .A2(n595), .B1(n601), .B2(n489), .ZN(n3020) );
  OAI22_X1 U1744 ( .A1(n3820), .A2(n595), .B1(n601), .B2(n488), .ZN(n3021) );
  OAI22_X1 U1745 ( .A1(n3819), .A2(n595), .B1(n602), .B2(n487), .ZN(n3022) );
  OAI22_X1 U1746 ( .A1(n3818), .A2(n595), .B1(n602), .B2(n486), .ZN(n3023) );
  OAI22_X1 U1747 ( .A1(n3817), .A2(n595), .B1(n602), .B2(n485), .ZN(n3024) );
  OAI22_X1 U1748 ( .A1(n3816), .A2(n595), .B1(n602), .B2(n484), .ZN(n3025) );
  OAI22_X1 U1749 ( .A1(n3815), .A2(n595), .B1(n602), .B2(n483), .ZN(n3026) );
  OAI22_X1 U1750 ( .A1(n3814), .A2(n595), .B1(n603), .B2(n482), .ZN(n3027) );
  OAI22_X1 U1751 ( .A1(n3813), .A2(n595), .B1(n603), .B2(n481), .ZN(n3028) );
  OAI22_X1 U1752 ( .A1(n3821), .A2(n586), .B1(n592), .B2(n457), .ZN(n3052) );
  OAI22_X1 U1753 ( .A1(n3820), .A2(n586), .B1(n592), .B2(n456), .ZN(n3053) );
  OAI22_X1 U1754 ( .A1(n3819), .A2(n586), .B1(n593), .B2(n455), .ZN(n3054) );
  OAI22_X1 U1755 ( .A1(n3818), .A2(n586), .B1(n593), .B2(n454), .ZN(n3055) );
  OAI22_X1 U1756 ( .A1(n3817), .A2(n586), .B1(n593), .B2(n453), .ZN(n3056) );
  OAI22_X1 U1757 ( .A1(n3816), .A2(n586), .B1(n593), .B2(n452), .ZN(n3057) );
  OAI22_X1 U1758 ( .A1(n3815), .A2(n586), .B1(n593), .B2(n451), .ZN(n3058) );
  OAI22_X1 U1759 ( .A1(n3814), .A2(n586), .B1(n594), .B2(n450), .ZN(n3059) );
  OAI22_X1 U1760 ( .A1(n3813), .A2(n586), .B1(n594), .B2(n449), .ZN(n3060) );
  OAI22_X1 U1761 ( .A1(n3821), .A2(n577), .B1(n583), .B2(n425), .ZN(n3084) );
  OAI22_X1 U1762 ( .A1(n3820), .A2(n577), .B1(n583), .B2(n424), .ZN(n3085) );
  OAI22_X1 U1763 ( .A1(n3819), .A2(n577), .B1(n584), .B2(n423), .ZN(n3086) );
  OAI22_X1 U1764 ( .A1(n3818), .A2(n577), .B1(n584), .B2(n422), .ZN(n3087) );
  OAI22_X1 U1765 ( .A1(n3817), .A2(n577), .B1(n584), .B2(n421), .ZN(n3088) );
  OAI22_X1 U1766 ( .A1(n3816), .A2(n577), .B1(n584), .B2(n420), .ZN(n3089) );
  OAI22_X1 U1767 ( .A1(n3815), .A2(n577), .B1(n584), .B2(n419), .ZN(n3090) );
  OAI22_X1 U1768 ( .A1(n3814), .A2(n577), .B1(n585), .B2(n418), .ZN(n3091) );
  OAI22_X1 U1769 ( .A1(n3813), .A2(n577), .B1(n585), .B2(n417), .ZN(n3092) );
  OAI22_X1 U1770 ( .A1(n3821), .A2(n550), .B1(n556), .B2(n329), .ZN(n3116) );
  OAI22_X1 U1771 ( .A1(n3820), .A2(n550), .B1(n556), .B2(n328), .ZN(n3117) );
  OAI22_X1 U1772 ( .A1(n3819), .A2(n550), .B1(n557), .B2(n327), .ZN(n3118) );
  OAI22_X1 U1773 ( .A1(n3818), .A2(n550), .B1(n557), .B2(n326), .ZN(n3119) );
  OAI22_X1 U1774 ( .A1(n3817), .A2(n550), .B1(n557), .B2(n325), .ZN(n3120) );
  OAI22_X1 U1775 ( .A1(n3816), .A2(n550), .B1(n557), .B2(n324), .ZN(n3121) );
  OAI22_X1 U1776 ( .A1(n3815), .A2(n550), .B1(n557), .B2(n323), .ZN(n3122) );
  OAI22_X1 U1777 ( .A1(n3814), .A2(n550), .B1(n558), .B2(n322), .ZN(n3123) );
  OAI22_X1 U1778 ( .A1(n3813), .A2(n550), .B1(n558), .B2(n321), .ZN(n3124) );
  OAI22_X1 U1779 ( .A1(n3821), .A2(n413), .B1(n547), .B2(n297), .ZN(n3148) );
  OAI22_X1 U1780 ( .A1(n3820), .A2(n413), .B1(n547), .B2(n296), .ZN(n3149) );
  OAI22_X1 U1781 ( .A1(n3819), .A2(n413), .B1(n548), .B2(n295), .ZN(n3150) );
  OAI22_X1 U1782 ( .A1(n3818), .A2(n413), .B1(n548), .B2(n294), .ZN(n3151) );
  OAI22_X1 U1783 ( .A1(n3817), .A2(n413), .B1(n548), .B2(n293), .ZN(n3152) );
  OAI22_X1 U1784 ( .A1(n3816), .A2(n413), .B1(n548), .B2(n292), .ZN(n3153) );
  OAI22_X1 U1785 ( .A1(n3815), .A2(n413), .B1(n548), .B2(n291), .ZN(n3154) );
  OAI22_X1 U1786 ( .A1(n3814), .A2(n413), .B1(n549), .B2(n290), .ZN(n3155) );
  OAI22_X1 U1787 ( .A1(n3813), .A2(n413), .B1(n549), .B2(n289), .ZN(n3156) );
  OAI22_X1 U1788 ( .A1(n3821), .A2(n903), .B1(n909), .B2(n137), .ZN(n3180) );
  OAI22_X1 U1789 ( .A1(n3820), .A2(n903), .B1(n909), .B2(n136), .ZN(n3181) );
  OAI22_X1 U1790 ( .A1(n3819), .A2(n903), .B1(n910), .B2(n135), .ZN(n3182) );
  OAI22_X1 U1791 ( .A1(n3818), .A2(n903), .B1(n910), .B2(n134), .ZN(n3183) );
  OAI22_X1 U1792 ( .A1(n3817), .A2(n903), .B1(n910), .B2(n133), .ZN(n3184) );
  OAI22_X1 U1793 ( .A1(n3816), .A2(n903), .B1(n910), .B2(n132), .ZN(n3185) );
  OAI22_X1 U1794 ( .A1(n3815), .A2(n903), .B1(n910), .B2(n131), .ZN(n3186) );
  OAI22_X1 U1795 ( .A1(n3814), .A2(n903), .B1(n911), .B2(n130), .ZN(n3187) );
  OAI22_X1 U1796 ( .A1(n3813), .A2(n903), .B1(n911), .B2(n129), .ZN(n3188) );
  OAI22_X1 U1797 ( .A1(n3821), .A2(n894), .B1(n900), .B2(n105), .ZN(n3212) );
  OAI22_X1 U1798 ( .A1(n3820), .A2(n894), .B1(n900), .B2(n104), .ZN(n3213) );
  OAI22_X1 U1799 ( .A1(n3819), .A2(n894), .B1(n901), .B2(n103), .ZN(n3214) );
  OAI22_X1 U1800 ( .A1(n3818), .A2(n894), .B1(n901), .B2(n102), .ZN(n3215) );
  OAI22_X1 U1801 ( .A1(n3817), .A2(n894), .B1(n901), .B2(n101), .ZN(n3216) );
  OAI22_X1 U1802 ( .A1(n3816), .A2(n894), .B1(n901), .B2(n100), .ZN(n3217) );
  OAI22_X1 U1803 ( .A1(n3815), .A2(n894), .B1(n901), .B2(n99), .ZN(n3218) );
  OAI22_X1 U1804 ( .A1(n3814), .A2(n894), .B1(n902), .B2(n98), .ZN(n3219) );
  OAI22_X1 U1805 ( .A1(n3813), .A2(n894), .B1(n902), .B2(n97), .ZN(n3220) );
  OAI22_X1 U1806 ( .A1(n3821), .A2(n885), .B1(n891), .B2(n73), .ZN(n3244) );
  OAI22_X1 U1807 ( .A1(n3820), .A2(n885), .B1(n891), .B2(n72), .ZN(n3245) );
  OAI22_X1 U1808 ( .A1(n3819), .A2(n885), .B1(n892), .B2(n71), .ZN(n3246) );
  OAI22_X1 U1809 ( .A1(n3818), .A2(n885), .B1(n892), .B2(n70), .ZN(n3247) );
  OAI22_X1 U1810 ( .A1(n3817), .A2(n885), .B1(n892), .B2(n69), .ZN(n3248) );
  OAI22_X1 U1811 ( .A1(n3816), .A2(n885), .B1(n892), .B2(n68), .ZN(n3249) );
  OAI22_X1 U1812 ( .A1(n3815), .A2(n885), .B1(n892), .B2(n67), .ZN(n3250) );
  OAI22_X1 U1813 ( .A1(n3814), .A2(n885), .B1(n893), .B2(n66), .ZN(n3251) );
  OAI22_X1 U1814 ( .A1(n3813), .A2(n885), .B1(n893), .B2(n65), .ZN(n3252) );
  OAI22_X1 U1815 ( .A1(n3821), .A2(n876), .B1(n882), .B2(n41), .ZN(n3276) );
  OAI22_X1 U1816 ( .A1(n3820), .A2(n876), .B1(n882), .B2(n40), .ZN(n3277) );
  OAI22_X1 U1817 ( .A1(n3819), .A2(n876), .B1(n883), .B2(n39), .ZN(n3278) );
  OAI22_X1 U1818 ( .A1(n3818), .A2(n876), .B1(n883), .B2(n38), .ZN(n3279) );
  OAI22_X1 U1819 ( .A1(n3817), .A2(n876), .B1(n883), .B2(n37), .ZN(n3280) );
  OAI22_X1 U1820 ( .A1(n3816), .A2(n876), .B1(n883), .B2(n36), .ZN(n3281) );
  OAI22_X1 U1821 ( .A1(n3815), .A2(n876), .B1(n883), .B2(n35), .ZN(n3282) );
  OAI22_X1 U1822 ( .A1(n3814), .A2(n876), .B1(n884), .B2(n34), .ZN(n3283) );
  OAI22_X1 U1823 ( .A1(n3813), .A2(n876), .B1(n884), .B2(n33), .ZN(n3284) );
  AOI22_X1 U1824 ( .A1(n374), .A2(\registers[23][0] ), .B1(n371), .B2(
        \registers[22][0] ), .ZN(n2162) );
  AOI22_X1 U1825 ( .A1(n362), .A2(\registers[25][0] ), .B1(n359), .B2(
        \registers[24][0] ), .ZN(n2166) );
  AOI22_X1 U1826 ( .A1(n286), .A2(\registers[29][0] ), .B1(n283), .B2(
        \registers[28][0] ), .ZN(n2169) );
  AOI22_X1 U1827 ( .A1(n374), .A2(\registers[23][1] ), .B1(n371), .B2(
        \registers[22][1] ), .ZN(n2141) );
  AOI22_X1 U1828 ( .A1(n362), .A2(\registers[25][1] ), .B1(n359), .B2(
        \registers[24][1] ), .ZN(n2142) );
  AOI22_X1 U1829 ( .A1(n286), .A2(\registers[29][1] ), .B1(n283), .B2(
        \registers[28][1] ), .ZN(n2143) );
  AOI22_X1 U1830 ( .A1(n374), .A2(\registers[23][2] ), .B1(n371), .B2(
        \registers[22][2] ), .ZN(n2124) );
  AOI22_X1 U1831 ( .A1(n362), .A2(\registers[25][2] ), .B1(n359), .B2(
        \registers[24][2] ), .ZN(n2125) );
  AOI22_X1 U1832 ( .A1(n286), .A2(\registers[29][2] ), .B1(n283), .B2(
        \registers[28][2] ), .ZN(n2126) );
  AOI22_X1 U1833 ( .A1(n374), .A2(\registers[23][3] ), .B1(n371), .B2(
        \registers[22][3] ), .ZN(n2107) );
  AOI22_X1 U1834 ( .A1(n362), .A2(\registers[25][3] ), .B1(n359), .B2(
        \registers[24][3] ), .ZN(n2108) );
  AOI22_X1 U1835 ( .A1(n286), .A2(\registers[29][3] ), .B1(n283), .B2(
        \registers[28][3] ), .ZN(n2109) );
  AOI22_X1 U1836 ( .A1(n374), .A2(\registers[23][4] ), .B1(n371), .B2(
        \registers[22][4] ), .ZN(n2090) );
  AOI22_X1 U1837 ( .A1(n362), .A2(\registers[25][4] ), .B1(n359), .B2(
        \registers[24][4] ), .ZN(n2091) );
  AOI22_X1 U1838 ( .A1(n286), .A2(\registers[29][4] ), .B1(n283), .B2(
        \registers[28][4] ), .ZN(n2092) );
  AOI22_X1 U1839 ( .A1(n374), .A2(\registers[23][5] ), .B1(n371), .B2(
        \registers[22][5] ), .ZN(n2073) );
  AOI22_X1 U1840 ( .A1(n362), .A2(\registers[25][5] ), .B1(n359), .B2(
        \registers[24][5] ), .ZN(n2074) );
  AOI22_X1 U1841 ( .A1(n286), .A2(\registers[29][5] ), .B1(n283), .B2(
        \registers[28][5] ), .ZN(n2075) );
  AOI22_X1 U1842 ( .A1(n374), .A2(\registers[23][6] ), .B1(n371), .B2(
        \registers[22][6] ), .ZN(n2056) );
  AOI22_X1 U1843 ( .A1(n362), .A2(\registers[25][6] ), .B1(n359), .B2(
        \registers[24][6] ), .ZN(n2057) );
  AOI22_X1 U1844 ( .A1(n286), .A2(\registers[29][6] ), .B1(n283), .B2(
        \registers[28][6] ), .ZN(n2058) );
  AOI22_X1 U1845 ( .A1(n374), .A2(\registers[23][7] ), .B1(n371), .B2(
        \registers[22][7] ), .ZN(n2039) );
  AOI22_X1 U1846 ( .A1(n362), .A2(\registers[25][7] ), .B1(n359), .B2(
        \registers[24][7] ), .ZN(n2040) );
  AOI22_X1 U1847 ( .A1(n286), .A2(\registers[29][7] ), .B1(n283), .B2(
        \registers[28][7] ), .ZN(n2041) );
  AOI22_X1 U1848 ( .A1(n374), .A2(\registers[23][8] ), .B1(n371), .B2(
        \registers[22][8] ), .ZN(n2022) );
  AOI22_X1 U1849 ( .A1(n362), .A2(\registers[25][8] ), .B1(n359), .B2(
        \registers[24][8] ), .ZN(n2023) );
  AOI22_X1 U1850 ( .A1(n286), .A2(\registers[29][8] ), .B1(n283), .B2(
        \registers[28][8] ), .ZN(n2024) );
  AOI22_X1 U1851 ( .A1(n374), .A2(\registers[23][9] ), .B1(n371), .B2(
        \registers[22][9] ), .ZN(n2005) );
  AOI22_X1 U1852 ( .A1(n362), .A2(\registers[25][9] ), .B1(n359), .B2(
        \registers[24][9] ), .ZN(n2006) );
  AOI22_X1 U1853 ( .A1(n286), .A2(\registers[29][9] ), .B1(n283), .B2(
        \registers[28][9] ), .ZN(n2007) );
  AOI22_X1 U1854 ( .A1(n374), .A2(\registers[23][10] ), .B1(n371), .B2(
        \registers[22][10] ), .ZN(n1988) );
  AOI22_X1 U1855 ( .A1(n362), .A2(\registers[25][10] ), .B1(n359), .B2(
        \registers[24][10] ), .ZN(n1989) );
  AOI22_X1 U1856 ( .A1(n286), .A2(\registers[29][10] ), .B1(n283), .B2(
        \registers[28][10] ), .ZN(n1990) );
  AOI22_X1 U1857 ( .A1(n375), .A2(\registers[23][11] ), .B1(n372), .B2(
        \registers[22][11] ), .ZN(n1971) );
  AOI22_X1 U1858 ( .A1(n363), .A2(\registers[25][11] ), .B1(n360), .B2(
        \registers[24][11] ), .ZN(n1972) );
  AOI22_X1 U1859 ( .A1(n287), .A2(\registers[29][11] ), .B1(n284), .B2(
        \registers[28][11] ), .ZN(n1973) );
  AOI22_X1 U1860 ( .A1(n375), .A2(\registers[23][12] ), .B1(n372), .B2(
        \registers[22][12] ), .ZN(n1954) );
  AOI22_X1 U1861 ( .A1(n363), .A2(\registers[25][12] ), .B1(n360), .B2(
        \registers[24][12] ), .ZN(n1955) );
  AOI22_X1 U1862 ( .A1(n287), .A2(\registers[29][12] ), .B1(n284), .B2(
        \registers[28][12] ), .ZN(n1956) );
  AOI22_X1 U1863 ( .A1(n375), .A2(\registers[23][13] ), .B1(n372), .B2(
        \registers[22][13] ), .ZN(n1937) );
  AOI22_X1 U1864 ( .A1(n363), .A2(\registers[25][13] ), .B1(n360), .B2(
        \registers[24][13] ), .ZN(n1938) );
  AOI22_X1 U1865 ( .A1(n287), .A2(\registers[29][13] ), .B1(n284), .B2(
        \registers[28][13] ), .ZN(n1939) );
  AOI22_X1 U1866 ( .A1(n375), .A2(\registers[23][14] ), .B1(n372), .B2(
        \registers[22][14] ), .ZN(n1920) );
  AOI22_X1 U1867 ( .A1(n363), .A2(\registers[25][14] ), .B1(n360), .B2(
        \registers[24][14] ), .ZN(n1921) );
  AOI22_X1 U1868 ( .A1(n287), .A2(\registers[29][14] ), .B1(n284), .B2(
        \registers[28][14] ), .ZN(n1922) );
  AOI22_X1 U1869 ( .A1(n375), .A2(\registers[23][15] ), .B1(n372), .B2(
        \registers[22][15] ), .ZN(n1903) );
  AOI22_X1 U1870 ( .A1(n363), .A2(\registers[25][15] ), .B1(n360), .B2(
        \registers[24][15] ), .ZN(n1904) );
  AOI22_X1 U1871 ( .A1(n287), .A2(\registers[29][15] ), .B1(n284), .B2(
        \registers[28][15] ), .ZN(n1905) );
  AOI22_X1 U1872 ( .A1(n375), .A2(\registers[23][16] ), .B1(n372), .B2(
        \registers[22][16] ), .ZN(n1886) );
  AOI22_X1 U1873 ( .A1(n363), .A2(\registers[25][16] ), .B1(n360), .B2(
        \registers[24][16] ), .ZN(n1887) );
  AOI22_X1 U1874 ( .A1(n287), .A2(\registers[29][16] ), .B1(n284), .B2(
        \registers[28][16] ), .ZN(n1888) );
  AOI22_X1 U1875 ( .A1(n375), .A2(\registers[23][17] ), .B1(n372), .B2(
        \registers[22][17] ), .ZN(n1869) );
  AOI22_X1 U1876 ( .A1(n363), .A2(\registers[25][17] ), .B1(n360), .B2(
        \registers[24][17] ), .ZN(n1870) );
  AOI22_X1 U1877 ( .A1(n287), .A2(\registers[29][17] ), .B1(n284), .B2(
        \registers[28][17] ), .ZN(n1871) );
  AOI22_X1 U1878 ( .A1(n375), .A2(\registers[23][18] ), .B1(n372), .B2(
        \registers[22][18] ), .ZN(n1852) );
  AOI22_X1 U1879 ( .A1(n363), .A2(\registers[25][18] ), .B1(n360), .B2(
        \registers[24][18] ), .ZN(n1853) );
  AOI22_X1 U1880 ( .A1(n287), .A2(\registers[29][18] ), .B1(n284), .B2(
        \registers[28][18] ), .ZN(n1854) );
  AOI22_X1 U1881 ( .A1(n375), .A2(\registers[23][19] ), .B1(n372), .B2(
        \registers[22][19] ), .ZN(n1835) );
  AOI22_X1 U1882 ( .A1(n363), .A2(\registers[25][19] ), .B1(n360), .B2(
        \registers[24][19] ), .ZN(n1836) );
  AOI22_X1 U1883 ( .A1(n287), .A2(\registers[29][19] ), .B1(n284), .B2(
        \registers[28][19] ), .ZN(n1837) );
  AOI22_X1 U1884 ( .A1(n375), .A2(\registers[23][20] ), .B1(n372), .B2(
        \registers[22][20] ), .ZN(n1818) );
  AOI22_X1 U1885 ( .A1(n363), .A2(\registers[25][20] ), .B1(n360), .B2(
        \registers[24][20] ), .ZN(n1819) );
  AOI22_X1 U1886 ( .A1(n287), .A2(\registers[29][20] ), .B1(n284), .B2(
        \registers[28][20] ), .ZN(n1820) );
  AOI22_X1 U1887 ( .A1(n375), .A2(\registers[23][21] ), .B1(n372), .B2(
        \registers[22][21] ), .ZN(n1801) );
  AOI22_X1 U1888 ( .A1(n363), .A2(\registers[25][21] ), .B1(n360), .B2(
        \registers[24][21] ), .ZN(n1802) );
  AOI22_X1 U1889 ( .A1(n287), .A2(\registers[29][21] ), .B1(n284), .B2(
        \registers[28][21] ), .ZN(n1803) );
  AOI22_X1 U1890 ( .A1(n376), .A2(\registers[23][22] ), .B1(n373), .B2(
        \registers[22][22] ), .ZN(n1784) );
  AOI22_X1 U1891 ( .A1(n364), .A2(\registers[25][22] ), .B1(n361), .B2(
        \registers[24][22] ), .ZN(n1785) );
  AOI22_X1 U1892 ( .A1(n288), .A2(\registers[29][22] ), .B1(n285), .B2(
        \registers[28][22] ), .ZN(n1786) );
  AOI22_X1 U1893 ( .A1(n376), .A2(\registers[23][23] ), .B1(n373), .B2(
        \registers[22][23] ), .ZN(n1767) );
  AOI22_X1 U1894 ( .A1(n364), .A2(\registers[25][23] ), .B1(n361), .B2(
        \registers[24][23] ), .ZN(n1768) );
  AOI22_X1 U1895 ( .A1(n288), .A2(\registers[29][23] ), .B1(n285), .B2(
        \registers[28][23] ), .ZN(n1769) );
  AOI22_X1 U1896 ( .A1(n376), .A2(\registers[23][24] ), .B1(n373), .B2(
        \registers[22][24] ), .ZN(n1750) );
  AOI22_X1 U1897 ( .A1(n364), .A2(\registers[25][24] ), .B1(n361), .B2(
        \registers[24][24] ), .ZN(n1751) );
  AOI22_X1 U1898 ( .A1(n288), .A2(\registers[29][24] ), .B1(n285), .B2(
        \registers[28][24] ), .ZN(n1752) );
  AOI22_X1 U1899 ( .A1(n376), .A2(\registers[23][25] ), .B1(n373), .B2(
        \registers[22][25] ), .ZN(n1733) );
  AOI22_X1 U1900 ( .A1(n364), .A2(\registers[25][25] ), .B1(n361), .B2(
        \registers[24][25] ), .ZN(n1734) );
  AOI22_X1 U1901 ( .A1(n288), .A2(\registers[29][25] ), .B1(n285), .B2(
        \registers[28][25] ), .ZN(n1735) );
  AOI22_X1 U1902 ( .A1(n376), .A2(\registers[23][26] ), .B1(n373), .B2(
        \registers[22][26] ), .ZN(n1716) );
  AOI22_X1 U1903 ( .A1(n364), .A2(\registers[25][26] ), .B1(n361), .B2(
        \registers[24][26] ), .ZN(n1717) );
  AOI22_X1 U1904 ( .A1(n288), .A2(\registers[29][26] ), .B1(n285), .B2(
        \registers[28][26] ), .ZN(n1718) );
  AOI22_X1 U1905 ( .A1(n376), .A2(\registers[23][27] ), .B1(n373), .B2(
        \registers[22][27] ), .ZN(n1699) );
  AOI22_X1 U1906 ( .A1(n364), .A2(\registers[25][27] ), .B1(n361), .B2(
        \registers[24][27] ), .ZN(n1700) );
  AOI22_X1 U1907 ( .A1(n288), .A2(\registers[29][27] ), .B1(n285), .B2(
        \registers[28][27] ), .ZN(n1701) );
  AOI22_X1 U1908 ( .A1(n376), .A2(\registers[23][28] ), .B1(n373), .B2(
        \registers[22][28] ), .ZN(n1682) );
  AOI22_X1 U1909 ( .A1(n364), .A2(\registers[25][28] ), .B1(n361), .B2(
        \registers[24][28] ), .ZN(n1683) );
  AOI22_X1 U1910 ( .A1(n288), .A2(\registers[29][28] ), .B1(n285), .B2(
        \registers[28][28] ), .ZN(n1684) );
  AOI22_X1 U1911 ( .A1(n376), .A2(\registers[23][29] ), .B1(n373), .B2(
        \registers[22][29] ), .ZN(n1665) );
  AOI22_X1 U1912 ( .A1(n364), .A2(\registers[25][29] ), .B1(n361), .B2(
        \registers[24][29] ), .ZN(n1666) );
  AOI22_X1 U1913 ( .A1(n288), .A2(\registers[29][29] ), .B1(n285), .B2(
        \registers[28][29] ), .ZN(n1667) );
  AOI22_X1 U1914 ( .A1(n376), .A2(\registers[23][30] ), .B1(n373), .B2(
        \registers[22][30] ), .ZN(n1648) );
  AOI22_X1 U1915 ( .A1(n364), .A2(\registers[25][30] ), .B1(n361), .B2(
        \registers[24][30] ), .ZN(n1649) );
  AOI22_X1 U1916 ( .A1(n288), .A2(\registers[29][30] ), .B1(n285), .B2(
        \registers[28][30] ), .ZN(n1650) );
  AOI22_X1 U1917 ( .A1(n376), .A2(\registers[23][31] ), .B1(n373), .B2(
        \registers[22][31] ), .ZN(n1606) );
  AOI22_X1 U1918 ( .A1(n364), .A2(\registers[25][31] ), .B1(n361), .B2(
        \registers[24][31] ), .ZN(n1611) );
  AOI22_X1 U1919 ( .A1(n288), .A2(\registers[29][31] ), .B1(n285), .B2(
        \registers[28][31] ), .ZN(n1616) );
  AOI22_X1 U1920 ( .A1(n217), .A2(\registers[23][0] ), .B1(n214), .B2(
        \registers[22][0] ), .ZN(n2753) );
  AOI22_X1 U1921 ( .A1(n205), .A2(\registers[25][0] ), .B1(n202), .B2(
        \registers[24][0] ), .ZN(n2757) );
  AOI22_X1 U1922 ( .A1(n193), .A2(\registers[29][0] ), .B1(n190), .B2(
        \registers[28][0] ), .ZN(n2760) );
  AOI22_X1 U1923 ( .A1(n217), .A2(\registers[23][1] ), .B1(n214), .B2(
        \registers[22][1] ), .ZN(n2732) );
  AOI22_X1 U1924 ( .A1(n205), .A2(\registers[25][1] ), .B1(n202), .B2(
        \registers[24][1] ), .ZN(n2733) );
  AOI22_X1 U1925 ( .A1(n193), .A2(\registers[29][1] ), .B1(n190), .B2(
        \registers[28][1] ), .ZN(n2734) );
  AOI22_X1 U1926 ( .A1(n217), .A2(\registers[23][2] ), .B1(n214), .B2(
        \registers[22][2] ), .ZN(n2715) );
  AOI22_X1 U1927 ( .A1(n205), .A2(\registers[25][2] ), .B1(n202), .B2(
        \registers[24][2] ), .ZN(n2716) );
  AOI22_X1 U1928 ( .A1(n193), .A2(\registers[29][2] ), .B1(n190), .B2(
        \registers[28][2] ), .ZN(n2717) );
  AOI22_X1 U1929 ( .A1(n217), .A2(\registers[23][3] ), .B1(n214), .B2(
        \registers[22][3] ), .ZN(n2698) );
  AOI22_X1 U1930 ( .A1(n205), .A2(\registers[25][3] ), .B1(n202), .B2(
        \registers[24][3] ), .ZN(n2699) );
  AOI22_X1 U1931 ( .A1(n193), .A2(\registers[29][3] ), .B1(n190), .B2(
        \registers[28][3] ), .ZN(n2700) );
  AOI22_X1 U1932 ( .A1(n217), .A2(\registers[23][4] ), .B1(n214), .B2(
        \registers[22][4] ), .ZN(n2681) );
  AOI22_X1 U1933 ( .A1(n205), .A2(\registers[25][4] ), .B1(n202), .B2(
        \registers[24][4] ), .ZN(n2682) );
  AOI22_X1 U1934 ( .A1(n193), .A2(\registers[29][4] ), .B1(n190), .B2(
        \registers[28][4] ), .ZN(n2683) );
  AOI22_X1 U1935 ( .A1(n217), .A2(\registers[23][5] ), .B1(n214), .B2(
        \registers[22][5] ), .ZN(n2664) );
  AOI22_X1 U1936 ( .A1(n205), .A2(\registers[25][5] ), .B1(n202), .B2(
        \registers[24][5] ), .ZN(n2665) );
  AOI22_X1 U1937 ( .A1(n193), .A2(\registers[29][5] ), .B1(n190), .B2(
        \registers[28][5] ), .ZN(n2666) );
  AOI22_X1 U1938 ( .A1(n217), .A2(\registers[23][6] ), .B1(n214), .B2(
        \registers[22][6] ), .ZN(n2647) );
  AOI22_X1 U1939 ( .A1(n205), .A2(\registers[25][6] ), .B1(n202), .B2(
        \registers[24][6] ), .ZN(n2648) );
  AOI22_X1 U1940 ( .A1(n193), .A2(\registers[29][6] ), .B1(n190), .B2(
        \registers[28][6] ), .ZN(n2649) );
  AOI22_X1 U1941 ( .A1(n217), .A2(\registers[23][7] ), .B1(n214), .B2(
        \registers[22][7] ), .ZN(n2630) );
  AOI22_X1 U1942 ( .A1(n205), .A2(\registers[25][7] ), .B1(n202), .B2(
        \registers[24][7] ), .ZN(n2631) );
  AOI22_X1 U1943 ( .A1(n193), .A2(\registers[29][7] ), .B1(n190), .B2(
        \registers[28][7] ), .ZN(n2632) );
  AOI22_X1 U1944 ( .A1(n217), .A2(\registers[23][8] ), .B1(n214), .B2(
        \registers[22][8] ), .ZN(n2613) );
  AOI22_X1 U1945 ( .A1(n205), .A2(\registers[25][8] ), .B1(n202), .B2(
        \registers[24][8] ), .ZN(n2614) );
  AOI22_X1 U1946 ( .A1(n193), .A2(\registers[29][8] ), .B1(n190), .B2(
        \registers[28][8] ), .ZN(n2615) );
  AOI22_X1 U1947 ( .A1(n217), .A2(\registers[23][9] ), .B1(n214), .B2(
        \registers[22][9] ), .ZN(n2596) );
  AOI22_X1 U1948 ( .A1(n205), .A2(\registers[25][9] ), .B1(n202), .B2(
        \registers[24][9] ), .ZN(n2597) );
  AOI22_X1 U1949 ( .A1(n193), .A2(\registers[29][9] ), .B1(n190), .B2(
        \registers[28][9] ), .ZN(n2598) );
  AOI22_X1 U1950 ( .A1(n217), .A2(\registers[23][10] ), .B1(n214), .B2(
        \registers[22][10] ), .ZN(n2579) );
  AOI22_X1 U1951 ( .A1(n205), .A2(\registers[25][10] ), .B1(n202), .B2(
        \registers[24][10] ), .ZN(n2580) );
  AOI22_X1 U1952 ( .A1(n193), .A2(\registers[29][10] ), .B1(n190), .B2(
        \registers[28][10] ), .ZN(n2581) );
  AOI22_X1 U1953 ( .A1(n218), .A2(\registers[23][11] ), .B1(n215), .B2(
        \registers[22][11] ), .ZN(n2562) );
  AOI22_X1 U1954 ( .A1(n206), .A2(\registers[25][11] ), .B1(n203), .B2(
        \registers[24][11] ), .ZN(n2563) );
  AOI22_X1 U1955 ( .A1(n194), .A2(\registers[29][11] ), .B1(n191), .B2(
        \registers[28][11] ), .ZN(n2564) );
  AOI22_X1 U1956 ( .A1(n218), .A2(\registers[23][12] ), .B1(n215), .B2(
        \registers[22][12] ), .ZN(n2545) );
  AOI22_X1 U1957 ( .A1(n206), .A2(\registers[25][12] ), .B1(n203), .B2(
        \registers[24][12] ), .ZN(n2546) );
  AOI22_X1 U1958 ( .A1(n194), .A2(\registers[29][12] ), .B1(n191), .B2(
        \registers[28][12] ), .ZN(n2547) );
  AOI22_X1 U1959 ( .A1(n218), .A2(\registers[23][13] ), .B1(n215), .B2(
        \registers[22][13] ), .ZN(n2528) );
  AOI22_X1 U1960 ( .A1(n206), .A2(\registers[25][13] ), .B1(n203), .B2(
        \registers[24][13] ), .ZN(n2529) );
  AOI22_X1 U1961 ( .A1(n194), .A2(\registers[29][13] ), .B1(n191), .B2(
        \registers[28][13] ), .ZN(n2530) );
  AOI22_X1 U1962 ( .A1(n218), .A2(\registers[23][14] ), .B1(n215), .B2(
        \registers[22][14] ), .ZN(n2511) );
  AOI22_X1 U1963 ( .A1(n206), .A2(\registers[25][14] ), .B1(n203), .B2(
        \registers[24][14] ), .ZN(n2512) );
  AOI22_X1 U1964 ( .A1(n194), .A2(\registers[29][14] ), .B1(n191), .B2(
        \registers[28][14] ), .ZN(n2513) );
  AOI22_X1 U1965 ( .A1(n218), .A2(\registers[23][15] ), .B1(n215), .B2(
        \registers[22][15] ), .ZN(n2494) );
  AOI22_X1 U1966 ( .A1(n206), .A2(\registers[25][15] ), .B1(n203), .B2(
        \registers[24][15] ), .ZN(n2495) );
  AOI22_X1 U1967 ( .A1(n194), .A2(\registers[29][15] ), .B1(n191), .B2(
        \registers[28][15] ), .ZN(n2496) );
  AOI22_X1 U1968 ( .A1(n218), .A2(\registers[23][16] ), .B1(n215), .B2(
        \registers[22][16] ), .ZN(n2477) );
  AOI22_X1 U1969 ( .A1(n206), .A2(\registers[25][16] ), .B1(n203), .B2(
        \registers[24][16] ), .ZN(n2478) );
  AOI22_X1 U1970 ( .A1(n194), .A2(\registers[29][16] ), .B1(n191), .B2(
        \registers[28][16] ), .ZN(n2479) );
  AOI22_X1 U1971 ( .A1(n218), .A2(\registers[23][17] ), .B1(n215), .B2(
        \registers[22][17] ), .ZN(n2460) );
  AOI22_X1 U1972 ( .A1(n206), .A2(\registers[25][17] ), .B1(n203), .B2(
        \registers[24][17] ), .ZN(n2461) );
  AOI22_X1 U1973 ( .A1(n194), .A2(\registers[29][17] ), .B1(n191), .B2(
        \registers[28][17] ), .ZN(n2462) );
  AOI22_X1 U1974 ( .A1(n218), .A2(\registers[23][18] ), .B1(n215), .B2(
        \registers[22][18] ), .ZN(n2443) );
  AOI22_X1 U1975 ( .A1(n206), .A2(\registers[25][18] ), .B1(n203), .B2(
        \registers[24][18] ), .ZN(n2444) );
  AOI22_X1 U1976 ( .A1(n194), .A2(\registers[29][18] ), .B1(n191), .B2(
        \registers[28][18] ), .ZN(n2445) );
  AOI22_X1 U1977 ( .A1(n218), .A2(\registers[23][19] ), .B1(n215), .B2(
        \registers[22][19] ), .ZN(n2426) );
  AOI22_X1 U1978 ( .A1(n206), .A2(\registers[25][19] ), .B1(n203), .B2(
        \registers[24][19] ), .ZN(n2427) );
  AOI22_X1 U1979 ( .A1(n194), .A2(\registers[29][19] ), .B1(n191), .B2(
        \registers[28][19] ), .ZN(n2428) );
  AOI22_X1 U1980 ( .A1(n218), .A2(\registers[23][20] ), .B1(n215), .B2(
        \registers[22][20] ), .ZN(n2409) );
  AOI22_X1 U1981 ( .A1(n206), .A2(\registers[25][20] ), .B1(n203), .B2(
        \registers[24][20] ), .ZN(n2410) );
  AOI22_X1 U1982 ( .A1(n194), .A2(\registers[29][20] ), .B1(n191), .B2(
        \registers[28][20] ), .ZN(n2411) );
  AOI22_X1 U1983 ( .A1(n218), .A2(\registers[23][21] ), .B1(n215), .B2(
        \registers[22][21] ), .ZN(n2392) );
  AOI22_X1 U1984 ( .A1(n206), .A2(\registers[25][21] ), .B1(n203), .B2(
        \registers[24][21] ), .ZN(n2393) );
  AOI22_X1 U1985 ( .A1(n194), .A2(\registers[29][21] ), .B1(n191), .B2(
        \registers[28][21] ), .ZN(n2394) );
  AOI22_X1 U1986 ( .A1(n219), .A2(\registers[23][22] ), .B1(n216), .B2(
        \registers[22][22] ), .ZN(n2375) );
  AOI22_X1 U1987 ( .A1(n207), .A2(\registers[25][22] ), .B1(n204), .B2(
        \registers[24][22] ), .ZN(n2376) );
  AOI22_X1 U1988 ( .A1(n195), .A2(\registers[29][22] ), .B1(n192), .B2(
        \registers[28][22] ), .ZN(n2377) );
  AOI22_X1 U1989 ( .A1(n219), .A2(\registers[23][23] ), .B1(n216), .B2(
        \registers[22][23] ), .ZN(n2358) );
  AOI22_X1 U1990 ( .A1(n207), .A2(\registers[25][23] ), .B1(n204), .B2(
        \registers[24][23] ), .ZN(n2359) );
  AOI22_X1 U1991 ( .A1(n195), .A2(\registers[29][23] ), .B1(n192), .B2(
        \registers[28][23] ), .ZN(n2360) );
  AOI22_X1 U1992 ( .A1(n219), .A2(\registers[23][24] ), .B1(n216), .B2(
        \registers[22][24] ), .ZN(n2341) );
  AOI22_X1 U1993 ( .A1(n207), .A2(\registers[25][24] ), .B1(n204), .B2(
        \registers[24][24] ), .ZN(n2342) );
  AOI22_X1 U1994 ( .A1(n195), .A2(\registers[29][24] ), .B1(n192), .B2(
        \registers[28][24] ), .ZN(n2343) );
  AOI22_X1 U1995 ( .A1(n219), .A2(\registers[23][25] ), .B1(n216), .B2(
        \registers[22][25] ), .ZN(n2324) );
  AOI22_X1 U1996 ( .A1(n207), .A2(\registers[25][25] ), .B1(n204), .B2(
        \registers[24][25] ), .ZN(n2325) );
  AOI22_X1 U1997 ( .A1(n195), .A2(\registers[29][25] ), .B1(n192), .B2(
        \registers[28][25] ), .ZN(n2326) );
  AOI22_X1 U1998 ( .A1(n219), .A2(\registers[23][26] ), .B1(n216), .B2(
        \registers[22][26] ), .ZN(n2307) );
  AOI22_X1 U1999 ( .A1(n207), .A2(\registers[25][26] ), .B1(n204), .B2(
        \registers[24][26] ), .ZN(n2308) );
  AOI22_X1 U2000 ( .A1(n195), .A2(\registers[29][26] ), .B1(n192), .B2(
        \registers[28][26] ), .ZN(n2309) );
  AOI22_X1 U2001 ( .A1(n219), .A2(\registers[23][27] ), .B1(n216), .B2(
        \registers[22][27] ), .ZN(n2290) );
  AOI22_X1 U2002 ( .A1(n207), .A2(\registers[25][27] ), .B1(n204), .B2(
        \registers[24][27] ), .ZN(n2291) );
  AOI22_X1 U2003 ( .A1(n195), .A2(\registers[29][27] ), .B1(n192), .B2(
        \registers[28][27] ), .ZN(n2292) );
  AOI22_X1 U2004 ( .A1(n219), .A2(\registers[23][28] ), .B1(n216), .B2(
        \registers[22][28] ), .ZN(n2273) );
  AOI22_X1 U2005 ( .A1(n207), .A2(\registers[25][28] ), .B1(n204), .B2(
        \registers[24][28] ), .ZN(n2274) );
  AOI22_X1 U2006 ( .A1(n195), .A2(\registers[29][28] ), .B1(n192), .B2(
        \registers[28][28] ), .ZN(n2275) );
  AOI22_X1 U2007 ( .A1(n219), .A2(\registers[23][29] ), .B1(n216), .B2(
        \registers[22][29] ), .ZN(n2256) );
  AOI22_X1 U2008 ( .A1(n207), .A2(\registers[25][29] ), .B1(n204), .B2(
        \registers[24][29] ), .ZN(n2257) );
  AOI22_X1 U2009 ( .A1(n195), .A2(\registers[29][29] ), .B1(n192), .B2(
        \registers[28][29] ), .ZN(n2258) );
  AOI22_X1 U2010 ( .A1(n219), .A2(\registers[23][30] ), .B1(n216), .B2(
        \registers[22][30] ), .ZN(n2239) );
  AOI22_X1 U2011 ( .A1(n207), .A2(\registers[25][30] ), .B1(n204), .B2(
        \registers[24][30] ), .ZN(n2240) );
  AOI22_X1 U2012 ( .A1(n195), .A2(\registers[29][30] ), .B1(n192), .B2(
        \registers[28][30] ), .ZN(n2241) );
  AOI22_X1 U2013 ( .A1(n219), .A2(\registers[23][31] ), .B1(n216), .B2(
        \registers[22][31] ), .ZN(n2197) );
  AOI22_X1 U2014 ( .A1(n207), .A2(\registers[25][31] ), .B1(n204), .B2(
        \registers[24][31] ), .ZN(n2202) );
  AOI22_X1 U2015 ( .A1(n195), .A2(\registers[29][31] ), .B1(n192), .B2(
        \registers[28][31] ), .ZN(n2207) );
  OAI221_X1 U2016 ( .B1(n160), .B2(n178), .C1(n128), .C2(n175), .A(n2766), 
        .ZN(n2762) );
  AOI22_X1 U2017 ( .A1(n172), .A2(\registers[7][0] ), .B1(n169), .B2(
        \registers[6][0] ), .ZN(n2766) );
  OAI221_X1 U2018 ( .B1(n159), .B2(n178), .C1(n127), .C2(n175), .A(n2737), 
        .ZN(n2735) );
  AOI22_X1 U2019 ( .A1(n172), .A2(\registers[7][1] ), .B1(n169), .B2(
        \registers[6][1] ), .ZN(n2737) );
  OAI221_X1 U2020 ( .B1(n158), .B2(n178), .C1(n126), .C2(n175), .A(n2720), 
        .ZN(n2718) );
  AOI22_X1 U2021 ( .A1(n172), .A2(\registers[7][2] ), .B1(n169), .B2(
        \registers[6][2] ), .ZN(n2720) );
  OAI221_X1 U2022 ( .B1(n157), .B2(n178), .C1(n125), .C2(n175), .A(n2703), 
        .ZN(n2701) );
  AOI22_X1 U2023 ( .A1(n172), .A2(\registers[7][3] ), .B1(n169), .B2(
        \registers[6][3] ), .ZN(n2703) );
  OAI221_X1 U2024 ( .B1(n156), .B2(n178), .C1(n124), .C2(n175), .A(n2686), 
        .ZN(n2684) );
  AOI22_X1 U2025 ( .A1(n172), .A2(\registers[7][4] ), .B1(n169), .B2(
        \registers[6][4] ), .ZN(n2686) );
  OAI221_X1 U2026 ( .B1(n155), .B2(n178), .C1(n123), .C2(n175), .A(n2669), 
        .ZN(n2667) );
  AOI22_X1 U2027 ( .A1(n172), .A2(\registers[7][5] ), .B1(n169), .B2(
        \registers[6][5] ), .ZN(n2669) );
  OAI221_X1 U2028 ( .B1(n154), .B2(n178), .C1(n122), .C2(n175), .A(n2652), 
        .ZN(n2650) );
  AOI22_X1 U2029 ( .A1(n172), .A2(\registers[7][6] ), .B1(n169), .B2(
        \registers[6][6] ), .ZN(n2652) );
  OAI221_X1 U2030 ( .B1(n153), .B2(n178), .C1(n121), .C2(n175), .A(n2635), 
        .ZN(n2633) );
  AOI22_X1 U2031 ( .A1(n172), .A2(\registers[7][7] ), .B1(n169), .B2(
        \registers[6][7] ), .ZN(n2635) );
  OAI221_X1 U2032 ( .B1(n152), .B2(n178), .C1(n120), .C2(n175), .A(n2618), 
        .ZN(n2616) );
  AOI22_X1 U2033 ( .A1(n172), .A2(\registers[7][8] ), .B1(n169), .B2(
        \registers[6][8] ), .ZN(n2618) );
  OAI221_X1 U2034 ( .B1(n151), .B2(n178), .C1(n119), .C2(n175), .A(n2601), 
        .ZN(n2599) );
  AOI22_X1 U2035 ( .A1(n172), .A2(\registers[7][9] ), .B1(n169), .B2(
        \registers[6][9] ), .ZN(n2601) );
  OAI221_X1 U2036 ( .B1(n150), .B2(n178), .C1(n118), .C2(n175), .A(n2584), 
        .ZN(n2582) );
  AOI22_X1 U2037 ( .A1(n172), .A2(\registers[7][10] ), .B1(n169), .B2(
        \registers[6][10] ), .ZN(n2584) );
  OAI221_X1 U2038 ( .B1(n149), .B2(n179), .C1(n117), .C2(n176), .A(n2567), 
        .ZN(n2565) );
  AOI22_X1 U2039 ( .A1(n173), .A2(\registers[7][11] ), .B1(n170), .B2(
        \registers[6][11] ), .ZN(n2567) );
  OAI221_X1 U2040 ( .B1(n148), .B2(n179), .C1(n116), .C2(n176), .A(n2550), 
        .ZN(n2548) );
  AOI22_X1 U2041 ( .A1(n173), .A2(\registers[7][12] ), .B1(n170), .B2(
        \registers[6][12] ), .ZN(n2550) );
  OAI221_X1 U2042 ( .B1(n147), .B2(n179), .C1(n115), .C2(n176), .A(n2533), 
        .ZN(n2531) );
  AOI22_X1 U2043 ( .A1(n173), .A2(\registers[7][13] ), .B1(n170), .B2(
        \registers[6][13] ), .ZN(n2533) );
  OAI221_X1 U2044 ( .B1(n146), .B2(n179), .C1(n114), .C2(n176), .A(n2516), 
        .ZN(n2514) );
  AOI22_X1 U2045 ( .A1(n173), .A2(\registers[7][14] ), .B1(n170), .B2(
        \registers[6][14] ), .ZN(n2516) );
  OAI221_X1 U2046 ( .B1(n145), .B2(n179), .C1(n113), .C2(n176), .A(n2499), 
        .ZN(n2497) );
  AOI22_X1 U2047 ( .A1(n173), .A2(\registers[7][15] ), .B1(n170), .B2(
        \registers[6][15] ), .ZN(n2499) );
  OAI221_X1 U2048 ( .B1(n144), .B2(n179), .C1(n112), .C2(n176), .A(n2482), 
        .ZN(n2480) );
  AOI22_X1 U2049 ( .A1(n173), .A2(\registers[7][16] ), .B1(n170), .B2(
        \registers[6][16] ), .ZN(n2482) );
  OAI221_X1 U2050 ( .B1(n143), .B2(n179), .C1(n111), .C2(n176), .A(n2465), 
        .ZN(n2463) );
  AOI22_X1 U2051 ( .A1(n173), .A2(\registers[7][17] ), .B1(n170), .B2(
        \registers[6][17] ), .ZN(n2465) );
  OAI221_X1 U2052 ( .B1(n142), .B2(n179), .C1(n110), .C2(n176), .A(n2448), 
        .ZN(n2446) );
  AOI22_X1 U2053 ( .A1(n173), .A2(\registers[7][18] ), .B1(n170), .B2(
        \registers[6][18] ), .ZN(n2448) );
  OAI221_X1 U2054 ( .B1(n141), .B2(n179), .C1(n109), .C2(n176), .A(n2431), 
        .ZN(n2429) );
  AOI22_X1 U2055 ( .A1(n173), .A2(\registers[7][19] ), .B1(n170), .B2(
        \registers[6][19] ), .ZN(n2431) );
  OAI221_X1 U2056 ( .B1(n140), .B2(n179), .C1(n108), .C2(n176), .A(n2414), 
        .ZN(n2412) );
  AOI22_X1 U2057 ( .A1(n173), .A2(\registers[7][20] ), .B1(n170), .B2(
        \registers[6][20] ), .ZN(n2414) );
  OAI221_X1 U2058 ( .B1(n139), .B2(n179), .C1(n107), .C2(n176), .A(n2397), 
        .ZN(n2395) );
  AOI22_X1 U2059 ( .A1(n173), .A2(\registers[7][21] ), .B1(n170), .B2(
        \registers[6][21] ), .ZN(n2397) );
  AND2_X1 U2060 ( .A1(ADD_RD2[0]), .A2(n2170), .ZN(n2168) );
  AND2_X1 U2061 ( .A1(ADD_RD1[0]), .A2(n2761), .ZN(n2759) );
  NAND4_X1 U2062 ( .A1(n2149), .A2(n2150), .A3(n2151), .A4(n2152), .ZN(N320)
         );
  AOI221_X1 U2063 ( .B1(n247), .B2(\registers[9][0] ), .C1(n244), .C2(
        \registers[8][0] ), .A(n2180), .ZN(n2149) );
  AOI221_X1 U2064 ( .B1(n259), .B2(\registers[13][0] ), .C1(n256), .C2(
        \registers[12][0] ), .A(n2177), .ZN(n2150) );
  AOI211_X1 U2065 ( .C1(n280), .C2(\registers[1][0] ), .A(n2171), .B(n2172), 
        .ZN(n2151) );
  NAND4_X1 U2066 ( .A1(n2132), .A2(n2133), .A3(n2134), .A4(n2135), .ZN(N321)
         );
  AOI221_X1 U2067 ( .B1(n247), .B2(\registers[9][1] ), .C1(n244), .C2(
        \registers[8][1] ), .A(n2148), .ZN(n2132) );
  AOI221_X1 U2068 ( .B1(n259), .B2(\registers[13][1] ), .C1(n256), .C2(
        \registers[12][1] ), .A(n2147), .ZN(n2133) );
  AOI211_X1 U2069 ( .C1(n280), .C2(\registers[1][1] ), .A(n2144), .B(n2145), 
        .ZN(n2134) );
  NAND4_X1 U2070 ( .A1(n2115), .A2(n2116), .A3(n2117), .A4(n2118), .ZN(N322)
         );
  AOI221_X1 U2071 ( .B1(n247), .B2(\registers[9][2] ), .C1(n244), .C2(
        \registers[8][2] ), .A(n2131), .ZN(n2115) );
  AOI221_X1 U2072 ( .B1(n259), .B2(\registers[13][2] ), .C1(n256), .C2(
        \registers[12][2] ), .A(n2130), .ZN(n2116) );
  AOI211_X1 U2073 ( .C1(n280), .C2(\registers[1][2] ), .A(n2127), .B(n2128), 
        .ZN(n2117) );
  NAND4_X1 U2074 ( .A1(n2098), .A2(n2099), .A3(n2100), .A4(n2101), .ZN(N323)
         );
  AOI221_X1 U2075 ( .B1(n247), .B2(\registers[9][3] ), .C1(n244), .C2(
        \registers[8][3] ), .A(n2114), .ZN(n2098) );
  AOI221_X1 U2076 ( .B1(n259), .B2(\registers[13][3] ), .C1(n256), .C2(
        \registers[12][3] ), .A(n2113), .ZN(n2099) );
  AOI211_X1 U2077 ( .C1(n280), .C2(\registers[1][3] ), .A(n2110), .B(n2111), 
        .ZN(n2100) );
  NAND4_X1 U2078 ( .A1(n2081), .A2(n2082), .A3(n2083), .A4(n2084), .ZN(N324)
         );
  AOI221_X1 U2079 ( .B1(n247), .B2(\registers[9][4] ), .C1(n244), .C2(
        \registers[8][4] ), .A(n2097), .ZN(n2081) );
  AOI221_X1 U2080 ( .B1(n259), .B2(\registers[13][4] ), .C1(n256), .C2(
        \registers[12][4] ), .A(n2096), .ZN(n2082) );
  AOI211_X1 U2081 ( .C1(n280), .C2(\registers[1][4] ), .A(n2093), .B(n2094), 
        .ZN(n2083) );
  NAND4_X1 U2082 ( .A1(n2064), .A2(n2065), .A3(n2066), .A4(n2067), .ZN(N325)
         );
  AOI221_X1 U2083 ( .B1(n247), .B2(\registers[9][5] ), .C1(n244), .C2(
        \registers[8][5] ), .A(n2080), .ZN(n2064) );
  AOI221_X1 U2084 ( .B1(n259), .B2(\registers[13][5] ), .C1(n256), .C2(
        \registers[12][5] ), .A(n2079), .ZN(n2065) );
  AOI211_X1 U2085 ( .C1(n280), .C2(\registers[1][5] ), .A(n2076), .B(n2077), 
        .ZN(n2066) );
  NAND4_X1 U2086 ( .A1(n2047), .A2(n2048), .A3(n2049), .A4(n2050), .ZN(N326)
         );
  AOI221_X1 U2087 ( .B1(n247), .B2(\registers[9][6] ), .C1(n244), .C2(
        \registers[8][6] ), .A(n2063), .ZN(n2047) );
  AOI221_X1 U2088 ( .B1(n259), .B2(\registers[13][6] ), .C1(n256), .C2(
        \registers[12][6] ), .A(n2062), .ZN(n2048) );
  AOI211_X1 U2089 ( .C1(n280), .C2(\registers[1][6] ), .A(n2059), .B(n2060), 
        .ZN(n2049) );
  NAND4_X1 U2090 ( .A1(n2030), .A2(n2031), .A3(n2032), .A4(n2033), .ZN(N327)
         );
  AOI221_X1 U2091 ( .B1(n247), .B2(\registers[9][7] ), .C1(n244), .C2(
        \registers[8][7] ), .A(n2046), .ZN(n2030) );
  AOI221_X1 U2092 ( .B1(n259), .B2(\registers[13][7] ), .C1(n256), .C2(
        \registers[12][7] ), .A(n2045), .ZN(n2031) );
  AOI211_X1 U2093 ( .C1(n280), .C2(\registers[1][7] ), .A(n2042), .B(n2043), 
        .ZN(n2032) );
  NAND4_X1 U2094 ( .A1(n2013), .A2(n2014), .A3(n2015), .A4(n2016), .ZN(N328)
         );
  AOI221_X1 U2095 ( .B1(n247), .B2(\registers[9][8] ), .C1(n244), .C2(
        \registers[8][8] ), .A(n2029), .ZN(n2013) );
  AOI221_X1 U2096 ( .B1(n259), .B2(\registers[13][8] ), .C1(n256), .C2(
        \registers[12][8] ), .A(n2028), .ZN(n2014) );
  AOI211_X1 U2097 ( .C1(n280), .C2(\registers[1][8] ), .A(n2025), .B(n2026), 
        .ZN(n2015) );
  NAND4_X1 U2098 ( .A1(n1996), .A2(n1997), .A3(n1998), .A4(n1999), .ZN(N329)
         );
  AOI221_X1 U2099 ( .B1(n247), .B2(\registers[9][9] ), .C1(n244), .C2(
        \registers[8][9] ), .A(n2012), .ZN(n1996) );
  AOI221_X1 U2100 ( .B1(n259), .B2(\registers[13][9] ), .C1(n256), .C2(
        \registers[12][9] ), .A(n2011), .ZN(n1997) );
  AOI211_X1 U2101 ( .C1(n280), .C2(\registers[1][9] ), .A(n2008), .B(n2009), 
        .ZN(n1998) );
  NAND4_X1 U2102 ( .A1(n1979), .A2(n1980), .A3(n1981), .A4(n1982), .ZN(N330)
         );
  AOI221_X1 U2103 ( .B1(n247), .B2(\registers[9][10] ), .C1(n244), .C2(
        \registers[8][10] ), .A(n1995), .ZN(n1979) );
  AOI221_X1 U2104 ( .B1(n259), .B2(\registers[13][10] ), .C1(n256), .C2(
        \registers[12][10] ), .A(n1994), .ZN(n1980) );
  AOI211_X1 U2105 ( .C1(n280), .C2(\registers[1][10] ), .A(n1991), .B(n1992), 
        .ZN(n1981) );
  NAND4_X1 U2106 ( .A1(n1962), .A2(n1963), .A3(n1964), .A4(n1965), .ZN(N331)
         );
  AOI221_X1 U2107 ( .B1(n248), .B2(\registers[9][11] ), .C1(n245), .C2(
        \registers[8][11] ), .A(n1978), .ZN(n1962) );
  AOI221_X1 U2108 ( .B1(n260), .B2(\registers[13][11] ), .C1(n257), .C2(
        \registers[12][11] ), .A(n1977), .ZN(n1963) );
  AOI211_X1 U2109 ( .C1(n281), .C2(\registers[1][11] ), .A(n1974), .B(n1975), 
        .ZN(n1964) );
  NAND4_X1 U2110 ( .A1(n1945), .A2(n1946), .A3(n1947), .A4(n1948), .ZN(N332)
         );
  AOI221_X1 U2111 ( .B1(n248), .B2(\registers[9][12] ), .C1(n245), .C2(
        \registers[8][12] ), .A(n1961), .ZN(n1945) );
  AOI221_X1 U2112 ( .B1(n260), .B2(\registers[13][12] ), .C1(n257), .C2(
        \registers[12][12] ), .A(n1960), .ZN(n1946) );
  AOI211_X1 U2113 ( .C1(n281), .C2(\registers[1][12] ), .A(n1957), .B(n1958), 
        .ZN(n1947) );
  NAND4_X1 U2114 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .ZN(N333)
         );
  AOI221_X1 U2115 ( .B1(n248), .B2(\registers[9][13] ), .C1(n245), .C2(
        \registers[8][13] ), .A(n1944), .ZN(n1928) );
  AOI221_X1 U2116 ( .B1(n260), .B2(\registers[13][13] ), .C1(n257), .C2(
        \registers[12][13] ), .A(n1943), .ZN(n1929) );
  AOI211_X1 U2117 ( .C1(n281), .C2(\registers[1][13] ), .A(n1940), .B(n1941), 
        .ZN(n1930) );
  NAND4_X1 U2118 ( .A1(n1911), .A2(n1912), .A3(n1913), .A4(n1914), .ZN(N334)
         );
  AOI221_X1 U2119 ( .B1(n248), .B2(\registers[9][14] ), .C1(n245), .C2(
        \registers[8][14] ), .A(n1927), .ZN(n1911) );
  AOI221_X1 U2120 ( .B1(n260), .B2(\registers[13][14] ), .C1(n257), .C2(
        \registers[12][14] ), .A(n1926), .ZN(n1912) );
  AOI211_X1 U2121 ( .C1(n281), .C2(\registers[1][14] ), .A(n1923), .B(n1924), 
        .ZN(n1913) );
  NAND4_X1 U2122 ( .A1(n1894), .A2(n1895), .A3(n1896), .A4(n1897), .ZN(N335)
         );
  AOI221_X1 U2123 ( .B1(n248), .B2(\registers[9][15] ), .C1(n245), .C2(
        \registers[8][15] ), .A(n1910), .ZN(n1894) );
  AOI221_X1 U2124 ( .B1(n260), .B2(\registers[13][15] ), .C1(n257), .C2(
        \registers[12][15] ), .A(n1909), .ZN(n1895) );
  AOI211_X1 U2125 ( .C1(n281), .C2(\registers[1][15] ), .A(n1906), .B(n1907), 
        .ZN(n1896) );
  NAND4_X1 U2126 ( .A1(n1877), .A2(n1878), .A3(n1879), .A4(n1880), .ZN(N336)
         );
  AOI221_X1 U2127 ( .B1(n248), .B2(\registers[9][16] ), .C1(n245), .C2(
        \registers[8][16] ), .A(n1893), .ZN(n1877) );
  AOI221_X1 U2128 ( .B1(n260), .B2(\registers[13][16] ), .C1(n257), .C2(
        \registers[12][16] ), .A(n1892), .ZN(n1878) );
  AOI211_X1 U2129 ( .C1(n281), .C2(\registers[1][16] ), .A(n1889), .B(n1890), 
        .ZN(n1879) );
  NAND4_X1 U2130 ( .A1(n1860), .A2(n1861), .A3(n1862), .A4(n1863), .ZN(N337)
         );
  AOI221_X1 U2131 ( .B1(n248), .B2(\registers[9][17] ), .C1(n245), .C2(
        \registers[8][17] ), .A(n1876), .ZN(n1860) );
  AOI221_X1 U2132 ( .B1(n260), .B2(\registers[13][17] ), .C1(n257), .C2(
        \registers[12][17] ), .A(n1875), .ZN(n1861) );
  AOI211_X1 U2133 ( .C1(n281), .C2(\registers[1][17] ), .A(n1872), .B(n1873), 
        .ZN(n1862) );
  NAND4_X1 U2134 ( .A1(n1843), .A2(n1844), .A3(n1845), .A4(n1846), .ZN(N338)
         );
  AOI221_X1 U2135 ( .B1(n248), .B2(\registers[9][18] ), .C1(n245), .C2(
        \registers[8][18] ), .A(n1859), .ZN(n1843) );
  AOI221_X1 U2136 ( .B1(n260), .B2(\registers[13][18] ), .C1(n257), .C2(
        \registers[12][18] ), .A(n1858), .ZN(n1844) );
  AOI211_X1 U2137 ( .C1(n281), .C2(\registers[1][18] ), .A(n1855), .B(n1856), 
        .ZN(n1845) );
  NAND4_X1 U2138 ( .A1(n1826), .A2(n1827), .A3(n1828), .A4(n1829), .ZN(N339)
         );
  AOI221_X1 U2139 ( .B1(n248), .B2(\registers[9][19] ), .C1(n245), .C2(
        \registers[8][19] ), .A(n1842), .ZN(n1826) );
  AOI221_X1 U2140 ( .B1(n260), .B2(\registers[13][19] ), .C1(n257), .C2(
        \registers[12][19] ), .A(n1841), .ZN(n1827) );
  AOI211_X1 U2141 ( .C1(n281), .C2(\registers[1][19] ), .A(n1838), .B(n1839), 
        .ZN(n1828) );
  NAND4_X1 U2142 ( .A1(n1809), .A2(n1810), .A3(n1811), .A4(n1812), .ZN(N340)
         );
  AOI221_X1 U2143 ( .B1(n248), .B2(\registers[9][20] ), .C1(n245), .C2(
        \registers[8][20] ), .A(n1825), .ZN(n1809) );
  AOI221_X1 U2144 ( .B1(n260), .B2(\registers[13][20] ), .C1(n257), .C2(
        \registers[12][20] ), .A(n1824), .ZN(n1810) );
  AOI211_X1 U2145 ( .C1(n281), .C2(\registers[1][20] ), .A(n1821), .B(n1822), 
        .ZN(n1811) );
  NAND4_X1 U2146 ( .A1(n1792), .A2(n1793), .A3(n1794), .A4(n1795), .ZN(N341)
         );
  AOI221_X1 U2147 ( .B1(n248), .B2(\registers[9][21] ), .C1(n245), .C2(
        \registers[8][21] ), .A(n1808), .ZN(n1792) );
  AOI221_X1 U2148 ( .B1(n260), .B2(\registers[13][21] ), .C1(n257), .C2(
        \registers[12][21] ), .A(n1807), .ZN(n1793) );
  AOI211_X1 U2149 ( .C1(n281), .C2(\registers[1][21] ), .A(n1804), .B(n1805), 
        .ZN(n1794) );
  NAND4_X1 U2150 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .ZN(N342)
         );
  AOI221_X1 U2151 ( .B1(n249), .B2(\registers[9][22] ), .C1(n246), .C2(
        \registers[8][22] ), .A(n1791), .ZN(n1775) );
  AOI221_X1 U2152 ( .B1(n261), .B2(\registers[13][22] ), .C1(n258), .C2(
        \registers[12][22] ), .A(n1790), .ZN(n1776) );
  AOI211_X1 U2153 ( .C1(n282), .C2(\registers[1][22] ), .A(n1787), .B(n1788), 
        .ZN(n1777) );
  NAND4_X1 U2154 ( .A1(n1758), .A2(n1759), .A3(n1760), .A4(n1761), .ZN(N343)
         );
  AOI221_X1 U2155 ( .B1(n249), .B2(\registers[9][23] ), .C1(n246), .C2(
        \registers[8][23] ), .A(n1774), .ZN(n1758) );
  AOI221_X1 U2156 ( .B1(n261), .B2(\registers[13][23] ), .C1(n258), .C2(
        \registers[12][23] ), .A(n1773), .ZN(n1759) );
  AOI211_X1 U2157 ( .C1(n282), .C2(\registers[1][23] ), .A(n1770), .B(n1771), 
        .ZN(n1760) );
  NAND4_X1 U2158 ( .A1(n1741), .A2(n1742), .A3(n1743), .A4(n1744), .ZN(N344)
         );
  AOI221_X1 U2159 ( .B1(n261), .B2(\registers[13][24] ), .C1(n258), .C2(
        \registers[12][24] ), .A(n1756), .ZN(n1742) );
  AOI221_X1 U2160 ( .B1(n249), .B2(\registers[9][24] ), .C1(n246), .C2(
        \registers[8][24] ), .A(n1757), .ZN(n1741) );
  AOI211_X1 U2161 ( .C1(n282), .C2(\registers[1][24] ), .A(n1753), .B(n1754), 
        .ZN(n1743) );
  NAND4_X1 U2162 ( .A1(n1724), .A2(n1725), .A3(n1726), .A4(n1727), .ZN(N345)
         );
  AOI221_X1 U2163 ( .B1(n261), .B2(\registers[13][25] ), .C1(n258), .C2(
        \registers[12][25] ), .A(n1739), .ZN(n1725) );
  AOI221_X1 U2164 ( .B1(n249), .B2(\registers[9][25] ), .C1(n246), .C2(
        \registers[8][25] ), .A(n1740), .ZN(n1724) );
  AOI211_X1 U2165 ( .C1(n282), .C2(\registers[1][25] ), .A(n1736), .B(n1737), 
        .ZN(n1726) );
  NAND4_X1 U2166 ( .A1(n1707), .A2(n1708), .A3(n1709), .A4(n1710), .ZN(N346)
         );
  AOI221_X1 U2167 ( .B1(n261), .B2(\registers[13][26] ), .C1(n258), .C2(
        \registers[12][26] ), .A(n1722), .ZN(n1708) );
  AOI221_X1 U2168 ( .B1(n249), .B2(\registers[9][26] ), .C1(n246), .C2(
        \registers[8][26] ), .A(n1723), .ZN(n1707) );
  AOI211_X1 U2169 ( .C1(n282), .C2(\registers[1][26] ), .A(n1719), .B(n1720), 
        .ZN(n1709) );
  NAND4_X1 U2170 ( .A1(n1690), .A2(n1691), .A3(n1692), .A4(n1693), .ZN(N347)
         );
  AOI221_X1 U2171 ( .B1(n261), .B2(\registers[13][27] ), .C1(n258), .C2(
        \registers[12][27] ), .A(n1705), .ZN(n1691) );
  AOI221_X1 U2172 ( .B1(n249), .B2(\registers[9][27] ), .C1(n246), .C2(
        \registers[8][27] ), .A(n1706), .ZN(n1690) );
  AOI211_X1 U2173 ( .C1(n282), .C2(\registers[1][27] ), .A(n1702), .B(n1703), 
        .ZN(n1692) );
  NAND4_X1 U2174 ( .A1(n1673), .A2(n1674), .A3(n1675), .A4(n1676), .ZN(N348)
         );
  AOI221_X1 U2175 ( .B1(n261), .B2(\registers[13][28] ), .C1(n258), .C2(
        \registers[12][28] ), .A(n1688), .ZN(n1674) );
  AOI221_X1 U2176 ( .B1(n249), .B2(\registers[9][28] ), .C1(n246), .C2(
        \registers[8][28] ), .A(n1689), .ZN(n1673) );
  AOI211_X1 U2177 ( .C1(n282), .C2(\registers[1][28] ), .A(n1685), .B(n1686), 
        .ZN(n1675) );
  NAND4_X1 U2178 ( .A1(n1656), .A2(n1657), .A3(n1658), .A4(n1659), .ZN(N349)
         );
  AOI221_X1 U2179 ( .B1(n261), .B2(\registers[13][29] ), .C1(n258), .C2(
        \registers[12][29] ), .A(n1671), .ZN(n1657) );
  AOI221_X1 U2180 ( .B1(n249), .B2(\registers[9][29] ), .C1(n246), .C2(
        \registers[8][29] ), .A(n1672), .ZN(n1656) );
  AOI211_X1 U2181 ( .C1(n282), .C2(\registers[1][29] ), .A(n1668), .B(n1669), 
        .ZN(n1658) );
  NAND4_X1 U2182 ( .A1(n1639), .A2(n1640), .A3(n1641), .A4(n1642), .ZN(N350)
         );
  AOI221_X1 U2183 ( .B1(n261), .B2(\registers[13][30] ), .C1(n258), .C2(
        \registers[12][30] ), .A(n1654), .ZN(n1640) );
  AOI221_X1 U2184 ( .B1(n249), .B2(\registers[9][30] ), .C1(n246), .C2(
        \registers[8][30] ), .A(n1655), .ZN(n1639) );
  AOI211_X1 U2185 ( .C1(n282), .C2(\registers[1][30] ), .A(n1651), .B(n1652), 
        .ZN(n1641) );
  NAND4_X1 U2186 ( .A1(n1591), .A2(n1592), .A3(n1593), .A4(n1594), .ZN(N351)
         );
  AOI221_X1 U2187 ( .B1(n261), .B2(\registers[13][31] ), .C1(n258), .C2(
        \registers[12][31] ), .A(n1631), .ZN(n1592) );
  AOI221_X1 U2188 ( .B1(n249), .B2(\registers[9][31] ), .C1(n246), .C2(
        \registers[8][31] ), .A(n1636), .ZN(n1591) );
  AOI211_X1 U2189 ( .C1(n282), .C2(\registers[1][31] ), .A(n1620), .B(n1621), 
        .ZN(n1593) );
  NAND4_X1 U2190 ( .A1(n2740), .A2(n2741), .A3(n2742), .A4(n2743), .ZN(N185)
         );
  AOI221_X1 U2191 ( .B1(n166), .B2(\registers[13][0] ), .C1(n163), .C2(
        \registers[12][0] ), .A(n2768), .ZN(n2741) );
  AOI221_X1 U2192 ( .B1(n26), .B2(\registers[9][0] ), .C1(n23), .C2(
        \registers[8][0] ), .A(n2771), .ZN(n2740) );
  AOI211_X1 U2193 ( .C1(n187), .C2(\registers[1][0] ), .A(n2762), .B(n2763), 
        .ZN(n2742) );
  NAND4_X1 U2194 ( .A1(n2723), .A2(n2724), .A3(n2725), .A4(n2726), .ZN(N186)
         );
  AOI221_X1 U2195 ( .B1(n166), .B2(\registers[13][1] ), .C1(n163), .C2(
        \registers[12][1] ), .A(n2738), .ZN(n2724) );
  AOI221_X1 U2196 ( .B1(n26), .B2(\registers[9][1] ), .C1(n23), .C2(
        \registers[8][1] ), .A(n2739), .ZN(n2723) );
  AOI211_X1 U2197 ( .C1(n187), .C2(\registers[1][1] ), .A(n2735), .B(n2736), 
        .ZN(n2725) );
  NAND4_X1 U2198 ( .A1(n2706), .A2(n2707), .A3(n2708), .A4(n2709), .ZN(N187)
         );
  AOI221_X1 U2199 ( .B1(n166), .B2(\registers[13][2] ), .C1(n163), .C2(
        \registers[12][2] ), .A(n2721), .ZN(n2707) );
  AOI221_X1 U2200 ( .B1(n26), .B2(\registers[9][2] ), .C1(n23), .C2(
        \registers[8][2] ), .A(n2722), .ZN(n2706) );
  AOI211_X1 U2201 ( .C1(n187), .C2(\registers[1][2] ), .A(n2718), .B(n2719), 
        .ZN(n2708) );
  NAND4_X1 U2202 ( .A1(n2689), .A2(n2690), .A3(n2691), .A4(n2692), .ZN(N188)
         );
  AOI221_X1 U2203 ( .B1(n166), .B2(\registers[13][3] ), .C1(n163), .C2(
        \registers[12][3] ), .A(n2704), .ZN(n2690) );
  AOI221_X1 U2204 ( .B1(n26), .B2(\registers[9][3] ), .C1(n23), .C2(
        \registers[8][3] ), .A(n2705), .ZN(n2689) );
  AOI211_X1 U2205 ( .C1(n187), .C2(\registers[1][3] ), .A(n2701), .B(n2702), 
        .ZN(n2691) );
  NAND4_X1 U2206 ( .A1(n2672), .A2(n2673), .A3(n2674), .A4(n2675), .ZN(N189)
         );
  AOI221_X1 U2207 ( .B1(n166), .B2(\registers[13][4] ), .C1(n163), .C2(
        \registers[12][4] ), .A(n2687), .ZN(n2673) );
  AOI221_X1 U2208 ( .B1(n26), .B2(\registers[9][4] ), .C1(n23), .C2(
        \registers[8][4] ), .A(n2688), .ZN(n2672) );
  AOI211_X1 U2209 ( .C1(n187), .C2(\registers[1][4] ), .A(n2684), .B(n2685), 
        .ZN(n2674) );
  NAND4_X1 U2210 ( .A1(n2655), .A2(n2656), .A3(n2657), .A4(n2658), .ZN(N190)
         );
  AOI221_X1 U2211 ( .B1(n166), .B2(\registers[13][5] ), .C1(n163), .C2(
        \registers[12][5] ), .A(n2670), .ZN(n2656) );
  AOI221_X1 U2212 ( .B1(n26), .B2(\registers[9][5] ), .C1(n23), .C2(
        \registers[8][5] ), .A(n2671), .ZN(n2655) );
  AOI211_X1 U2213 ( .C1(n187), .C2(\registers[1][5] ), .A(n2667), .B(n2668), 
        .ZN(n2657) );
  NAND4_X1 U2214 ( .A1(n2638), .A2(n2639), .A3(n2640), .A4(n2641), .ZN(N191)
         );
  AOI221_X1 U2215 ( .B1(n166), .B2(\registers[13][6] ), .C1(n163), .C2(
        \registers[12][6] ), .A(n2653), .ZN(n2639) );
  AOI221_X1 U2216 ( .B1(n26), .B2(\registers[9][6] ), .C1(n23), .C2(
        \registers[8][6] ), .A(n2654), .ZN(n2638) );
  AOI211_X1 U2217 ( .C1(n187), .C2(\registers[1][6] ), .A(n2650), .B(n2651), 
        .ZN(n2640) );
  NAND4_X1 U2218 ( .A1(n2621), .A2(n2622), .A3(n2623), .A4(n2624), .ZN(N192)
         );
  AOI221_X1 U2219 ( .B1(n166), .B2(\registers[13][7] ), .C1(n163), .C2(
        \registers[12][7] ), .A(n2636), .ZN(n2622) );
  AOI221_X1 U2220 ( .B1(n26), .B2(\registers[9][7] ), .C1(n23), .C2(
        \registers[8][7] ), .A(n2637), .ZN(n2621) );
  AOI211_X1 U2221 ( .C1(n187), .C2(\registers[1][7] ), .A(n2633), .B(n2634), 
        .ZN(n2623) );
  NAND4_X1 U2222 ( .A1(n2604), .A2(n2605), .A3(n2606), .A4(n2607), .ZN(N193)
         );
  AOI221_X1 U2223 ( .B1(n166), .B2(\registers[13][8] ), .C1(n163), .C2(
        \registers[12][8] ), .A(n2619), .ZN(n2605) );
  AOI221_X1 U2224 ( .B1(n26), .B2(\registers[9][8] ), .C1(n23), .C2(
        \registers[8][8] ), .A(n2620), .ZN(n2604) );
  AOI211_X1 U2225 ( .C1(n187), .C2(\registers[1][8] ), .A(n2616), .B(n2617), 
        .ZN(n2606) );
  NAND4_X1 U2226 ( .A1(n2587), .A2(n2588), .A3(n2589), .A4(n2590), .ZN(N194)
         );
  AOI221_X1 U2227 ( .B1(n166), .B2(\registers[13][9] ), .C1(n163), .C2(
        \registers[12][9] ), .A(n2602), .ZN(n2588) );
  AOI221_X1 U2228 ( .B1(n26), .B2(\registers[9][9] ), .C1(n23), .C2(
        \registers[8][9] ), .A(n2603), .ZN(n2587) );
  AOI211_X1 U2229 ( .C1(n187), .C2(\registers[1][9] ), .A(n2599), .B(n2600), 
        .ZN(n2589) );
  NAND4_X1 U2230 ( .A1(n2570), .A2(n2571), .A3(n2572), .A4(n2573), .ZN(N195)
         );
  AOI221_X1 U2231 ( .B1(n166), .B2(\registers[13][10] ), .C1(n163), .C2(
        \registers[12][10] ), .A(n2585), .ZN(n2571) );
  AOI221_X1 U2232 ( .B1(n26), .B2(\registers[9][10] ), .C1(n23), .C2(
        \registers[8][10] ), .A(n2586), .ZN(n2570) );
  AOI211_X1 U2233 ( .C1(n187), .C2(\registers[1][10] ), .A(n2582), .B(n2583), 
        .ZN(n2572) );
  NAND4_X1 U2234 ( .A1(n2553), .A2(n2554), .A3(n2555), .A4(n2556), .ZN(N196)
         );
  AOI221_X1 U2235 ( .B1(n167), .B2(\registers[13][11] ), .C1(n164), .C2(
        \registers[12][11] ), .A(n2568), .ZN(n2554) );
  AOI221_X1 U2236 ( .B1(n27), .B2(\registers[9][11] ), .C1(n24), .C2(
        \registers[8][11] ), .A(n2569), .ZN(n2553) );
  AOI211_X1 U2237 ( .C1(n188), .C2(\registers[1][11] ), .A(n2565), .B(n2566), 
        .ZN(n2555) );
  NAND4_X1 U2238 ( .A1(n2536), .A2(n2537), .A3(n2538), .A4(n2539), .ZN(N197)
         );
  AOI221_X1 U2239 ( .B1(n167), .B2(\registers[13][12] ), .C1(n164), .C2(
        \registers[12][12] ), .A(n2551), .ZN(n2537) );
  AOI221_X1 U2240 ( .B1(n27), .B2(\registers[9][12] ), .C1(n24), .C2(
        \registers[8][12] ), .A(n2552), .ZN(n2536) );
  AOI211_X1 U2241 ( .C1(n188), .C2(\registers[1][12] ), .A(n2548), .B(n2549), 
        .ZN(n2538) );
  NAND4_X1 U2242 ( .A1(n2519), .A2(n2520), .A3(n2521), .A4(n2522), .ZN(N198)
         );
  AOI221_X1 U2243 ( .B1(n167), .B2(\registers[13][13] ), .C1(n164), .C2(
        \registers[12][13] ), .A(n2534), .ZN(n2520) );
  AOI221_X1 U2244 ( .B1(n27), .B2(\registers[9][13] ), .C1(n24), .C2(
        \registers[8][13] ), .A(n2535), .ZN(n2519) );
  AOI211_X1 U2245 ( .C1(n188), .C2(\registers[1][13] ), .A(n2531), .B(n2532), 
        .ZN(n2521) );
  NAND4_X1 U2246 ( .A1(n2502), .A2(n2503), .A3(n2504), .A4(n2505), .ZN(N199)
         );
  AOI221_X1 U2247 ( .B1(n167), .B2(\registers[13][14] ), .C1(n164), .C2(
        \registers[12][14] ), .A(n2517), .ZN(n2503) );
  AOI221_X1 U2248 ( .B1(n27), .B2(\registers[9][14] ), .C1(n24), .C2(
        \registers[8][14] ), .A(n2518), .ZN(n2502) );
  AOI211_X1 U2249 ( .C1(n188), .C2(\registers[1][14] ), .A(n2514), .B(n2515), 
        .ZN(n2504) );
  NAND4_X1 U2250 ( .A1(n2485), .A2(n2486), .A3(n2487), .A4(n2488), .ZN(N200)
         );
  AOI221_X1 U2251 ( .B1(n167), .B2(\registers[13][15] ), .C1(n164), .C2(
        \registers[12][15] ), .A(n2500), .ZN(n2486) );
  AOI221_X1 U2252 ( .B1(n27), .B2(\registers[9][15] ), .C1(n24), .C2(
        \registers[8][15] ), .A(n2501), .ZN(n2485) );
  AOI211_X1 U2253 ( .C1(n188), .C2(\registers[1][15] ), .A(n2497), .B(n2498), 
        .ZN(n2487) );
  NAND4_X1 U2254 ( .A1(n2468), .A2(n2469), .A3(n2470), .A4(n2471), .ZN(N201)
         );
  AOI221_X1 U2255 ( .B1(n167), .B2(\registers[13][16] ), .C1(n164), .C2(
        \registers[12][16] ), .A(n2483), .ZN(n2469) );
  AOI221_X1 U2256 ( .B1(n27), .B2(\registers[9][16] ), .C1(n24), .C2(
        \registers[8][16] ), .A(n2484), .ZN(n2468) );
  AOI211_X1 U2257 ( .C1(n188), .C2(\registers[1][16] ), .A(n2480), .B(n2481), 
        .ZN(n2470) );
  NAND4_X1 U2258 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(N202)
         );
  AOI221_X1 U2259 ( .B1(n167), .B2(\registers[13][17] ), .C1(n164), .C2(
        \registers[12][17] ), .A(n2466), .ZN(n2452) );
  AOI221_X1 U2260 ( .B1(n27), .B2(\registers[9][17] ), .C1(n24), .C2(
        \registers[8][17] ), .A(n2467), .ZN(n2451) );
  AOI211_X1 U2261 ( .C1(n188), .C2(\registers[1][17] ), .A(n2463), .B(n2464), 
        .ZN(n2453) );
  NAND4_X1 U2262 ( .A1(n2434), .A2(n2435), .A3(n2436), .A4(n2437), .ZN(N203)
         );
  AOI221_X1 U2263 ( .B1(n167), .B2(\registers[13][18] ), .C1(n164), .C2(
        \registers[12][18] ), .A(n2449), .ZN(n2435) );
  AOI221_X1 U2264 ( .B1(n27), .B2(\registers[9][18] ), .C1(n24), .C2(
        \registers[8][18] ), .A(n2450), .ZN(n2434) );
  AOI211_X1 U2265 ( .C1(n188), .C2(\registers[1][18] ), .A(n2446), .B(n2447), 
        .ZN(n2436) );
  NAND4_X1 U2266 ( .A1(n2417), .A2(n2418), .A3(n2419), .A4(n2420), .ZN(N204)
         );
  AOI221_X1 U2267 ( .B1(n167), .B2(\registers[13][19] ), .C1(n164), .C2(
        \registers[12][19] ), .A(n2432), .ZN(n2418) );
  AOI221_X1 U2268 ( .B1(n27), .B2(\registers[9][19] ), .C1(n24), .C2(
        \registers[8][19] ), .A(n2433), .ZN(n2417) );
  AOI211_X1 U2269 ( .C1(n188), .C2(\registers[1][19] ), .A(n2429), .B(n2430), 
        .ZN(n2419) );
  NAND4_X1 U2270 ( .A1(n2400), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(N205)
         );
  AOI221_X1 U2271 ( .B1(n167), .B2(\registers[13][20] ), .C1(n164), .C2(
        \registers[12][20] ), .A(n2415), .ZN(n2401) );
  AOI221_X1 U2272 ( .B1(n27), .B2(\registers[9][20] ), .C1(n24), .C2(
        \registers[8][20] ), .A(n2416), .ZN(n2400) );
  AOI211_X1 U2273 ( .C1(n188), .C2(\registers[1][20] ), .A(n2412), .B(n2413), 
        .ZN(n2402) );
  NAND4_X1 U2274 ( .A1(n2383), .A2(n2384), .A3(n2385), .A4(n2386), .ZN(N206)
         );
  AOI221_X1 U2275 ( .B1(n167), .B2(\registers[13][21] ), .C1(n164), .C2(
        \registers[12][21] ), .A(n2398), .ZN(n2384) );
  AOI221_X1 U2276 ( .B1(n27), .B2(\registers[9][21] ), .C1(n24), .C2(
        \registers[8][21] ), .A(n2399), .ZN(n2383) );
  AOI211_X1 U2277 ( .C1(n188), .C2(\registers[1][21] ), .A(n2395), .B(n2396), 
        .ZN(n2385) );
  NAND4_X1 U2278 ( .A1(n2366), .A2(n2367), .A3(n2368), .A4(n2369), .ZN(N207)
         );
  AOI221_X1 U2279 ( .B1(n168), .B2(\registers[13][22] ), .C1(n165), .C2(
        \registers[12][22] ), .A(n2381), .ZN(n2367) );
  AOI221_X1 U2280 ( .B1(n28), .B2(\registers[9][22] ), .C1(n25), .C2(
        \registers[8][22] ), .A(n2382), .ZN(n2366) );
  AOI211_X1 U2281 ( .C1(n189), .C2(\registers[1][22] ), .A(n2378), .B(n2379), 
        .ZN(n2368) );
  NAND4_X1 U2282 ( .A1(n2349), .A2(n2350), .A3(n2351), .A4(n2352), .ZN(N208)
         );
  AOI221_X1 U2283 ( .B1(n168), .B2(\registers[13][23] ), .C1(n165), .C2(
        \registers[12][23] ), .A(n2364), .ZN(n2350) );
  AOI221_X1 U2284 ( .B1(n28), .B2(\registers[9][23] ), .C1(n25), .C2(
        \registers[8][23] ), .A(n2365), .ZN(n2349) );
  AOI211_X1 U2285 ( .C1(n189), .C2(\registers[1][23] ), .A(n2361), .B(n2362), 
        .ZN(n2351) );
  NAND4_X1 U2286 ( .A1(n2332), .A2(n2333), .A3(n2334), .A4(n2335), .ZN(N209)
         );
  AOI221_X1 U2287 ( .B1(n168), .B2(\registers[13][24] ), .C1(n165), .C2(
        \registers[12][24] ), .A(n2347), .ZN(n2333) );
  AOI221_X1 U2288 ( .B1(n28), .B2(\registers[9][24] ), .C1(n25), .C2(
        \registers[8][24] ), .A(n2348), .ZN(n2332) );
  AOI211_X1 U2289 ( .C1(n189), .C2(\registers[1][24] ), .A(n2344), .B(n2345), 
        .ZN(n2334) );
  NAND4_X1 U2290 ( .A1(n2315), .A2(n2316), .A3(n2317), .A4(n2318), .ZN(N210)
         );
  AOI221_X1 U2291 ( .B1(n168), .B2(\registers[13][25] ), .C1(n165), .C2(
        \registers[12][25] ), .A(n2330), .ZN(n2316) );
  AOI221_X1 U2292 ( .B1(n28), .B2(\registers[9][25] ), .C1(n25), .C2(
        \registers[8][25] ), .A(n2331), .ZN(n2315) );
  AOI211_X1 U2293 ( .C1(n189), .C2(\registers[1][25] ), .A(n2327), .B(n2328), 
        .ZN(n2317) );
  NAND4_X1 U2294 ( .A1(n2298), .A2(n2299), .A3(n2300), .A4(n2301), .ZN(N211)
         );
  AOI221_X1 U2295 ( .B1(n168), .B2(\registers[13][26] ), .C1(n165), .C2(
        \registers[12][26] ), .A(n2313), .ZN(n2299) );
  AOI221_X1 U2296 ( .B1(n28), .B2(\registers[9][26] ), .C1(n25), .C2(
        \registers[8][26] ), .A(n2314), .ZN(n2298) );
  AOI211_X1 U2297 ( .C1(n189), .C2(\registers[1][26] ), .A(n2310), .B(n2311), 
        .ZN(n2300) );
  NAND4_X1 U2298 ( .A1(n2281), .A2(n2282), .A3(n2283), .A4(n2284), .ZN(N212)
         );
  AOI221_X1 U2299 ( .B1(n168), .B2(\registers[13][27] ), .C1(n165), .C2(
        \registers[12][27] ), .A(n2296), .ZN(n2282) );
  AOI221_X1 U2300 ( .B1(n28), .B2(\registers[9][27] ), .C1(n25), .C2(
        \registers[8][27] ), .A(n2297), .ZN(n2281) );
  AOI211_X1 U2301 ( .C1(n189), .C2(\registers[1][27] ), .A(n2293), .B(n2294), 
        .ZN(n2283) );
  NAND4_X1 U2302 ( .A1(n2264), .A2(n2265), .A3(n2266), .A4(n2267), .ZN(N213)
         );
  AOI221_X1 U2303 ( .B1(n168), .B2(\registers[13][28] ), .C1(n165), .C2(
        \registers[12][28] ), .A(n2279), .ZN(n2265) );
  AOI221_X1 U2304 ( .B1(n28), .B2(\registers[9][28] ), .C1(n25), .C2(
        \registers[8][28] ), .A(n2280), .ZN(n2264) );
  AOI211_X1 U2305 ( .C1(n189), .C2(\registers[1][28] ), .A(n2276), .B(n2277), 
        .ZN(n2266) );
  NAND4_X1 U2306 ( .A1(n2247), .A2(n2248), .A3(n2249), .A4(n2250), .ZN(N214)
         );
  AOI221_X1 U2307 ( .B1(n168), .B2(\registers[13][29] ), .C1(n165), .C2(
        \registers[12][29] ), .A(n2262), .ZN(n2248) );
  AOI221_X1 U2308 ( .B1(n28), .B2(\registers[9][29] ), .C1(n25), .C2(
        \registers[8][29] ), .A(n2263), .ZN(n2247) );
  AOI211_X1 U2309 ( .C1(n189), .C2(\registers[1][29] ), .A(n2259), .B(n2260), 
        .ZN(n2249) );
  NAND4_X1 U2310 ( .A1(n2230), .A2(n2231), .A3(n2232), .A4(n2233), .ZN(N215)
         );
  AOI221_X1 U2311 ( .B1(n168), .B2(\registers[13][30] ), .C1(n165), .C2(
        \registers[12][30] ), .A(n2245), .ZN(n2231) );
  AOI221_X1 U2312 ( .B1(n28), .B2(\registers[9][30] ), .C1(n25), .C2(
        \registers[8][30] ), .A(n2246), .ZN(n2230) );
  AOI211_X1 U2313 ( .C1(n189), .C2(\registers[1][30] ), .A(n2242), .B(n2243), 
        .ZN(n2232) );
  NAND4_X1 U2314 ( .A1(n2182), .A2(n2183), .A3(n2184), .A4(n2185), .ZN(N216)
         );
  AOI221_X1 U2315 ( .B1(n168), .B2(\registers[13][31] ), .C1(n165), .C2(
        \registers[12][31] ), .A(n2222), .ZN(n2183) );
  AOI221_X1 U2316 ( .B1(n28), .B2(\registers[9][31] ), .C1(n25), .C2(
        \registers[8][31] ), .A(n2227), .ZN(n2182) );
  AOI211_X1 U2317 ( .C1(n189), .C2(\registers[1][31] ), .A(n2211), .B(n2212), 
        .ZN(n2184) );
  NOR2_X1 U2318 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n2176) );
  NOR2_X1 U2319 ( .A1(n3810), .A2(ADD_RD2[4]), .ZN(n2181) );
  NOR2_X1 U2320 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n2767) );
  NOR2_X1 U2321 ( .A1(n3807), .A2(ADD_RD1[4]), .ZN(n2772) );
  AND2_X1 U2322 ( .A1(n2165), .A2(ADD_RD2[0]), .ZN(n2160) );
  AND2_X1 U2323 ( .A1(n2176), .A2(ADD_RD2[0]), .ZN(n2173) );
  AND2_X1 U2324 ( .A1(n2181), .A2(ADD_RD2[0]), .ZN(n2178) );
  AND2_X1 U2325 ( .A1(n2756), .A2(ADD_RD1[0]), .ZN(n2751) );
  AND2_X1 U2326 ( .A1(n2767), .A2(ADD_RD1[0]), .ZN(n2764) );
  AND2_X1 U2327 ( .A1(n2772), .A2(ADD_RD1[0]), .ZN(n2769) );
  INV_X1 U2328 ( .A(ADD_RD2[0]), .ZN(n3812) );
  INV_X1 U2329 ( .A(ADD_RD1[0]), .ZN(n3809) );
  AND2_X1 U2330 ( .A1(WR), .A2(ENABLE), .ZN(n1293) );
  INV_X1 U2331 ( .A(ADD_RD2[3]), .ZN(n3810) );
  INV_X1 U2332 ( .A(ADD_RD2[1]), .ZN(n3811) );
  INV_X1 U2333 ( .A(ADD_RD1[3]), .ZN(n3807) );
  INV_X1 U2334 ( .A(ADD_RD1[1]), .ZN(n3808) );
  AND2_X1 U2335 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n2170) );
  AND2_X1 U2336 ( .A1(ADD_RD2[4]), .A2(n3810), .ZN(n2165) );
  AND2_X1 U2337 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2761) );
  AND2_X1 U2338 ( .A1(ADD_RD1[4]), .A2(n3807), .ZN(n2756) );
  INV_X1 U2339 ( .A(n1159), .ZN(n3771) );
  AOI22_X1 U2340 ( .A1(DATAIN[0]), .A2(n777), .B1(n778), .B2(
        \registers[29][0] ), .ZN(n1159) );
  INV_X1 U2341 ( .A(n1161), .ZN(n3772) );
  AOI22_X1 U2342 ( .A1(DATAIN[1]), .A2(n776), .B1(n778), .B2(
        \registers[29][1] ), .ZN(n1161) );
  INV_X1 U2343 ( .A(n1162), .ZN(n3773) );
  AOI22_X1 U2344 ( .A1(DATAIN[2]), .A2(n777), .B1(n778), .B2(
        \registers[29][2] ), .ZN(n1162) );
  INV_X1 U2345 ( .A(n1163), .ZN(n3774) );
  AOI22_X1 U2346 ( .A1(DATAIN[3]), .A2(n776), .B1(n778), .B2(
        \registers[29][3] ), .ZN(n1163) );
  INV_X1 U2347 ( .A(n1164), .ZN(n3775) );
  AOI22_X1 U2348 ( .A1(DATAIN[4]), .A2(n777), .B1(n778), .B2(
        \registers[29][4] ), .ZN(n1164) );
  INV_X1 U2349 ( .A(n1165), .ZN(n3776) );
  AOI22_X1 U2350 ( .A1(DATAIN[5]), .A2(n776), .B1(n779), .B2(
        \registers[29][5] ), .ZN(n1165) );
  INV_X1 U2351 ( .A(n1166), .ZN(n3777) );
  AOI22_X1 U2352 ( .A1(DATAIN[6]), .A2(n777), .B1(n779), .B2(
        \registers[29][6] ), .ZN(n1166) );
  INV_X1 U2353 ( .A(n1167), .ZN(n3778) );
  AOI22_X1 U2354 ( .A1(DATAIN[7]), .A2(n776), .B1(n779), .B2(
        \registers[29][7] ), .ZN(n1167) );
  INV_X1 U2355 ( .A(n1168), .ZN(n3779) );
  AOI22_X1 U2356 ( .A1(DATAIN[8]), .A2(n777), .B1(n779), .B2(
        \registers[29][8] ), .ZN(n1168) );
  INV_X1 U2357 ( .A(n1169), .ZN(n3780) );
  AOI22_X1 U2358 ( .A1(DATAIN[9]), .A2(n777), .B1(n779), .B2(
        \registers[29][9] ), .ZN(n1169) );
  INV_X1 U2359 ( .A(n1170), .ZN(n3781) );
  AOI22_X1 U2360 ( .A1(DATAIN[10]), .A2(n777), .B1(n780), .B2(
        \registers[29][10] ), .ZN(n1170) );
  INV_X1 U2361 ( .A(n1171), .ZN(n3782) );
  AOI22_X1 U2362 ( .A1(DATAIN[11]), .A2(n777), .B1(n780), .B2(
        \registers[29][11] ), .ZN(n1171) );
  INV_X1 U2363 ( .A(n1172), .ZN(n3783) );
  AOI22_X1 U2364 ( .A1(DATAIN[12]), .A2(n777), .B1(n780), .B2(
        \registers[29][12] ), .ZN(n1172) );
  INV_X1 U2365 ( .A(n1173), .ZN(n3784) );
  AOI22_X1 U2366 ( .A1(DATAIN[13]), .A2(n777), .B1(n780), .B2(
        \registers[29][13] ), .ZN(n1173) );
  INV_X1 U2367 ( .A(n1174), .ZN(n3785) );
  AOI22_X1 U2368 ( .A1(DATAIN[14]), .A2(n777), .B1(n780), .B2(
        \registers[29][14] ), .ZN(n1174) );
  INV_X1 U2369 ( .A(n1175), .ZN(n3786) );
  AOI22_X1 U2370 ( .A1(DATAIN[15]), .A2(n777), .B1(n781), .B2(
        \registers[29][15] ), .ZN(n1175) );
  INV_X1 U2371 ( .A(n1176), .ZN(n3787) );
  AOI22_X1 U2372 ( .A1(DATAIN[16]), .A2(n777), .B1(n781), .B2(
        \registers[29][16] ), .ZN(n1176) );
  INV_X1 U2373 ( .A(n1177), .ZN(n3788) );
  AOI22_X1 U2374 ( .A1(DATAIN[17]), .A2(n777), .B1(n781), .B2(
        \registers[29][17] ), .ZN(n1177) );
  INV_X1 U2375 ( .A(n1178), .ZN(n3789) );
  AOI22_X1 U2376 ( .A1(DATAIN[18]), .A2(n777), .B1(n781), .B2(
        \registers[29][18] ), .ZN(n1178) );
  INV_X1 U2377 ( .A(n1179), .ZN(n3790) );
  AOI22_X1 U2378 ( .A1(DATAIN[19]), .A2(n777), .B1(n781), .B2(
        \registers[29][19] ), .ZN(n1179) );
  INV_X1 U2379 ( .A(n1180), .ZN(n3791) );
  AOI22_X1 U2380 ( .A1(DATAIN[20]), .A2(n776), .B1(n782), .B2(
        \registers[29][20] ), .ZN(n1180) );
  INV_X1 U2381 ( .A(n1181), .ZN(n3792) );
  AOI22_X1 U2382 ( .A1(DATAIN[21]), .A2(n776), .B1(n782), .B2(
        \registers[29][21] ), .ZN(n1181) );
  INV_X1 U2383 ( .A(n1182), .ZN(n3793) );
  AOI22_X1 U2384 ( .A1(DATAIN[22]), .A2(n776), .B1(n782), .B2(
        \registers[29][22] ), .ZN(n1182) );
  INV_X1 U2385 ( .A(n1192), .ZN(n3739) );
  AOI22_X1 U2386 ( .A1(DATAIN[0]), .A2(n768), .B1(n769), .B2(
        \registers[28][0] ), .ZN(n1192) );
  INV_X1 U2387 ( .A(n1194), .ZN(n3740) );
  AOI22_X1 U2388 ( .A1(DATAIN[1]), .A2(n767), .B1(n769), .B2(
        \registers[28][1] ), .ZN(n1194) );
  INV_X1 U2389 ( .A(n1195), .ZN(n3741) );
  AOI22_X1 U2390 ( .A1(DATAIN[2]), .A2(n768), .B1(n769), .B2(
        \registers[28][2] ), .ZN(n1195) );
  INV_X1 U2391 ( .A(n1196), .ZN(n3742) );
  AOI22_X1 U2392 ( .A1(DATAIN[3]), .A2(n767), .B1(n769), .B2(
        \registers[28][3] ), .ZN(n1196) );
  INV_X1 U2393 ( .A(n1197), .ZN(n3743) );
  AOI22_X1 U2394 ( .A1(DATAIN[4]), .A2(n768), .B1(n769), .B2(
        \registers[28][4] ), .ZN(n1197) );
  INV_X1 U2395 ( .A(n1198), .ZN(n3744) );
  AOI22_X1 U2396 ( .A1(DATAIN[5]), .A2(n767), .B1(n770), .B2(
        \registers[28][5] ), .ZN(n1198) );
  INV_X1 U2397 ( .A(n1199), .ZN(n3745) );
  AOI22_X1 U2398 ( .A1(DATAIN[6]), .A2(n768), .B1(n770), .B2(
        \registers[28][6] ), .ZN(n1199) );
  INV_X1 U2399 ( .A(n1200), .ZN(n3746) );
  AOI22_X1 U2400 ( .A1(DATAIN[7]), .A2(n767), .B1(n770), .B2(
        \registers[28][7] ), .ZN(n1200) );
  INV_X1 U2401 ( .A(n1201), .ZN(n3747) );
  AOI22_X1 U2402 ( .A1(DATAIN[8]), .A2(n768), .B1(n770), .B2(
        \registers[28][8] ), .ZN(n1201) );
  INV_X1 U2403 ( .A(n1202), .ZN(n3748) );
  AOI22_X1 U2404 ( .A1(DATAIN[9]), .A2(n768), .B1(n770), .B2(
        \registers[28][9] ), .ZN(n1202) );
  INV_X1 U2405 ( .A(n1203), .ZN(n3749) );
  AOI22_X1 U2406 ( .A1(DATAIN[10]), .A2(n768), .B1(n771), .B2(
        \registers[28][10] ), .ZN(n1203) );
  INV_X1 U2407 ( .A(n1204), .ZN(n3750) );
  AOI22_X1 U2408 ( .A1(DATAIN[11]), .A2(n768), .B1(n771), .B2(
        \registers[28][11] ), .ZN(n1204) );
  INV_X1 U2409 ( .A(n1205), .ZN(n3751) );
  AOI22_X1 U2410 ( .A1(DATAIN[12]), .A2(n768), .B1(n771), .B2(
        \registers[28][12] ), .ZN(n1205) );
  INV_X1 U2411 ( .A(n1206), .ZN(n3752) );
  AOI22_X1 U2412 ( .A1(DATAIN[13]), .A2(n768), .B1(n771), .B2(
        \registers[28][13] ), .ZN(n1206) );
  INV_X1 U2413 ( .A(n1207), .ZN(n3753) );
  AOI22_X1 U2414 ( .A1(DATAIN[14]), .A2(n768), .B1(n771), .B2(
        \registers[28][14] ), .ZN(n1207) );
  INV_X1 U2415 ( .A(n1208), .ZN(n3754) );
  AOI22_X1 U2416 ( .A1(DATAIN[15]), .A2(n768), .B1(n772), .B2(
        \registers[28][15] ), .ZN(n1208) );
  INV_X1 U2417 ( .A(n1209), .ZN(n3755) );
  AOI22_X1 U2418 ( .A1(DATAIN[16]), .A2(n768), .B1(n772), .B2(
        \registers[28][16] ), .ZN(n1209) );
  INV_X1 U2419 ( .A(n1210), .ZN(n3756) );
  AOI22_X1 U2420 ( .A1(DATAIN[17]), .A2(n768), .B1(n772), .B2(
        \registers[28][17] ), .ZN(n1210) );
  INV_X1 U2421 ( .A(n1211), .ZN(n3757) );
  AOI22_X1 U2422 ( .A1(DATAIN[18]), .A2(n768), .B1(n772), .B2(
        \registers[28][18] ), .ZN(n1211) );
  INV_X1 U2423 ( .A(n1212), .ZN(n3758) );
  AOI22_X1 U2424 ( .A1(DATAIN[19]), .A2(n768), .B1(n772), .B2(
        \registers[28][19] ), .ZN(n1212) );
  INV_X1 U2425 ( .A(n1213), .ZN(n3759) );
  AOI22_X1 U2426 ( .A1(DATAIN[20]), .A2(n767), .B1(n773), .B2(
        \registers[28][20] ), .ZN(n1213) );
  INV_X1 U2427 ( .A(n1214), .ZN(n3760) );
  AOI22_X1 U2428 ( .A1(DATAIN[21]), .A2(n767), .B1(n773), .B2(
        \registers[28][21] ), .ZN(n1214) );
  INV_X1 U2429 ( .A(n1215), .ZN(n3761) );
  AOI22_X1 U2430 ( .A1(DATAIN[22]), .A2(n767), .B1(n773), .B2(
        \registers[28][22] ), .ZN(n1215) );
  INV_X1 U2431 ( .A(n1227), .ZN(n3707) );
  AOI22_X1 U2432 ( .A1(DATAIN[0]), .A2(n741), .B1(n742), .B2(
        \registers[25][0] ), .ZN(n1227) );
  INV_X1 U2433 ( .A(n1229), .ZN(n3708) );
  AOI22_X1 U2434 ( .A1(DATAIN[1]), .A2(n740), .B1(n742), .B2(
        \registers[25][1] ), .ZN(n1229) );
  INV_X1 U2435 ( .A(n1230), .ZN(n3709) );
  AOI22_X1 U2436 ( .A1(DATAIN[2]), .A2(n741), .B1(n742), .B2(
        \registers[25][2] ), .ZN(n1230) );
  INV_X1 U2437 ( .A(n1231), .ZN(n3710) );
  AOI22_X1 U2438 ( .A1(DATAIN[3]), .A2(n740), .B1(n742), .B2(
        \registers[25][3] ), .ZN(n1231) );
  INV_X1 U2439 ( .A(n1232), .ZN(n3711) );
  AOI22_X1 U2440 ( .A1(DATAIN[4]), .A2(n741), .B1(n742), .B2(
        \registers[25][4] ), .ZN(n1232) );
  INV_X1 U2441 ( .A(n1233), .ZN(n3712) );
  AOI22_X1 U2442 ( .A1(DATAIN[5]), .A2(n740), .B1(n743), .B2(
        \registers[25][5] ), .ZN(n1233) );
  INV_X1 U2443 ( .A(n1234), .ZN(n3713) );
  AOI22_X1 U2444 ( .A1(DATAIN[6]), .A2(n741), .B1(n743), .B2(
        \registers[25][6] ), .ZN(n1234) );
  INV_X1 U2445 ( .A(n1235), .ZN(n3714) );
  AOI22_X1 U2446 ( .A1(DATAIN[7]), .A2(n740), .B1(n743), .B2(
        \registers[25][7] ), .ZN(n1235) );
  INV_X1 U2447 ( .A(n1236), .ZN(n3715) );
  AOI22_X1 U2448 ( .A1(DATAIN[8]), .A2(n741), .B1(n743), .B2(
        \registers[25][8] ), .ZN(n1236) );
  INV_X1 U2449 ( .A(n1237), .ZN(n3716) );
  AOI22_X1 U2450 ( .A1(DATAIN[9]), .A2(n741), .B1(n743), .B2(
        \registers[25][9] ), .ZN(n1237) );
  INV_X1 U2451 ( .A(n1238), .ZN(n3717) );
  AOI22_X1 U2452 ( .A1(DATAIN[10]), .A2(n741), .B1(n744), .B2(
        \registers[25][10] ), .ZN(n1238) );
  INV_X1 U2453 ( .A(n1239), .ZN(n3718) );
  AOI22_X1 U2454 ( .A1(DATAIN[11]), .A2(n741), .B1(n744), .B2(
        \registers[25][11] ), .ZN(n1239) );
  INV_X1 U2455 ( .A(n1240), .ZN(n3719) );
  AOI22_X1 U2456 ( .A1(DATAIN[12]), .A2(n741), .B1(n744), .B2(
        \registers[25][12] ), .ZN(n1240) );
  INV_X1 U2457 ( .A(n1241), .ZN(n3720) );
  AOI22_X1 U2458 ( .A1(DATAIN[13]), .A2(n741), .B1(n744), .B2(
        \registers[25][13] ), .ZN(n1241) );
  INV_X1 U2459 ( .A(n1242), .ZN(n3721) );
  AOI22_X1 U2460 ( .A1(DATAIN[14]), .A2(n741), .B1(n744), .B2(
        \registers[25][14] ), .ZN(n1242) );
  INV_X1 U2461 ( .A(n1243), .ZN(n3722) );
  AOI22_X1 U2462 ( .A1(DATAIN[15]), .A2(n741), .B1(n745), .B2(
        \registers[25][15] ), .ZN(n1243) );
  INV_X1 U2463 ( .A(n1244), .ZN(n3723) );
  AOI22_X1 U2464 ( .A1(DATAIN[16]), .A2(n741), .B1(n745), .B2(
        \registers[25][16] ), .ZN(n1244) );
  INV_X1 U2465 ( .A(n1245), .ZN(n3724) );
  AOI22_X1 U2466 ( .A1(DATAIN[17]), .A2(n741), .B1(n745), .B2(
        \registers[25][17] ), .ZN(n1245) );
  INV_X1 U2467 ( .A(n1246), .ZN(n3725) );
  AOI22_X1 U2468 ( .A1(DATAIN[18]), .A2(n741), .B1(n745), .B2(
        \registers[25][18] ), .ZN(n1246) );
  INV_X1 U2469 ( .A(n1247), .ZN(n3726) );
  AOI22_X1 U2470 ( .A1(DATAIN[19]), .A2(n741), .B1(n745), .B2(
        \registers[25][19] ), .ZN(n1247) );
  INV_X1 U2471 ( .A(n1248), .ZN(n3727) );
  AOI22_X1 U2472 ( .A1(DATAIN[20]), .A2(n740), .B1(n746), .B2(
        \registers[25][20] ), .ZN(n1248) );
  INV_X1 U2473 ( .A(n1249), .ZN(n3728) );
  AOI22_X1 U2474 ( .A1(DATAIN[21]), .A2(n740), .B1(n746), .B2(
        \registers[25][21] ), .ZN(n1249) );
  INV_X1 U2475 ( .A(n1250), .ZN(n3729) );
  AOI22_X1 U2476 ( .A1(DATAIN[22]), .A2(n740), .B1(n746), .B2(
        \registers[25][22] ), .ZN(n1250) );
  INV_X1 U2477 ( .A(n1260), .ZN(n3675) );
  AOI22_X1 U2478 ( .A1(DATAIN[0]), .A2(n732), .B1(n733), .B2(
        \registers[24][0] ), .ZN(n1260) );
  INV_X1 U2479 ( .A(n1262), .ZN(n3676) );
  AOI22_X1 U2480 ( .A1(DATAIN[1]), .A2(n731), .B1(n733), .B2(
        \registers[24][1] ), .ZN(n1262) );
  INV_X1 U2481 ( .A(n1263), .ZN(n3677) );
  AOI22_X1 U2482 ( .A1(DATAIN[2]), .A2(n732), .B1(n733), .B2(
        \registers[24][2] ), .ZN(n1263) );
  INV_X1 U2483 ( .A(n1264), .ZN(n3678) );
  AOI22_X1 U2484 ( .A1(DATAIN[3]), .A2(n731), .B1(n733), .B2(
        \registers[24][3] ), .ZN(n1264) );
  INV_X1 U2485 ( .A(n1265), .ZN(n3679) );
  AOI22_X1 U2486 ( .A1(DATAIN[4]), .A2(n732), .B1(n733), .B2(
        \registers[24][4] ), .ZN(n1265) );
  INV_X1 U2487 ( .A(n1266), .ZN(n3680) );
  AOI22_X1 U2488 ( .A1(DATAIN[5]), .A2(n731), .B1(n734), .B2(
        \registers[24][5] ), .ZN(n1266) );
  INV_X1 U2489 ( .A(n1267), .ZN(n3681) );
  AOI22_X1 U2490 ( .A1(DATAIN[6]), .A2(n732), .B1(n734), .B2(
        \registers[24][6] ), .ZN(n1267) );
  INV_X1 U2491 ( .A(n1268), .ZN(n3682) );
  AOI22_X1 U2492 ( .A1(DATAIN[7]), .A2(n731), .B1(n734), .B2(
        \registers[24][7] ), .ZN(n1268) );
  INV_X1 U2493 ( .A(n1269), .ZN(n3683) );
  AOI22_X1 U2494 ( .A1(DATAIN[8]), .A2(n732), .B1(n734), .B2(
        \registers[24][8] ), .ZN(n1269) );
  INV_X1 U2495 ( .A(n1270), .ZN(n3684) );
  AOI22_X1 U2496 ( .A1(DATAIN[9]), .A2(n732), .B1(n734), .B2(
        \registers[24][9] ), .ZN(n1270) );
  INV_X1 U2497 ( .A(n1271), .ZN(n3685) );
  AOI22_X1 U2498 ( .A1(DATAIN[10]), .A2(n732), .B1(n735), .B2(
        \registers[24][10] ), .ZN(n1271) );
  INV_X1 U2499 ( .A(n1272), .ZN(n3686) );
  AOI22_X1 U2500 ( .A1(DATAIN[11]), .A2(n732), .B1(n735), .B2(
        \registers[24][11] ), .ZN(n1272) );
  INV_X1 U2501 ( .A(n1273), .ZN(n3687) );
  AOI22_X1 U2502 ( .A1(DATAIN[12]), .A2(n732), .B1(n735), .B2(
        \registers[24][12] ), .ZN(n1273) );
  INV_X1 U2503 ( .A(n1274), .ZN(n3688) );
  AOI22_X1 U2504 ( .A1(DATAIN[13]), .A2(n732), .B1(n735), .B2(
        \registers[24][13] ), .ZN(n1274) );
  INV_X1 U2505 ( .A(n1275), .ZN(n3689) );
  AOI22_X1 U2506 ( .A1(DATAIN[14]), .A2(n732), .B1(n735), .B2(
        \registers[24][14] ), .ZN(n1275) );
  INV_X1 U2507 ( .A(n1276), .ZN(n3690) );
  AOI22_X1 U2508 ( .A1(DATAIN[15]), .A2(n732), .B1(n736), .B2(
        \registers[24][15] ), .ZN(n1276) );
  INV_X1 U2509 ( .A(n1277), .ZN(n3691) );
  AOI22_X1 U2510 ( .A1(DATAIN[16]), .A2(n732), .B1(n736), .B2(
        \registers[24][16] ), .ZN(n1277) );
  INV_X1 U2511 ( .A(n1278), .ZN(n3692) );
  AOI22_X1 U2512 ( .A1(DATAIN[17]), .A2(n732), .B1(n736), .B2(
        \registers[24][17] ), .ZN(n1278) );
  INV_X1 U2513 ( .A(n1279), .ZN(n3693) );
  AOI22_X1 U2514 ( .A1(DATAIN[18]), .A2(n732), .B1(n736), .B2(
        \registers[24][18] ), .ZN(n1279) );
  INV_X1 U2515 ( .A(n1280), .ZN(n3694) );
  AOI22_X1 U2516 ( .A1(DATAIN[19]), .A2(n732), .B1(n736), .B2(
        \registers[24][19] ), .ZN(n1280) );
  INV_X1 U2517 ( .A(n1281), .ZN(n3695) );
  AOI22_X1 U2518 ( .A1(DATAIN[20]), .A2(n731), .B1(n737), .B2(
        \registers[24][20] ), .ZN(n1281) );
  INV_X1 U2519 ( .A(n1282), .ZN(n3696) );
  AOI22_X1 U2520 ( .A1(DATAIN[21]), .A2(n731), .B1(n737), .B2(
        \registers[24][21] ), .ZN(n1282) );
  INV_X1 U2521 ( .A(n1283), .ZN(n3697) );
  AOI22_X1 U2522 ( .A1(DATAIN[22]), .A2(n731), .B1(n737), .B2(
        \registers[24][22] ), .ZN(n1283) );
  INV_X1 U2523 ( .A(n1294), .ZN(n3643) );
  AOI22_X1 U2524 ( .A1(DATAIN[0]), .A2(n723), .B1(n724), .B2(
        \registers[23][0] ), .ZN(n1294) );
  INV_X1 U2525 ( .A(n1296), .ZN(n3644) );
  AOI22_X1 U2526 ( .A1(DATAIN[1]), .A2(n722), .B1(n724), .B2(
        \registers[23][1] ), .ZN(n1296) );
  INV_X1 U2527 ( .A(n1297), .ZN(n3645) );
  AOI22_X1 U2528 ( .A1(DATAIN[2]), .A2(n723), .B1(n724), .B2(
        \registers[23][2] ), .ZN(n1297) );
  INV_X1 U2529 ( .A(n1298), .ZN(n3646) );
  AOI22_X1 U2530 ( .A1(DATAIN[3]), .A2(n722), .B1(n724), .B2(
        \registers[23][3] ), .ZN(n1298) );
  INV_X1 U2531 ( .A(n1299), .ZN(n3647) );
  AOI22_X1 U2532 ( .A1(DATAIN[4]), .A2(n723), .B1(n724), .B2(
        \registers[23][4] ), .ZN(n1299) );
  INV_X1 U2533 ( .A(n1300), .ZN(n3648) );
  AOI22_X1 U2534 ( .A1(DATAIN[5]), .A2(n722), .B1(n725), .B2(
        \registers[23][5] ), .ZN(n1300) );
  INV_X1 U2535 ( .A(n1301), .ZN(n3649) );
  AOI22_X1 U2536 ( .A1(DATAIN[6]), .A2(n723), .B1(n725), .B2(
        \registers[23][6] ), .ZN(n1301) );
  INV_X1 U2537 ( .A(n1302), .ZN(n3650) );
  AOI22_X1 U2538 ( .A1(DATAIN[7]), .A2(n722), .B1(n725), .B2(
        \registers[23][7] ), .ZN(n1302) );
  INV_X1 U2539 ( .A(n1303), .ZN(n3651) );
  AOI22_X1 U2540 ( .A1(DATAIN[8]), .A2(n723), .B1(n725), .B2(
        \registers[23][8] ), .ZN(n1303) );
  INV_X1 U2541 ( .A(n1304), .ZN(n3652) );
  AOI22_X1 U2542 ( .A1(DATAIN[9]), .A2(n723), .B1(n725), .B2(
        \registers[23][9] ), .ZN(n1304) );
  INV_X1 U2543 ( .A(n1305), .ZN(n3653) );
  AOI22_X1 U2544 ( .A1(DATAIN[10]), .A2(n723), .B1(n726), .B2(
        \registers[23][10] ), .ZN(n1305) );
  INV_X1 U2545 ( .A(n1306), .ZN(n3654) );
  AOI22_X1 U2546 ( .A1(DATAIN[11]), .A2(n723), .B1(n726), .B2(
        \registers[23][11] ), .ZN(n1306) );
  INV_X1 U2547 ( .A(n1307), .ZN(n3655) );
  AOI22_X1 U2548 ( .A1(DATAIN[12]), .A2(n723), .B1(n726), .B2(
        \registers[23][12] ), .ZN(n1307) );
  INV_X1 U2549 ( .A(n1308), .ZN(n3656) );
  AOI22_X1 U2550 ( .A1(DATAIN[13]), .A2(n723), .B1(n726), .B2(
        \registers[23][13] ), .ZN(n1308) );
  INV_X1 U2551 ( .A(n1309), .ZN(n3657) );
  AOI22_X1 U2552 ( .A1(DATAIN[14]), .A2(n723), .B1(n726), .B2(
        \registers[23][14] ), .ZN(n1309) );
  INV_X1 U2553 ( .A(n1310), .ZN(n3658) );
  AOI22_X1 U2554 ( .A1(DATAIN[15]), .A2(n723), .B1(n727), .B2(
        \registers[23][15] ), .ZN(n1310) );
  INV_X1 U2555 ( .A(n1311), .ZN(n3659) );
  AOI22_X1 U2556 ( .A1(DATAIN[16]), .A2(n723), .B1(n727), .B2(
        \registers[23][16] ), .ZN(n1311) );
  INV_X1 U2557 ( .A(n1312), .ZN(n3660) );
  AOI22_X1 U2558 ( .A1(DATAIN[17]), .A2(n723), .B1(n727), .B2(
        \registers[23][17] ), .ZN(n1312) );
  INV_X1 U2559 ( .A(n1313), .ZN(n3661) );
  AOI22_X1 U2560 ( .A1(DATAIN[18]), .A2(n723), .B1(n727), .B2(
        \registers[23][18] ), .ZN(n1313) );
  INV_X1 U2561 ( .A(n1314), .ZN(n3662) );
  AOI22_X1 U2562 ( .A1(DATAIN[19]), .A2(n723), .B1(n727), .B2(
        \registers[23][19] ), .ZN(n1314) );
  INV_X1 U2563 ( .A(n1315), .ZN(n3663) );
  AOI22_X1 U2564 ( .A1(DATAIN[20]), .A2(n722), .B1(n728), .B2(
        \registers[23][20] ), .ZN(n1315) );
  INV_X1 U2565 ( .A(n1316), .ZN(n3664) );
  AOI22_X1 U2566 ( .A1(DATAIN[21]), .A2(n722), .B1(n728), .B2(
        \registers[23][21] ), .ZN(n1316) );
  INV_X1 U2567 ( .A(n1317), .ZN(n3665) );
  AOI22_X1 U2568 ( .A1(DATAIN[22]), .A2(n722), .B1(n728), .B2(
        \registers[23][22] ), .ZN(n1317) );
  INV_X1 U2569 ( .A(n1328), .ZN(n3611) );
  AOI22_X1 U2570 ( .A1(DATAIN[0]), .A2(n714), .B1(n715), .B2(
        \registers[22][0] ), .ZN(n1328) );
  INV_X1 U2571 ( .A(n1330), .ZN(n3612) );
  AOI22_X1 U2572 ( .A1(DATAIN[1]), .A2(n713), .B1(n715), .B2(
        \registers[22][1] ), .ZN(n1330) );
  INV_X1 U2573 ( .A(n1331), .ZN(n3613) );
  AOI22_X1 U2574 ( .A1(DATAIN[2]), .A2(n714), .B1(n715), .B2(
        \registers[22][2] ), .ZN(n1331) );
  INV_X1 U2575 ( .A(n1332), .ZN(n3614) );
  AOI22_X1 U2576 ( .A1(DATAIN[3]), .A2(n713), .B1(n715), .B2(
        \registers[22][3] ), .ZN(n1332) );
  INV_X1 U2577 ( .A(n1333), .ZN(n3615) );
  AOI22_X1 U2578 ( .A1(DATAIN[4]), .A2(n714), .B1(n715), .B2(
        \registers[22][4] ), .ZN(n1333) );
  INV_X1 U2579 ( .A(n1334), .ZN(n3616) );
  AOI22_X1 U2580 ( .A1(DATAIN[5]), .A2(n713), .B1(n716), .B2(
        \registers[22][5] ), .ZN(n1334) );
  INV_X1 U2581 ( .A(n1335), .ZN(n3617) );
  AOI22_X1 U2582 ( .A1(DATAIN[6]), .A2(n714), .B1(n716), .B2(
        \registers[22][6] ), .ZN(n1335) );
  INV_X1 U2583 ( .A(n1336), .ZN(n3618) );
  AOI22_X1 U2584 ( .A1(DATAIN[7]), .A2(n713), .B1(n716), .B2(
        \registers[22][7] ), .ZN(n1336) );
  INV_X1 U2585 ( .A(n1337), .ZN(n3619) );
  AOI22_X1 U2586 ( .A1(DATAIN[8]), .A2(n714), .B1(n716), .B2(
        \registers[22][8] ), .ZN(n1337) );
  INV_X1 U2587 ( .A(n1338), .ZN(n3620) );
  AOI22_X1 U2588 ( .A1(DATAIN[9]), .A2(n714), .B1(n716), .B2(
        \registers[22][9] ), .ZN(n1338) );
  INV_X1 U2589 ( .A(n1339), .ZN(n3621) );
  AOI22_X1 U2590 ( .A1(DATAIN[10]), .A2(n714), .B1(n717), .B2(
        \registers[22][10] ), .ZN(n1339) );
  INV_X1 U2591 ( .A(n1340), .ZN(n3622) );
  AOI22_X1 U2592 ( .A1(DATAIN[11]), .A2(n714), .B1(n717), .B2(
        \registers[22][11] ), .ZN(n1340) );
  INV_X1 U2593 ( .A(n1341), .ZN(n3623) );
  AOI22_X1 U2594 ( .A1(DATAIN[12]), .A2(n714), .B1(n717), .B2(
        \registers[22][12] ), .ZN(n1341) );
  INV_X1 U2595 ( .A(n1342), .ZN(n3624) );
  AOI22_X1 U2596 ( .A1(DATAIN[13]), .A2(n714), .B1(n717), .B2(
        \registers[22][13] ), .ZN(n1342) );
  INV_X1 U2597 ( .A(n1343), .ZN(n3625) );
  AOI22_X1 U2598 ( .A1(DATAIN[14]), .A2(n714), .B1(n717), .B2(
        \registers[22][14] ), .ZN(n1343) );
  INV_X1 U2599 ( .A(n1344), .ZN(n3626) );
  AOI22_X1 U2600 ( .A1(DATAIN[15]), .A2(n714), .B1(n718), .B2(
        \registers[22][15] ), .ZN(n1344) );
  INV_X1 U2601 ( .A(n1345), .ZN(n3627) );
  AOI22_X1 U2602 ( .A1(DATAIN[16]), .A2(n714), .B1(n718), .B2(
        \registers[22][16] ), .ZN(n1345) );
  INV_X1 U2603 ( .A(n1346), .ZN(n3628) );
  AOI22_X1 U2604 ( .A1(DATAIN[17]), .A2(n714), .B1(n718), .B2(
        \registers[22][17] ), .ZN(n1346) );
  INV_X1 U2605 ( .A(n1347), .ZN(n3629) );
  AOI22_X1 U2606 ( .A1(DATAIN[18]), .A2(n714), .B1(n718), .B2(
        \registers[22][18] ), .ZN(n1347) );
  INV_X1 U2607 ( .A(n1348), .ZN(n3630) );
  AOI22_X1 U2608 ( .A1(DATAIN[19]), .A2(n714), .B1(n718), .B2(
        \registers[22][19] ), .ZN(n1348) );
  INV_X1 U2609 ( .A(n1349), .ZN(n3631) );
  AOI22_X1 U2610 ( .A1(DATAIN[20]), .A2(n713), .B1(n719), .B2(
        \registers[22][20] ), .ZN(n1349) );
  INV_X1 U2611 ( .A(n1350), .ZN(n3632) );
  AOI22_X1 U2612 ( .A1(DATAIN[21]), .A2(n713), .B1(n719), .B2(
        \registers[22][21] ), .ZN(n1350) );
  INV_X1 U2613 ( .A(n1351), .ZN(n3633) );
  AOI22_X1 U2614 ( .A1(DATAIN[22]), .A2(n713), .B1(n719), .B2(
        \registers[22][22] ), .ZN(n1351) );
  INV_X1 U2615 ( .A(n1363), .ZN(n3579) );
  AOI22_X1 U2616 ( .A1(DATAIN[0]), .A2(n687), .B1(n688), .B2(
        \registers[19][0] ), .ZN(n1363) );
  INV_X1 U2617 ( .A(n1365), .ZN(n3580) );
  AOI22_X1 U2618 ( .A1(DATAIN[1]), .A2(n686), .B1(n688), .B2(
        \registers[19][1] ), .ZN(n1365) );
  INV_X1 U2619 ( .A(n1366), .ZN(n3581) );
  AOI22_X1 U2620 ( .A1(DATAIN[2]), .A2(n687), .B1(n688), .B2(
        \registers[19][2] ), .ZN(n1366) );
  INV_X1 U2621 ( .A(n1367), .ZN(n3582) );
  AOI22_X1 U2622 ( .A1(DATAIN[3]), .A2(n686), .B1(n688), .B2(
        \registers[19][3] ), .ZN(n1367) );
  INV_X1 U2623 ( .A(n1368), .ZN(n3583) );
  AOI22_X1 U2624 ( .A1(DATAIN[4]), .A2(n687), .B1(n688), .B2(
        \registers[19][4] ), .ZN(n1368) );
  INV_X1 U2625 ( .A(n1369), .ZN(n3584) );
  AOI22_X1 U2626 ( .A1(DATAIN[5]), .A2(n686), .B1(n689), .B2(
        \registers[19][5] ), .ZN(n1369) );
  INV_X1 U2627 ( .A(n1370), .ZN(n3585) );
  AOI22_X1 U2628 ( .A1(DATAIN[6]), .A2(n687), .B1(n689), .B2(
        \registers[19][6] ), .ZN(n1370) );
  INV_X1 U2629 ( .A(n1371), .ZN(n3586) );
  AOI22_X1 U2630 ( .A1(DATAIN[7]), .A2(n686), .B1(n689), .B2(
        \registers[19][7] ), .ZN(n1371) );
  INV_X1 U2631 ( .A(n1372), .ZN(n3587) );
  AOI22_X1 U2632 ( .A1(DATAIN[8]), .A2(n687), .B1(n689), .B2(
        \registers[19][8] ), .ZN(n1372) );
  INV_X1 U2633 ( .A(n1373), .ZN(n3588) );
  AOI22_X1 U2634 ( .A1(DATAIN[9]), .A2(n687), .B1(n689), .B2(
        \registers[19][9] ), .ZN(n1373) );
  INV_X1 U2635 ( .A(n1374), .ZN(n3589) );
  AOI22_X1 U2636 ( .A1(DATAIN[10]), .A2(n687), .B1(n690), .B2(
        \registers[19][10] ), .ZN(n1374) );
  INV_X1 U2637 ( .A(n1375), .ZN(n3590) );
  AOI22_X1 U2638 ( .A1(DATAIN[11]), .A2(n687), .B1(n690), .B2(
        \registers[19][11] ), .ZN(n1375) );
  INV_X1 U2639 ( .A(n1376), .ZN(n3591) );
  AOI22_X1 U2640 ( .A1(DATAIN[12]), .A2(n687), .B1(n690), .B2(
        \registers[19][12] ), .ZN(n1376) );
  INV_X1 U2641 ( .A(n1377), .ZN(n3592) );
  AOI22_X1 U2642 ( .A1(DATAIN[13]), .A2(n687), .B1(n690), .B2(
        \registers[19][13] ), .ZN(n1377) );
  INV_X1 U2643 ( .A(n1378), .ZN(n3593) );
  AOI22_X1 U2644 ( .A1(DATAIN[14]), .A2(n687), .B1(n690), .B2(
        \registers[19][14] ), .ZN(n1378) );
  INV_X1 U2645 ( .A(n1379), .ZN(n3594) );
  AOI22_X1 U2646 ( .A1(DATAIN[15]), .A2(n687), .B1(n691), .B2(
        \registers[19][15] ), .ZN(n1379) );
  INV_X1 U2647 ( .A(n1380), .ZN(n3595) );
  AOI22_X1 U2648 ( .A1(DATAIN[16]), .A2(n687), .B1(n691), .B2(
        \registers[19][16] ), .ZN(n1380) );
  INV_X1 U2649 ( .A(n1381), .ZN(n3596) );
  AOI22_X1 U2650 ( .A1(DATAIN[17]), .A2(n687), .B1(n691), .B2(
        \registers[19][17] ), .ZN(n1381) );
  INV_X1 U2651 ( .A(n1382), .ZN(n3597) );
  AOI22_X1 U2652 ( .A1(DATAIN[18]), .A2(n687), .B1(n691), .B2(
        \registers[19][18] ), .ZN(n1382) );
  INV_X1 U2653 ( .A(n1383), .ZN(n3598) );
  AOI22_X1 U2654 ( .A1(DATAIN[19]), .A2(n687), .B1(n691), .B2(
        \registers[19][19] ), .ZN(n1383) );
  INV_X1 U2655 ( .A(n1384), .ZN(n3599) );
  AOI22_X1 U2656 ( .A1(DATAIN[20]), .A2(n686), .B1(n692), .B2(
        \registers[19][20] ), .ZN(n1384) );
  INV_X1 U2657 ( .A(n1385), .ZN(n3600) );
  AOI22_X1 U2658 ( .A1(DATAIN[21]), .A2(n686), .B1(n692), .B2(
        \registers[19][21] ), .ZN(n1385) );
  INV_X1 U2659 ( .A(n1386), .ZN(n3601) );
  AOI22_X1 U2660 ( .A1(DATAIN[22]), .A2(n686), .B1(n692), .B2(
        \registers[19][22] ), .ZN(n1386) );
  INV_X1 U2661 ( .A(n1396), .ZN(n3547) );
  AOI22_X1 U2662 ( .A1(DATAIN[0]), .A2(n678), .B1(n679), .B2(
        \registers[18][0] ), .ZN(n1396) );
  INV_X1 U2663 ( .A(n1398), .ZN(n3548) );
  AOI22_X1 U2664 ( .A1(DATAIN[1]), .A2(n677), .B1(n679), .B2(
        \registers[18][1] ), .ZN(n1398) );
  INV_X1 U2665 ( .A(n1399), .ZN(n3549) );
  AOI22_X1 U2666 ( .A1(DATAIN[2]), .A2(n678), .B1(n679), .B2(
        \registers[18][2] ), .ZN(n1399) );
  INV_X1 U2667 ( .A(n1400), .ZN(n3550) );
  AOI22_X1 U2668 ( .A1(DATAIN[3]), .A2(n677), .B1(n679), .B2(
        \registers[18][3] ), .ZN(n1400) );
  INV_X1 U2669 ( .A(n1401), .ZN(n3551) );
  AOI22_X1 U2670 ( .A1(DATAIN[4]), .A2(n678), .B1(n679), .B2(
        \registers[18][4] ), .ZN(n1401) );
  INV_X1 U2671 ( .A(n1402), .ZN(n3552) );
  AOI22_X1 U2672 ( .A1(DATAIN[5]), .A2(n677), .B1(n680), .B2(
        \registers[18][5] ), .ZN(n1402) );
  INV_X1 U2673 ( .A(n1403), .ZN(n3553) );
  AOI22_X1 U2674 ( .A1(DATAIN[6]), .A2(n678), .B1(n680), .B2(
        \registers[18][6] ), .ZN(n1403) );
  INV_X1 U2675 ( .A(n1404), .ZN(n3554) );
  AOI22_X1 U2676 ( .A1(DATAIN[7]), .A2(n677), .B1(n680), .B2(
        \registers[18][7] ), .ZN(n1404) );
  INV_X1 U2677 ( .A(n1405), .ZN(n3555) );
  AOI22_X1 U2678 ( .A1(DATAIN[8]), .A2(n678), .B1(n680), .B2(
        \registers[18][8] ), .ZN(n1405) );
  INV_X1 U2679 ( .A(n1406), .ZN(n3556) );
  AOI22_X1 U2680 ( .A1(DATAIN[9]), .A2(n678), .B1(n680), .B2(
        \registers[18][9] ), .ZN(n1406) );
  INV_X1 U2681 ( .A(n1407), .ZN(n3557) );
  AOI22_X1 U2682 ( .A1(DATAIN[10]), .A2(n678), .B1(n681), .B2(
        \registers[18][10] ), .ZN(n1407) );
  INV_X1 U2683 ( .A(n1408), .ZN(n3558) );
  AOI22_X1 U2684 ( .A1(DATAIN[11]), .A2(n678), .B1(n681), .B2(
        \registers[18][11] ), .ZN(n1408) );
  INV_X1 U2685 ( .A(n1409), .ZN(n3559) );
  AOI22_X1 U2686 ( .A1(DATAIN[12]), .A2(n678), .B1(n681), .B2(
        \registers[18][12] ), .ZN(n1409) );
  INV_X1 U2687 ( .A(n1410), .ZN(n3560) );
  AOI22_X1 U2688 ( .A1(DATAIN[13]), .A2(n678), .B1(n681), .B2(
        \registers[18][13] ), .ZN(n1410) );
  INV_X1 U2689 ( .A(n1411), .ZN(n3561) );
  AOI22_X1 U2690 ( .A1(DATAIN[14]), .A2(n678), .B1(n681), .B2(
        \registers[18][14] ), .ZN(n1411) );
  INV_X1 U2691 ( .A(n1412), .ZN(n3562) );
  AOI22_X1 U2692 ( .A1(DATAIN[15]), .A2(n678), .B1(n682), .B2(
        \registers[18][15] ), .ZN(n1412) );
  INV_X1 U2693 ( .A(n1413), .ZN(n3563) );
  AOI22_X1 U2694 ( .A1(DATAIN[16]), .A2(n678), .B1(n682), .B2(
        \registers[18][16] ), .ZN(n1413) );
  INV_X1 U2695 ( .A(n1414), .ZN(n3564) );
  AOI22_X1 U2696 ( .A1(DATAIN[17]), .A2(n678), .B1(n682), .B2(
        \registers[18][17] ), .ZN(n1414) );
  INV_X1 U2697 ( .A(n1415), .ZN(n3565) );
  AOI22_X1 U2698 ( .A1(DATAIN[18]), .A2(n678), .B1(n682), .B2(
        \registers[18][18] ), .ZN(n1415) );
  INV_X1 U2699 ( .A(n1416), .ZN(n3566) );
  AOI22_X1 U2700 ( .A1(DATAIN[19]), .A2(n678), .B1(n682), .B2(
        \registers[18][19] ), .ZN(n1416) );
  INV_X1 U2701 ( .A(n1417), .ZN(n3567) );
  AOI22_X1 U2702 ( .A1(DATAIN[20]), .A2(n677), .B1(n683), .B2(
        \registers[18][20] ), .ZN(n1417) );
  INV_X1 U2703 ( .A(n1418), .ZN(n3568) );
  AOI22_X1 U2704 ( .A1(DATAIN[21]), .A2(n677), .B1(n683), .B2(
        \registers[18][21] ), .ZN(n1418) );
  INV_X1 U2705 ( .A(n1419), .ZN(n3569) );
  AOI22_X1 U2706 ( .A1(DATAIN[22]), .A2(n677), .B1(n683), .B2(
        \registers[18][22] ), .ZN(n1419) );
  INV_X1 U2707 ( .A(n1434), .ZN(n3418) );
  AOI22_X1 U2708 ( .A1(DATAIN[0]), .A2(n569), .B1(n570), .B2(
        \registers[13][0] ), .ZN(n1434) );
  INV_X1 U2709 ( .A(n1436), .ZN(n3419) );
  AOI22_X1 U2710 ( .A1(DATAIN[1]), .A2(n568), .B1(n570), .B2(
        \registers[13][1] ), .ZN(n1436) );
  INV_X1 U2711 ( .A(n1437), .ZN(n3420) );
  AOI22_X1 U2712 ( .A1(DATAIN[2]), .A2(n569), .B1(n570), .B2(
        \registers[13][2] ), .ZN(n1437) );
  INV_X1 U2713 ( .A(n1438), .ZN(n3421) );
  AOI22_X1 U2714 ( .A1(DATAIN[3]), .A2(n568), .B1(n570), .B2(
        \registers[13][3] ), .ZN(n1438) );
  INV_X1 U2715 ( .A(n1439), .ZN(n3422) );
  AOI22_X1 U2716 ( .A1(DATAIN[4]), .A2(n569), .B1(n570), .B2(
        \registers[13][4] ), .ZN(n1439) );
  INV_X1 U2717 ( .A(n1440), .ZN(n3423) );
  AOI22_X1 U2718 ( .A1(DATAIN[5]), .A2(n568), .B1(n571), .B2(
        \registers[13][5] ), .ZN(n1440) );
  INV_X1 U2719 ( .A(n1441), .ZN(n3424) );
  AOI22_X1 U2720 ( .A1(DATAIN[6]), .A2(n569), .B1(n571), .B2(
        \registers[13][6] ), .ZN(n1441) );
  INV_X1 U2721 ( .A(n1442), .ZN(n3425) );
  AOI22_X1 U2722 ( .A1(DATAIN[7]), .A2(n568), .B1(n571), .B2(
        \registers[13][7] ), .ZN(n1442) );
  INV_X1 U2723 ( .A(n1443), .ZN(n3426) );
  AOI22_X1 U2724 ( .A1(DATAIN[8]), .A2(n569), .B1(n571), .B2(
        \registers[13][8] ), .ZN(n1443) );
  INV_X1 U2725 ( .A(n1444), .ZN(n3427) );
  AOI22_X1 U2726 ( .A1(DATAIN[9]), .A2(n569), .B1(n571), .B2(
        \registers[13][9] ), .ZN(n1444) );
  INV_X1 U2727 ( .A(n1445), .ZN(n3428) );
  AOI22_X1 U2728 ( .A1(DATAIN[10]), .A2(n569), .B1(n572), .B2(
        \registers[13][10] ), .ZN(n1445) );
  INV_X1 U2729 ( .A(n1446), .ZN(n3429) );
  AOI22_X1 U2730 ( .A1(DATAIN[11]), .A2(n569), .B1(n572), .B2(
        \registers[13][11] ), .ZN(n1446) );
  INV_X1 U2731 ( .A(n1447), .ZN(n3430) );
  AOI22_X1 U2732 ( .A1(DATAIN[12]), .A2(n569), .B1(n572), .B2(
        \registers[13][12] ), .ZN(n1447) );
  INV_X1 U2733 ( .A(n1448), .ZN(n3431) );
  AOI22_X1 U2734 ( .A1(DATAIN[13]), .A2(n569), .B1(n572), .B2(
        \registers[13][13] ), .ZN(n1448) );
  INV_X1 U2735 ( .A(n1449), .ZN(n3432) );
  AOI22_X1 U2736 ( .A1(DATAIN[14]), .A2(n569), .B1(n572), .B2(
        \registers[13][14] ), .ZN(n1449) );
  INV_X1 U2737 ( .A(n1450), .ZN(n3433) );
  AOI22_X1 U2738 ( .A1(DATAIN[15]), .A2(n569), .B1(n573), .B2(
        \registers[13][15] ), .ZN(n1450) );
  INV_X1 U2739 ( .A(n1451), .ZN(n3434) );
  AOI22_X1 U2740 ( .A1(DATAIN[16]), .A2(n569), .B1(n573), .B2(
        \registers[13][16] ), .ZN(n1451) );
  INV_X1 U2741 ( .A(n1452), .ZN(n3435) );
  AOI22_X1 U2742 ( .A1(DATAIN[17]), .A2(n569), .B1(n573), .B2(
        \registers[13][17] ), .ZN(n1452) );
  INV_X1 U2743 ( .A(n1453), .ZN(n3436) );
  AOI22_X1 U2744 ( .A1(DATAIN[18]), .A2(n569), .B1(n573), .B2(
        \registers[13][18] ), .ZN(n1453) );
  INV_X1 U2745 ( .A(n1454), .ZN(n3437) );
  AOI22_X1 U2746 ( .A1(DATAIN[19]), .A2(n569), .B1(n573), .B2(
        \registers[13][19] ), .ZN(n1454) );
  INV_X1 U2747 ( .A(n1455), .ZN(n3438) );
  AOI22_X1 U2748 ( .A1(DATAIN[20]), .A2(n568), .B1(n574), .B2(
        \registers[13][20] ), .ZN(n1455) );
  INV_X1 U2749 ( .A(n1456), .ZN(n3439) );
  AOI22_X1 U2750 ( .A1(DATAIN[21]), .A2(n568), .B1(n574), .B2(
        \registers[13][21] ), .ZN(n1456) );
  INV_X1 U2751 ( .A(n1457), .ZN(n3440) );
  AOI22_X1 U2752 ( .A1(DATAIN[22]), .A2(n568), .B1(n574), .B2(
        \registers[13][22] ), .ZN(n1457) );
  INV_X1 U2753 ( .A(n1467), .ZN(n3386) );
  AOI22_X1 U2754 ( .A1(DATAIN[0]), .A2(n560), .B1(n561), .B2(
        \registers[12][0] ), .ZN(n1467) );
  INV_X1 U2755 ( .A(n1469), .ZN(n3387) );
  AOI22_X1 U2756 ( .A1(DATAIN[1]), .A2(n559), .B1(n561), .B2(
        \registers[12][1] ), .ZN(n1469) );
  INV_X1 U2757 ( .A(n1470), .ZN(n3388) );
  AOI22_X1 U2758 ( .A1(DATAIN[2]), .A2(n560), .B1(n561), .B2(
        \registers[12][2] ), .ZN(n1470) );
  INV_X1 U2759 ( .A(n1471), .ZN(n3389) );
  AOI22_X1 U2760 ( .A1(DATAIN[3]), .A2(n559), .B1(n561), .B2(
        \registers[12][3] ), .ZN(n1471) );
  INV_X1 U2761 ( .A(n1472), .ZN(n3390) );
  AOI22_X1 U2762 ( .A1(DATAIN[4]), .A2(n560), .B1(n561), .B2(
        \registers[12][4] ), .ZN(n1472) );
  INV_X1 U2763 ( .A(n1473), .ZN(n3391) );
  AOI22_X1 U2764 ( .A1(DATAIN[5]), .A2(n559), .B1(n562), .B2(
        \registers[12][5] ), .ZN(n1473) );
  INV_X1 U2765 ( .A(n1474), .ZN(n3392) );
  AOI22_X1 U2766 ( .A1(DATAIN[6]), .A2(n560), .B1(n562), .B2(
        \registers[12][6] ), .ZN(n1474) );
  INV_X1 U2767 ( .A(n1475), .ZN(n3393) );
  AOI22_X1 U2768 ( .A1(DATAIN[7]), .A2(n559), .B1(n562), .B2(
        \registers[12][7] ), .ZN(n1475) );
  INV_X1 U2769 ( .A(n1476), .ZN(n3394) );
  AOI22_X1 U2770 ( .A1(DATAIN[8]), .A2(n560), .B1(n562), .B2(
        \registers[12][8] ), .ZN(n1476) );
  INV_X1 U2771 ( .A(n1477), .ZN(n3395) );
  AOI22_X1 U2772 ( .A1(DATAIN[9]), .A2(n560), .B1(n562), .B2(
        \registers[12][9] ), .ZN(n1477) );
  INV_X1 U2773 ( .A(n1478), .ZN(n3396) );
  AOI22_X1 U2774 ( .A1(DATAIN[10]), .A2(n560), .B1(n563), .B2(
        \registers[12][10] ), .ZN(n1478) );
  INV_X1 U2775 ( .A(n1479), .ZN(n3397) );
  AOI22_X1 U2776 ( .A1(DATAIN[11]), .A2(n560), .B1(n563), .B2(
        \registers[12][11] ), .ZN(n1479) );
  INV_X1 U2777 ( .A(n1480), .ZN(n3398) );
  AOI22_X1 U2778 ( .A1(DATAIN[12]), .A2(n560), .B1(n563), .B2(
        \registers[12][12] ), .ZN(n1480) );
  INV_X1 U2779 ( .A(n1481), .ZN(n3399) );
  AOI22_X1 U2780 ( .A1(DATAIN[13]), .A2(n560), .B1(n563), .B2(
        \registers[12][13] ), .ZN(n1481) );
  INV_X1 U2781 ( .A(n1482), .ZN(n3400) );
  AOI22_X1 U2782 ( .A1(DATAIN[14]), .A2(n560), .B1(n563), .B2(
        \registers[12][14] ), .ZN(n1482) );
  INV_X1 U2783 ( .A(n1483), .ZN(n3401) );
  AOI22_X1 U2784 ( .A1(DATAIN[15]), .A2(n560), .B1(n564), .B2(
        \registers[12][15] ), .ZN(n1483) );
  INV_X1 U2785 ( .A(n1484), .ZN(n3402) );
  AOI22_X1 U2786 ( .A1(DATAIN[16]), .A2(n560), .B1(n564), .B2(
        \registers[12][16] ), .ZN(n1484) );
  INV_X1 U2787 ( .A(n1485), .ZN(n3403) );
  AOI22_X1 U2788 ( .A1(DATAIN[17]), .A2(n560), .B1(n564), .B2(
        \registers[12][17] ), .ZN(n1485) );
  INV_X1 U2789 ( .A(n1486), .ZN(n3404) );
  AOI22_X1 U2790 ( .A1(DATAIN[18]), .A2(n560), .B1(n564), .B2(
        \registers[12][18] ), .ZN(n1486) );
  INV_X1 U2791 ( .A(n1487), .ZN(n3405) );
  AOI22_X1 U2792 ( .A1(DATAIN[19]), .A2(n560), .B1(n564), .B2(
        \registers[12][19] ), .ZN(n1487) );
  INV_X1 U2793 ( .A(n1488), .ZN(n3406) );
  AOI22_X1 U2794 ( .A1(DATAIN[20]), .A2(n559), .B1(n565), .B2(
        \registers[12][20] ), .ZN(n1488) );
  INV_X1 U2795 ( .A(n1489), .ZN(n3407) );
  AOI22_X1 U2796 ( .A1(DATAIN[21]), .A2(n559), .B1(n565), .B2(
        \registers[12][21] ), .ZN(n1489) );
  INV_X1 U2797 ( .A(n1490), .ZN(n3408) );
  AOI22_X1 U2798 ( .A1(DATAIN[22]), .A2(n559), .B1(n565), .B2(
        \registers[12][22] ), .ZN(n1490) );
  INV_X1 U2799 ( .A(n1502), .ZN(n3354) );
  AOI22_X1 U2800 ( .A1(DATAIN[0]), .A2(n405), .B1(n406), .B2(\registers[9][0] ), .ZN(n1502) );
  INV_X1 U2801 ( .A(n1504), .ZN(n3355) );
  AOI22_X1 U2802 ( .A1(DATAIN[1]), .A2(n404), .B1(n406), .B2(\registers[9][1] ), .ZN(n1504) );
  INV_X1 U2803 ( .A(n1505), .ZN(n3356) );
  AOI22_X1 U2804 ( .A1(DATAIN[2]), .A2(n405), .B1(n406), .B2(\registers[9][2] ), .ZN(n1505) );
  INV_X1 U2805 ( .A(n1506), .ZN(n3357) );
  AOI22_X1 U2806 ( .A1(DATAIN[3]), .A2(n404), .B1(n406), .B2(\registers[9][3] ), .ZN(n1506) );
  INV_X1 U2807 ( .A(n1507), .ZN(n3358) );
  AOI22_X1 U2808 ( .A1(DATAIN[4]), .A2(n405), .B1(n406), .B2(\registers[9][4] ), .ZN(n1507) );
  INV_X1 U2809 ( .A(n1508), .ZN(n3359) );
  AOI22_X1 U2810 ( .A1(DATAIN[5]), .A2(n404), .B1(n407), .B2(\registers[9][5] ), .ZN(n1508) );
  INV_X1 U2811 ( .A(n1509), .ZN(n3360) );
  AOI22_X1 U2812 ( .A1(DATAIN[6]), .A2(n405), .B1(n407), .B2(\registers[9][6] ), .ZN(n1509) );
  INV_X1 U2813 ( .A(n1510), .ZN(n3361) );
  AOI22_X1 U2814 ( .A1(DATAIN[7]), .A2(n404), .B1(n407), .B2(\registers[9][7] ), .ZN(n1510) );
  INV_X1 U2815 ( .A(n1511), .ZN(n3362) );
  AOI22_X1 U2816 ( .A1(DATAIN[8]), .A2(n405), .B1(n407), .B2(\registers[9][8] ), .ZN(n1511) );
  INV_X1 U2817 ( .A(n1512), .ZN(n3363) );
  AOI22_X1 U2818 ( .A1(DATAIN[9]), .A2(n405), .B1(n407), .B2(\registers[9][9] ), .ZN(n1512) );
  INV_X1 U2819 ( .A(n1513), .ZN(n3364) );
  AOI22_X1 U2820 ( .A1(DATAIN[10]), .A2(n405), .B1(n408), .B2(
        \registers[9][10] ), .ZN(n1513) );
  INV_X1 U2821 ( .A(n1514), .ZN(n3365) );
  AOI22_X1 U2822 ( .A1(DATAIN[11]), .A2(n405), .B1(n408), .B2(
        \registers[9][11] ), .ZN(n1514) );
  INV_X1 U2823 ( .A(n1515), .ZN(n3366) );
  AOI22_X1 U2824 ( .A1(DATAIN[12]), .A2(n405), .B1(n408), .B2(
        \registers[9][12] ), .ZN(n1515) );
  INV_X1 U2825 ( .A(n1516), .ZN(n3367) );
  AOI22_X1 U2826 ( .A1(DATAIN[13]), .A2(n405), .B1(n408), .B2(
        \registers[9][13] ), .ZN(n1516) );
  INV_X1 U2827 ( .A(n1517), .ZN(n3368) );
  AOI22_X1 U2828 ( .A1(DATAIN[14]), .A2(n405), .B1(n408), .B2(
        \registers[9][14] ), .ZN(n1517) );
  INV_X1 U2829 ( .A(n1518), .ZN(n3369) );
  AOI22_X1 U2830 ( .A1(DATAIN[15]), .A2(n405), .B1(n409), .B2(
        \registers[9][15] ), .ZN(n1518) );
  INV_X1 U2831 ( .A(n1519), .ZN(n3370) );
  AOI22_X1 U2832 ( .A1(DATAIN[16]), .A2(n405), .B1(n409), .B2(
        \registers[9][16] ), .ZN(n1519) );
  INV_X1 U2833 ( .A(n1520), .ZN(n3371) );
  AOI22_X1 U2834 ( .A1(DATAIN[17]), .A2(n405), .B1(n409), .B2(
        \registers[9][17] ), .ZN(n1520) );
  INV_X1 U2835 ( .A(n1521), .ZN(n3372) );
  AOI22_X1 U2836 ( .A1(DATAIN[18]), .A2(n405), .B1(n409), .B2(
        \registers[9][18] ), .ZN(n1521) );
  INV_X1 U2837 ( .A(n1522), .ZN(n3373) );
  AOI22_X1 U2838 ( .A1(DATAIN[19]), .A2(n405), .B1(n409), .B2(
        \registers[9][19] ), .ZN(n1522) );
  INV_X1 U2839 ( .A(n1523), .ZN(n3374) );
  AOI22_X1 U2840 ( .A1(DATAIN[20]), .A2(n404), .B1(n410), .B2(
        \registers[9][20] ), .ZN(n1523) );
  INV_X1 U2841 ( .A(n1524), .ZN(n3375) );
  AOI22_X1 U2842 ( .A1(DATAIN[21]), .A2(n404), .B1(n410), .B2(
        \registers[9][21] ), .ZN(n1524) );
  INV_X1 U2843 ( .A(n1525), .ZN(n3376) );
  AOI22_X1 U2844 ( .A1(DATAIN[22]), .A2(n404), .B1(n410), .B2(
        \registers[9][22] ), .ZN(n1525) );
  INV_X1 U2845 ( .A(n1535), .ZN(n3322) );
  AOI22_X1 U2846 ( .A1(DATAIN[0]), .A2(n396), .B1(n397), .B2(\registers[8][0] ), .ZN(n1535) );
  INV_X1 U2847 ( .A(n1537), .ZN(n3323) );
  AOI22_X1 U2848 ( .A1(DATAIN[1]), .A2(n395), .B1(n397), .B2(\registers[8][1] ), .ZN(n1537) );
  INV_X1 U2849 ( .A(n1538), .ZN(n3324) );
  AOI22_X1 U2850 ( .A1(DATAIN[2]), .A2(n396), .B1(n397), .B2(\registers[8][2] ), .ZN(n1538) );
  INV_X1 U2851 ( .A(n1539), .ZN(n3325) );
  AOI22_X1 U2852 ( .A1(DATAIN[3]), .A2(n395), .B1(n397), .B2(\registers[8][3] ), .ZN(n1539) );
  INV_X1 U2853 ( .A(n1540), .ZN(n3326) );
  AOI22_X1 U2854 ( .A1(DATAIN[4]), .A2(n396), .B1(n397), .B2(\registers[8][4] ), .ZN(n1540) );
  INV_X1 U2855 ( .A(n1541), .ZN(n3327) );
  AOI22_X1 U2856 ( .A1(DATAIN[5]), .A2(n395), .B1(n398), .B2(\registers[8][5] ), .ZN(n1541) );
  INV_X1 U2857 ( .A(n1542), .ZN(n3328) );
  AOI22_X1 U2858 ( .A1(DATAIN[6]), .A2(n396), .B1(n398), .B2(\registers[8][6] ), .ZN(n1542) );
  INV_X1 U2859 ( .A(n1543), .ZN(n3329) );
  AOI22_X1 U2860 ( .A1(DATAIN[7]), .A2(n395), .B1(n398), .B2(\registers[8][7] ), .ZN(n1543) );
  INV_X1 U2861 ( .A(n1544), .ZN(n3330) );
  AOI22_X1 U2862 ( .A1(DATAIN[8]), .A2(n396), .B1(n398), .B2(\registers[8][8] ), .ZN(n1544) );
  INV_X1 U2863 ( .A(n1545), .ZN(n3331) );
  AOI22_X1 U2864 ( .A1(DATAIN[9]), .A2(n396), .B1(n398), .B2(\registers[8][9] ), .ZN(n1545) );
  INV_X1 U2865 ( .A(n1546), .ZN(n3332) );
  AOI22_X1 U2866 ( .A1(DATAIN[10]), .A2(n396), .B1(n399), .B2(
        \registers[8][10] ), .ZN(n1546) );
  INV_X1 U2867 ( .A(n1547), .ZN(n3333) );
  AOI22_X1 U2868 ( .A1(DATAIN[11]), .A2(n396), .B1(n399), .B2(
        \registers[8][11] ), .ZN(n1547) );
  INV_X1 U2869 ( .A(n1548), .ZN(n3334) );
  AOI22_X1 U2870 ( .A1(DATAIN[12]), .A2(n396), .B1(n399), .B2(
        \registers[8][12] ), .ZN(n1548) );
  INV_X1 U2871 ( .A(n1549), .ZN(n3335) );
  AOI22_X1 U2872 ( .A1(DATAIN[13]), .A2(n396), .B1(n399), .B2(
        \registers[8][13] ), .ZN(n1549) );
  INV_X1 U2873 ( .A(n1550), .ZN(n3336) );
  AOI22_X1 U2874 ( .A1(DATAIN[14]), .A2(n396), .B1(n399), .B2(
        \registers[8][14] ), .ZN(n1550) );
  INV_X1 U2875 ( .A(n1551), .ZN(n3337) );
  AOI22_X1 U2876 ( .A1(DATAIN[15]), .A2(n396), .B1(n400), .B2(
        \registers[8][15] ), .ZN(n1551) );
  INV_X1 U2877 ( .A(n1552), .ZN(n3338) );
  AOI22_X1 U2878 ( .A1(DATAIN[16]), .A2(n396), .B1(n400), .B2(
        \registers[8][16] ), .ZN(n1552) );
  INV_X1 U2879 ( .A(n1553), .ZN(n3339) );
  AOI22_X1 U2880 ( .A1(DATAIN[17]), .A2(n396), .B1(n400), .B2(
        \registers[8][17] ), .ZN(n1553) );
  INV_X1 U2881 ( .A(n1554), .ZN(n3340) );
  AOI22_X1 U2882 ( .A1(DATAIN[18]), .A2(n396), .B1(n400), .B2(
        \registers[8][18] ), .ZN(n1554) );
  INV_X1 U2883 ( .A(n1555), .ZN(n3341) );
  AOI22_X1 U2884 ( .A1(DATAIN[19]), .A2(n396), .B1(n400), .B2(
        \registers[8][19] ), .ZN(n1555) );
  INV_X1 U2885 ( .A(n1556), .ZN(n3342) );
  AOI22_X1 U2886 ( .A1(DATAIN[20]), .A2(n395), .B1(n401), .B2(
        \registers[8][20] ), .ZN(n1556) );
  INV_X1 U2887 ( .A(n1557), .ZN(n3343) );
  AOI22_X1 U2888 ( .A1(DATAIN[21]), .A2(n395), .B1(n401), .B2(
        \registers[8][21] ), .ZN(n1557) );
  INV_X1 U2889 ( .A(n1558), .ZN(n3344) );
  AOI22_X1 U2890 ( .A1(DATAIN[22]), .A2(n395), .B1(n401), .B2(
        \registers[8][22] ), .ZN(n1558) );
  INV_X1 U2891 ( .A(n1120), .ZN(n3482) );
  AOI22_X1 U2892 ( .A1(DATAIN[0]), .A2(n868), .B1(n869), .B2(\registers[1][0] ), .ZN(n1120) );
  INV_X1 U2893 ( .A(n1122), .ZN(n3483) );
  AOI22_X1 U2894 ( .A1(DATAIN[1]), .A2(n867), .B1(n869), .B2(\registers[1][1] ), .ZN(n1122) );
  INV_X1 U2895 ( .A(n1123), .ZN(n3484) );
  AOI22_X1 U2896 ( .A1(DATAIN[2]), .A2(n868), .B1(n869), .B2(\registers[1][2] ), .ZN(n1123) );
  INV_X1 U2897 ( .A(n1124), .ZN(n3485) );
  AOI22_X1 U2898 ( .A1(DATAIN[3]), .A2(n867), .B1(n869), .B2(\registers[1][3] ), .ZN(n1124) );
  INV_X1 U2899 ( .A(n1125), .ZN(n3486) );
  AOI22_X1 U2900 ( .A1(DATAIN[4]), .A2(n868), .B1(n869), .B2(\registers[1][4] ), .ZN(n1125) );
  INV_X1 U2901 ( .A(n1126), .ZN(n3487) );
  AOI22_X1 U2902 ( .A1(DATAIN[5]), .A2(n867), .B1(n870), .B2(\registers[1][5] ), .ZN(n1126) );
  INV_X1 U2903 ( .A(n1127), .ZN(n3488) );
  AOI22_X1 U2904 ( .A1(DATAIN[6]), .A2(n868), .B1(n870), .B2(\registers[1][6] ), .ZN(n1127) );
  INV_X1 U2905 ( .A(n1128), .ZN(n3489) );
  AOI22_X1 U2906 ( .A1(DATAIN[7]), .A2(n867), .B1(n870), .B2(\registers[1][7] ), .ZN(n1128) );
  INV_X1 U2907 ( .A(n1129), .ZN(n3490) );
  AOI22_X1 U2908 ( .A1(DATAIN[8]), .A2(n868), .B1(n870), .B2(\registers[1][8] ), .ZN(n1129) );
  INV_X1 U2909 ( .A(n1130), .ZN(n3491) );
  AOI22_X1 U2910 ( .A1(DATAIN[9]), .A2(n868), .B1(n870), .B2(\registers[1][9] ), .ZN(n1130) );
  INV_X1 U2911 ( .A(n1131), .ZN(n3492) );
  AOI22_X1 U2912 ( .A1(DATAIN[10]), .A2(n868), .B1(n871), .B2(
        \registers[1][10] ), .ZN(n1131) );
  INV_X1 U2913 ( .A(n1132), .ZN(n3493) );
  AOI22_X1 U2914 ( .A1(DATAIN[11]), .A2(n868), .B1(n871), .B2(
        \registers[1][11] ), .ZN(n1132) );
  INV_X1 U2915 ( .A(n1133), .ZN(n3494) );
  AOI22_X1 U2916 ( .A1(DATAIN[12]), .A2(n868), .B1(n871), .B2(
        \registers[1][12] ), .ZN(n1133) );
  INV_X1 U2917 ( .A(n1134), .ZN(n3495) );
  AOI22_X1 U2918 ( .A1(DATAIN[13]), .A2(n868), .B1(n871), .B2(
        \registers[1][13] ), .ZN(n1134) );
  INV_X1 U2919 ( .A(n1135), .ZN(n3496) );
  AOI22_X1 U2920 ( .A1(DATAIN[14]), .A2(n868), .B1(n871), .B2(
        \registers[1][14] ), .ZN(n1135) );
  INV_X1 U2921 ( .A(n1136), .ZN(n3497) );
  AOI22_X1 U2922 ( .A1(DATAIN[15]), .A2(n868), .B1(n872), .B2(
        \registers[1][15] ), .ZN(n1136) );
  INV_X1 U2923 ( .A(n1137), .ZN(n3498) );
  AOI22_X1 U2924 ( .A1(DATAIN[16]), .A2(n868), .B1(n872), .B2(
        \registers[1][16] ), .ZN(n1137) );
  INV_X1 U2925 ( .A(n1138), .ZN(n3499) );
  AOI22_X1 U2926 ( .A1(DATAIN[17]), .A2(n868), .B1(n872), .B2(
        \registers[1][17] ), .ZN(n1138) );
  INV_X1 U2927 ( .A(n1139), .ZN(n3500) );
  AOI22_X1 U2928 ( .A1(DATAIN[18]), .A2(n868), .B1(n872), .B2(
        \registers[1][18] ), .ZN(n1139) );
  INV_X1 U2929 ( .A(n1140), .ZN(n3501) );
  AOI22_X1 U2930 ( .A1(DATAIN[19]), .A2(n868), .B1(n872), .B2(
        \registers[1][19] ), .ZN(n1140) );
  INV_X1 U2931 ( .A(n1141), .ZN(n3502) );
  AOI22_X1 U2932 ( .A1(DATAIN[20]), .A2(n867), .B1(n873), .B2(
        \registers[1][20] ), .ZN(n1141) );
  INV_X1 U2933 ( .A(n1142), .ZN(n3503) );
  AOI22_X1 U2934 ( .A1(DATAIN[21]), .A2(n867), .B1(n873), .B2(
        \registers[1][21] ), .ZN(n1142) );
  INV_X1 U2935 ( .A(n1143), .ZN(n3504) );
  AOI22_X1 U2936 ( .A1(DATAIN[22]), .A2(n867), .B1(n873), .B2(
        \registers[1][22] ), .ZN(n1143) );
  INV_X1 U2937 ( .A(n1183), .ZN(n3794) );
  AOI22_X1 U2938 ( .A1(DATAIN[23]), .A2(n776), .B1(n782), .B2(
        \registers[29][23] ), .ZN(n1183) );
  INV_X1 U2939 ( .A(n1184), .ZN(n3795) );
  AOI22_X1 U2940 ( .A1(DATAIN[24]), .A2(n776), .B1(n782), .B2(
        \registers[29][24] ), .ZN(n1184) );
  INV_X1 U2941 ( .A(n1185), .ZN(n3796) );
  AOI22_X1 U2942 ( .A1(DATAIN[25]), .A2(n776), .B1(n783), .B2(
        \registers[29][25] ), .ZN(n1185) );
  INV_X1 U2943 ( .A(n1186), .ZN(n3797) );
  AOI22_X1 U2944 ( .A1(DATAIN[26]), .A2(n776), .B1(n783), .B2(
        \registers[29][26] ), .ZN(n1186) );
  INV_X1 U2945 ( .A(n1187), .ZN(n3798) );
  AOI22_X1 U2946 ( .A1(DATAIN[27]), .A2(n776), .B1(n783), .B2(
        \registers[29][27] ), .ZN(n1187) );
  INV_X1 U2947 ( .A(n1188), .ZN(n3799) );
  AOI22_X1 U2948 ( .A1(DATAIN[28]), .A2(n776), .B1(n783), .B2(
        \registers[29][28] ), .ZN(n1188) );
  INV_X1 U2949 ( .A(n1189), .ZN(n3800) );
  AOI22_X1 U2950 ( .A1(DATAIN[29]), .A2(n776), .B1(n783), .B2(
        \registers[29][29] ), .ZN(n1189) );
  INV_X1 U2951 ( .A(n1190), .ZN(n3801) );
  AOI22_X1 U2952 ( .A1(DATAIN[30]), .A2(n776), .B1(n784), .B2(
        \registers[29][30] ), .ZN(n1190) );
  INV_X1 U2953 ( .A(n1191), .ZN(n3802) );
  AOI22_X1 U2954 ( .A1(DATAIN[31]), .A2(n776), .B1(n784), .B2(
        \registers[29][31] ), .ZN(n1191) );
  INV_X1 U2955 ( .A(n1216), .ZN(n3762) );
  AOI22_X1 U2956 ( .A1(DATAIN[23]), .A2(n767), .B1(n773), .B2(
        \registers[28][23] ), .ZN(n1216) );
  INV_X1 U2957 ( .A(n1217), .ZN(n3763) );
  AOI22_X1 U2958 ( .A1(DATAIN[24]), .A2(n767), .B1(n773), .B2(
        \registers[28][24] ), .ZN(n1217) );
  INV_X1 U2959 ( .A(n1218), .ZN(n3764) );
  AOI22_X1 U2960 ( .A1(DATAIN[25]), .A2(n767), .B1(n774), .B2(
        \registers[28][25] ), .ZN(n1218) );
  INV_X1 U2961 ( .A(n1219), .ZN(n3765) );
  AOI22_X1 U2962 ( .A1(DATAIN[26]), .A2(n767), .B1(n774), .B2(
        \registers[28][26] ), .ZN(n1219) );
  INV_X1 U2963 ( .A(n1220), .ZN(n3766) );
  AOI22_X1 U2964 ( .A1(DATAIN[27]), .A2(n767), .B1(n774), .B2(
        \registers[28][27] ), .ZN(n1220) );
  INV_X1 U2965 ( .A(n1221), .ZN(n3767) );
  AOI22_X1 U2966 ( .A1(DATAIN[28]), .A2(n767), .B1(n774), .B2(
        \registers[28][28] ), .ZN(n1221) );
  INV_X1 U2967 ( .A(n1222), .ZN(n3768) );
  AOI22_X1 U2968 ( .A1(DATAIN[29]), .A2(n767), .B1(n774), .B2(
        \registers[28][29] ), .ZN(n1222) );
  INV_X1 U2969 ( .A(n1223), .ZN(n3769) );
  AOI22_X1 U2970 ( .A1(DATAIN[30]), .A2(n767), .B1(n775), .B2(
        \registers[28][30] ), .ZN(n1223) );
  INV_X1 U2971 ( .A(n1224), .ZN(n3770) );
  AOI22_X1 U2972 ( .A1(DATAIN[31]), .A2(n767), .B1(n775), .B2(
        \registers[28][31] ), .ZN(n1224) );
  INV_X1 U2973 ( .A(n1251), .ZN(n3730) );
  AOI22_X1 U2974 ( .A1(DATAIN[23]), .A2(n740), .B1(n746), .B2(
        \registers[25][23] ), .ZN(n1251) );
  INV_X1 U2975 ( .A(n1252), .ZN(n3731) );
  AOI22_X1 U2976 ( .A1(DATAIN[24]), .A2(n740), .B1(n746), .B2(
        \registers[25][24] ), .ZN(n1252) );
  INV_X1 U2977 ( .A(n1253), .ZN(n3732) );
  AOI22_X1 U2978 ( .A1(DATAIN[25]), .A2(n740), .B1(n747), .B2(
        \registers[25][25] ), .ZN(n1253) );
  INV_X1 U2979 ( .A(n1254), .ZN(n3733) );
  AOI22_X1 U2980 ( .A1(DATAIN[26]), .A2(n740), .B1(n747), .B2(
        \registers[25][26] ), .ZN(n1254) );
  INV_X1 U2981 ( .A(n1255), .ZN(n3734) );
  AOI22_X1 U2982 ( .A1(DATAIN[27]), .A2(n740), .B1(n747), .B2(
        \registers[25][27] ), .ZN(n1255) );
  INV_X1 U2983 ( .A(n1256), .ZN(n3735) );
  AOI22_X1 U2984 ( .A1(DATAIN[28]), .A2(n740), .B1(n747), .B2(
        \registers[25][28] ), .ZN(n1256) );
  INV_X1 U2985 ( .A(n1257), .ZN(n3736) );
  AOI22_X1 U2986 ( .A1(DATAIN[29]), .A2(n740), .B1(n747), .B2(
        \registers[25][29] ), .ZN(n1257) );
  INV_X1 U2987 ( .A(n1258), .ZN(n3737) );
  AOI22_X1 U2988 ( .A1(DATAIN[30]), .A2(n740), .B1(n748), .B2(
        \registers[25][30] ), .ZN(n1258) );
  INV_X1 U2989 ( .A(n1259), .ZN(n3738) );
  AOI22_X1 U2990 ( .A1(DATAIN[31]), .A2(n740), .B1(n748), .B2(
        \registers[25][31] ), .ZN(n1259) );
  INV_X1 U2991 ( .A(n1284), .ZN(n3698) );
  AOI22_X1 U2992 ( .A1(DATAIN[23]), .A2(n731), .B1(n737), .B2(
        \registers[24][23] ), .ZN(n1284) );
  INV_X1 U2993 ( .A(n1285), .ZN(n3699) );
  AOI22_X1 U2994 ( .A1(DATAIN[24]), .A2(n731), .B1(n737), .B2(
        \registers[24][24] ), .ZN(n1285) );
  INV_X1 U2995 ( .A(n1286), .ZN(n3700) );
  AOI22_X1 U2996 ( .A1(DATAIN[25]), .A2(n731), .B1(n738), .B2(
        \registers[24][25] ), .ZN(n1286) );
  INV_X1 U2997 ( .A(n1287), .ZN(n3701) );
  AOI22_X1 U2998 ( .A1(DATAIN[26]), .A2(n731), .B1(n738), .B2(
        \registers[24][26] ), .ZN(n1287) );
  INV_X1 U2999 ( .A(n1288), .ZN(n3702) );
  AOI22_X1 U3000 ( .A1(DATAIN[27]), .A2(n731), .B1(n738), .B2(
        \registers[24][27] ), .ZN(n1288) );
  INV_X1 U3001 ( .A(n1289), .ZN(n3703) );
  AOI22_X1 U3002 ( .A1(DATAIN[28]), .A2(n731), .B1(n738), .B2(
        \registers[24][28] ), .ZN(n1289) );
  INV_X1 U3003 ( .A(n1290), .ZN(n3704) );
  AOI22_X1 U3004 ( .A1(DATAIN[29]), .A2(n731), .B1(n738), .B2(
        \registers[24][29] ), .ZN(n1290) );
  INV_X1 U3005 ( .A(n1291), .ZN(n3705) );
  AOI22_X1 U3006 ( .A1(DATAIN[30]), .A2(n731), .B1(n739), .B2(
        \registers[24][30] ), .ZN(n1291) );
  INV_X1 U3007 ( .A(n1292), .ZN(n3706) );
  AOI22_X1 U3008 ( .A1(DATAIN[31]), .A2(n731), .B1(n739), .B2(
        \registers[24][31] ), .ZN(n1292) );
  INV_X1 U3009 ( .A(n1318), .ZN(n3666) );
  AOI22_X1 U3010 ( .A1(DATAIN[23]), .A2(n722), .B1(n728), .B2(
        \registers[23][23] ), .ZN(n1318) );
  INV_X1 U3011 ( .A(n1319), .ZN(n3667) );
  AOI22_X1 U3012 ( .A1(DATAIN[24]), .A2(n722), .B1(n728), .B2(
        \registers[23][24] ), .ZN(n1319) );
  INV_X1 U3013 ( .A(n1320), .ZN(n3668) );
  AOI22_X1 U3014 ( .A1(DATAIN[25]), .A2(n722), .B1(n729), .B2(
        \registers[23][25] ), .ZN(n1320) );
  INV_X1 U3015 ( .A(n1321), .ZN(n3669) );
  AOI22_X1 U3016 ( .A1(DATAIN[26]), .A2(n722), .B1(n729), .B2(
        \registers[23][26] ), .ZN(n1321) );
  INV_X1 U3017 ( .A(n1322), .ZN(n3670) );
  AOI22_X1 U3018 ( .A1(DATAIN[27]), .A2(n722), .B1(n729), .B2(
        \registers[23][27] ), .ZN(n1322) );
  INV_X1 U3019 ( .A(n1323), .ZN(n3671) );
  AOI22_X1 U3020 ( .A1(DATAIN[28]), .A2(n722), .B1(n729), .B2(
        \registers[23][28] ), .ZN(n1323) );
  INV_X1 U3021 ( .A(n1324), .ZN(n3672) );
  AOI22_X1 U3022 ( .A1(DATAIN[29]), .A2(n722), .B1(n729), .B2(
        \registers[23][29] ), .ZN(n1324) );
  INV_X1 U3023 ( .A(n1325), .ZN(n3673) );
  AOI22_X1 U3024 ( .A1(DATAIN[30]), .A2(n722), .B1(n730), .B2(
        \registers[23][30] ), .ZN(n1325) );
  INV_X1 U3025 ( .A(n1326), .ZN(n3674) );
  AOI22_X1 U3026 ( .A1(DATAIN[31]), .A2(n722), .B1(n730), .B2(
        \registers[23][31] ), .ZN(n1326) );
  INV_X1 U3027 ( .A(n1352), .ZN(n3634) );
  AOI22_X1 U3028 ( .A1(DATAIN[23]), .A2(n713), .B1(n719), .B2(
        \registers[22][23] ), .ZN(n1352) );
  INV_X1 U3029 ( .A(n1353), .ZN(n3635) );
  AOI22_X1 U3030 ( .A1(DATAIN[24]), .A2(n713), .B1(n719), .B2(
        \registers[22][24] ), .ZN(n1353) );
  INV_X1 U3031 ( .A(n1354), .ZN(n3636) );
  AOI22_X1 U3032 ( .A1(DATAIN[25]), .A2(n713), .B1(n720), .B2(
        \registers[22][25] ), .ZN(n1354) );
  INV_X1 U3033 ( .A(n1355), .ZN(n3637) );
  AOI22_X1 U3034 ( .A1(DATAIN[26]), .A2(n713), .B1(n720), .B2(
        \registers[22][26] ), .ZN(n1355) );
  INV_X1 U3035 ( .A(n1356), .ZN(n3638) );
  AOI22_X1 U3036 ( .A1(DATAIN[27]), .A2(n713), .B1(n720), .B2(
        \registers[22][27] ), .ZN(n1356) );
  INV_X1 U3037 ( .A(n1357), .ZN(n3639) );
  AOI22_X1 U3038 ( .A1(DATAIN[28]), .A2(n713), .B1(n720), .B2(
        \registers[22][28] ), .ZN(n1357) );
  INV_X1 U3039 ( .A(n1358), .ZN(n3640) );
  AOI22_X1 U3040 ( .A1(DATAIN[29]), .A2(n713), .B1(n720), .B2(
        \registers[22][29] ), .ZN(n1358) );
  INV_X1 U3041 ( .A(n1359), .ZN(n3641) );
  AOI22_X1 U3042 ( .A1(DATAIN[30]), .A2(n713), .B1(n721), .B2(
        \registers[22][30] ), .ZN(n1359) );
  INV_X1 U3043 ( .A(n1360), .ZN(n3642) );
  AOI22_X1 U3044 ( .A1(DATAIN[31]), .A2(n713), .B1(n721), .B2(
        \registers[22][31] ), .ZN(n1360) );
  INV_X1 U3045 ( .A(n1387), .ZN(n3602) );
  AOI22_X1 U3046 ( .A1(DATAIN[23]), .A2(n686), .B1(n692), .B2(
        \registers[19][23] ), .ZN(n1387) );
  INV_X1 U3047 ( .A(n1388), .ZN(n3603) );
  AOI22_X1 U3048 ( .A1(DATAIN[24]), .A2(n686), .B1(n692), .B2(
        \registers[19][24] ), .ZN(n1388) );
  INV_X1 U3049 ( .A(n1389), .ZN(n3604) );
  AOI22_X1 U3050 ( .A1(DATAIN[25]), .A2(n686), .B1(n693), .B2(
        \registers[19][25] ), .ZN(n1389) );
  INV_X1 U3051 ( .A(n1390), .ZN(n3605) );
  AOI22_X1 U3052 ( .A1(DATAIN[26]), .A2(n686), .B1(n693), .B2(
        \registers[19][26] ), .ZN(n1390) );
  INV_X1 U3053 ( .A(n1391), .ZN(n3606) );
  AOI22_X1 U3054 ( .A1(DATAIN[27]), .A2(n686), .B1(n693), .B2(
        \registers[19][27] ), .ZN(n1391) );
  INV_X1 U3055 ( .A(n1392), .ZN(n3607) );
  AOI22_X1 U3056 ( .A1(DATAIN[28]), .A2(n686), .B1(n693), .B2(
        \registers[19][28] ), .ZN(n1392) );
  INV_X1 U3057 ( .A(n1393), .ZN(n3608) );
  AOI22_X1 U3058 ( .A1(DATAIN[29]), .A2(n686), .B1(n693), .B2(
        \registers[19][29] ), .ZN(n1393) );
  INV_X1 U3059 ( .A(n1394), .ZN(n3609) );
  AOI22_X1 U3060 ( .A1(DATAIN[30]), .A2(n686), .B1(n694), .B2(
        \registers[19][30] ), .ZN(n1394) );
  INV_X1 U3061 ( .A(n1395), .ZN(n3610) );
  AOI22_X1 U3062 ( .A1(DATAIN[31]), .A2(n686), .B1(n694), .B2(
        \registers[19][31] ), .ZN(n1395) );
  INV_X1 U3063 ( .A(n1420), .ZN(n3570) );
  AOI22_X1 U3064 ( .A1(DATAIN[23]), .A2(n677), .B1(n683), .B2(
        \registers[18][23] ), .ZN(n1420) );
  INV_X1 U3065 ( .A(n1421), .ZN(n3571) );
  AOI22_X1 U3066 ( .A1(DATAIN[24]), .A2(n677), .B1(n683), .B2(
        \registers[18][24] ), .ZN(n1421) );
  INV_X1 U3067 ( .A(n1422), .ZN(n3572) );
  AOI22_X1 U3068 ( .A1(DATAIN[25]), .A2(n677), .B1(n684), .B2(
        \registers[18][25] ), .ZN(n1422) );
  INV_X1 U3069 ( .A(n1423), .ZN(n3573) );
  AOI22_X1 U3070 ( .A1(DATAIN[26]), .A2(n677), .B1(n684), .B2(
        \registers[18][26] ), .ZN(n1423) );
  INV_X1 U3071 ( .A(n1424), .ZN(n3574) );
  AOI22_X1 U3072 ( .A1(DATAIN[27]), .A2(n677), .B1(n684), .B2(
        \registers[18][27] ), .ZN(n1424) );
  INV_X1 U3073 ( .A(n1425), .ZN(n3575) );
  AOI22_X1 U3074 ( .A1(DATAIN[28]), .A2(n677), .B1(n684), .B2(
        \registers[18][28] ), .ZN(n1425) );
  INV_X1 U3075 ( .A(n1426), .ZN(n3576) );
  AOI22_X1 U3076 ( .A1(DATAIN[29]), .A2(n677), .B1(n684), .B2(
        \registers[18][29] ), .ZN(n1426) );
  INV_X1 U3077 ( .A(n1427), .ZN(n3577) );
  AOI22_X1 U3078 ( .A1(DATAIN[30]), .A2(n677), .B1(n685), .B2(
        \registers[18][30] ), .ZN(n1427) );
  INV_X1 U3079 ( .A(n1428), .ZN(n3578) );
  AOI22_X1 U3080 ( .A1(DATAIN[31]), .A2(n677), .B1(n685), .B2(
        \registers[18][31] ), .ZN(n1428) );
  INV_X1 U3081 ( .A(n1458), .ZN(n3441) );
  AOI22_X1 U3082 ( .A1(DATAIN[23]), .A2(n568), .B1(n574), .B2(
        \registers[13][23] ), .ZN(n1458) );
  INV_X1 U3083 ( .A(n1459), .ZN(n3442) );
  AOI22_X1 U3084 ( .A1(DATAIN[24]), .A2(n568), .B1(n574), .B2(
        \registers[13][24] ), .ZN(n1459) );
  INV_X1 U3085 ( .A(n1460), .ZN(n3443) );
  AOI22_X1 U3086 ( .A1(DATAIN[25]), .A2(n568), .B1(n575), .B2(
        \registers[13][25] ), .ZN(n1460) );
  INV_X1 U3087 ( .A(n1461), .ZN(n3444) );
  AOI22_X1 U3088 ( .A1(DATAIN[26]), .A2(n568), .B1(n575), .B2(
        \registers[13][26] ), .ZN(n1461) );
  INV_X1 U3089 ( .A(n1462), .ZN(n3445) );
  AOI22_X1 U3090 ( .A1(DATAIN[27]), .A2(n568), .B1(n575), .B2(
        \registers[13][27] ), .ZN(n1462) );
  INV_X1 U3091 ( .A(n1463), .ZN(n3446) );
  AOI22_X1 U3092 ( .A1(DATAIN[28]), .A2(n568), .B1(n575), .B2(
        \registers[13][28] ), .ZN(n1463) );
  INV_X1 U3093 ( .A(n1464), .ZN(n3447) );
  AOI22_X1 U3094 ( .A1(DATAIN[29]), .A2(n568), .B1(n575), .B2(
        \registers[13][29] ), .ZN(n1464) );
  INV_X1 U3095 ( .A(n1465), .ZN(n3448) );
  AOI22_X1 U3096 ( .A1(DATAIN[30]), .A2(n568), .B1(n576), .B2(
        \registers[13][30] ), .ZN(n1465) );
  INV_X1 U3097 ( .A(n1466), .ZN(n3449) );
  AOI22_X1 U3098 ( .A1(DATAIN[31]), .A2(n568), .B1(n576), .B2(
        \registers[13][31] ), .ZN(n1466) );
  INV_X1 U3099 ( .A(n1491), .ZN(n3409) );
  AOI22_X1 U3100 ( .A1(DATAIN[23]), .A2(n559), .B1(n565), .B2(
        \registers[12][23] ), .ZN(n1491) );
  INV_X1 U3101 ( .A(n1492), .ZN(n3410) );
  AOI22_X1 U3102 ( .A1(DATAIN[24]), .A2(n559), .B1(n565), .B2(
        \registers[12][24] ), .ZN(n1492) );
  INV_X1 U3103 ( .A(n1493), .ZN(n3411) );
  AOI22_X1 U3104 ( .A1(DATAIN[25]), .A2(n559), .B1(n566), .B2(
        \registers[12][25] ), .ZN(n1493) );
  INV_X1 U3105 ( .A(n1494), .ZN(n3412) );
  AOI22_X1 U3106 ( .A1(DATAIN[26]), .A2(n559), .B1(n566), .B2(
        \registers[12][26] ), .ZN(n1494) );
  INV_X1 U3107 ( .A(n1495), .ZN(n3413) );
  AOI22_X1 U3108 ( .A1(DATAIN[27]), .A2(n559), .B1(n566), .B2(
        \registers[12][27] ), .ZN(n1495) );
  INV_X1 U3109 ( .A(n1496), .ZN(n3414) );
  AOI22_X1 U3110 ( .A1(DATAIN[28]), .A2(n559), .B1(n566), .B2(
        \registers[12][28] ), .ZN(n1496) );
  INV_X1 U3111 ( .A(n1497), .ZN(n3415) );
  AOI22_X1 U3112 ( .A1(DATAIN[29]), .A2(n559), .B1(n566), .B2(
        \registers[12][29] ), .ZN(n1497) );
  INV_X1 U3113 ( .A(n1498), .ZN(n3416) );
  AOI22_X1 U3114 ( .A1(DATAIN[30]), .A2(n559), .B1(n567), .B2(
        \registers[12][30] ), .ZN(n1498) );
  INV_X1 U3115 ( .A(n1499), .ZN(n3417) );
  AOI22_X1 U3116 ( .A1(DATAIN[31]), .A2(n559), .B1(n567), .B2(
        \registers[12][31] ), .ZN(n1499) );
  INV_X1 U3117 ( .A(n1526), .ZN(n3377) );
  AOI22_X1 U3118 ( .A1(DATAIN[23]), .A2(n404), .B1(n410), .B2(
        \registers[9][23] ), .ZN(n1526) );
  INV_X1 U3119 ( .A(n1527), .ZN(n3378) );
  AOI22_X1 U3120 ( .A1(DATAIN[24]), .A2(n404), .B1(n410), .B2(
        \registers[9][24] ), .ZN(n1527) );
  INV_X1 U3121 ( .A(n1528), .ZN(n3379) );
  AOI22_X1 U3122 ( .A1(DATAIN[25]), .A2(n404), .B1(n411), .B2(
        \registers[9][25] ), .ZN(n1528) );
  INV_X1 U3123 ( .A(n1529), .ZN(n3380) );
  AOI22_X1 U3124 ( .A1(DATAIN[26]), .A2(n404), .B1(n411), .B2(
        \registers[9][26] ), .ZN(n1529) );
  INV_X1 U3125 ( .A(n1530), .ZN(n3381) );
  AOI22_X1 U3126 ( .A1(DATAIN[27]), .A2(n404), .B1(n411), .B2(
        \registers[9][27] ), .ZN(n1530) );
  INV_X1 U3127 ( .A(n1531), .ZN(n3382) );
  AOI22_X1 U3128 ( .A1(DATAIN[28]), .A2(n404), .B1(n411), .B2(
        \registers[9][28] ), .ZN(n1531) );
  INV_X1 U3129 ( .A(n1532), .ZN(n3383) );
  AOI22_X1 U3130 ( .A1(DATAIN[29]), .A2(n404), .B1(n411), .B2(
        \registers[9][29] ), .ZN(n1532) );
  INV_X1 U3131 ( .A(n1533), .ZN(n3384) );
  AOI22_X1 U3132 ( .A1(DATAIN[30]), .A2(n404), .B1(n412), .B2(
        \registers[9][30] ), .ZN(n1533) );
  INV_X1 U3133 ( .A(n1534), .ZN(n3385) );
  AOI22_X1 U3134 ( .A1(DATAIN[31]), .A2(n404), .B1(n412), .B2(
        \registers[9][31] ), .ZN(n1534) );
  INV_X1 U3135 ( .A(n1559), .ZN(n3345) );
  AOI22_X1 U3136 ( .A1(DATAIN[23]), .A2(n395), .B1(n401), .B2(
        \registers[8][23] ), .ZN(n1559) );
  INV_X1 U3137 ( .A(n1560), .ZN(n3346) );
  AOI22_X1 U3138 ( .A1(DATAIN[24]), .A2(n395), .B1(n401), .B2(
        \registers[8][24] ), .ZN(n1560) );
  INV_X1 U3139 ( .A(n1561), .ZN(n3347) );
  AOI22_X1 U3140 ( .A1(DATAIN[25]), .A2(n395), .B1(n402), .B2(
        \registers[8][25] ), .ZN(n1561) );
  INV_X1 U3141 ( .A(n1562), .ZN(n3348) );
  AOI22_X1 U3142 ( .A1(DATAIN[26]), .A2(n395), .B1(n402), .B2(
        \registers[8][26] ), .ZN(n1562) );
  INV_X1 U3143 ( .A(n1563), .ZN(n3349) );
  AOI22_X1 U3144 ( .A1(DATAIN[27]), .A2(n395), .B1(n402), .B2(
        \registers[8][27] ), .ZN(n1563) );
  INV_X1 U3145 ( .A(n1564), .ZN(n3350) );
  AOI22_X1 U3146 ( .A1(DATAIN[28]), .A2(n395), .B1(n402), .B2(
        \registers[8][28] ), .ZN(n1564) );
  INV_X1 U3147 ( .A(n1565), .ZN(n3351) );
  AOI22_X1 U3148 ( .A1(DATAIN[29]), .A2(n395), .B1(n402), .B2(
        \registers[8][29] ), .ZN(n1565) );
  INV_X1 U3149 ( .A(n1566), .ZN(n3352) );
  AOI22_X1 U3150 ( .A1(DATAIN[30]), .A2(n395), .B1(n403), .B2(
        \registers[8][30] ), .ZN(n1566) );
  INV_X1 U3151 ( .A(n1567), .ZN(n3353) );
  AOI22_X1 U3152 ( .A1(DATAIN[31]), .A2(n395), .B1(n403), .B2(
        \registers[8][31] ), .ZN(n1567) );
  INV_X1 U3153 ( .A(n1101), .ZN(n3537) );
  AOI22_X1 U3154 ( .A1(DATAIN[23]), .A2(n912), .B1(n918), .B2(
        \registers[6][23] ), .ZN(n1101) );
  INV_X1 U3155 ( .A(n1102), .ZN(n3538) );
  AOI22_X1 U3156 ( .A1(DATAIN[24]), .A2(n912), .B1(n918), .B2(
        \registers[6][24] ), .ZN(n1102) );
  INV_X1 U3157 ( .A(n1103), .ZN(n3539) );
  AOI22_X1 U3158 ( .A1(DATAIN[25]), .A2(n912), .B1(n919), .B2(
        \registers[6][25] ), .ZN(n1103) );
  INV_X1 U3159 ( .A(n1104), .ZN(n3540) );
  AOI22_X1 U3160 ( .A1(DATAIN[26]), .A2(n912), .B1(n919), .B2(
        \registers[6][26] ), .ZN(n1104) );
  INV_X1 U3161 ( .A(n1105), .ZN(n3541) );
  AOI22_X1 U3162 ( .A1(DATAIN[27]), .A2(n912), .B1(n919), .B2(
        \registers[6][27] ), .ZN(n1105) );
  INV_X1 U3163 ( .A(n1106), .ZN(n3542) );
  AOI22_X1 U3164 ( .A1(DATAIN[28]), .A2(n912), .B1(n919), .B2(
        \registers[6][28] ), .ZN(n1106) );
  INV_X1 U3165 ( .A(n1107), .ZN(n3543) );
  AOI22_X1 U3166 ( .A1(DATAIN[29]), .A2(n912), .B1(n919), .B2(
        \registers[6][29] ), .ZN(n1107) );
  INV_X1 U3167 ( .A(n1108), .ZN(n3544) );
  AOI22_X1 U3168 ( .A1(DATAIN[30]), .A2(n912), .B1(n920), .B2(
        \registers[6][30] ), .ZN(n1108) );
  INV_X1 U3169 ( .A(n1109), .ZN(n3545) );
  AOI22_X1 U3170 ( .A1(DATAIN[31]), .A2(n912), .B1(n920), .B2(
        \registers[6][31] ), .ZN(n1109) );
  INV_X1 U3171 ( .A(n1144), .ZN(n3505) );
  AOI22_X1 U3172 ( .A1(DATAIN[23]), .A2(n867), .B1(n873), .B2(
        \registers[1][23] ), .ZN(n1144) );
  INV_X1 U3173 ( .A(n1145), .ZN(n3506) );
  AOI22_X1 U3174 ( .A1(DATAIN[24]), .A2(n867), .B1(n873), .B2(
        \registers[1][24] ), .ZN(n1145) );
  INV_X1 U3175 ( .A(n1146), .ZN(n3507) );
  AOI22_X1 U3176 ( .A1(DATAIN[25]), .A2(n867), .B1(n874), .B2(
        \registers[1][25] ), .ZN(n1146) );
  INV_X1 U3177 ( .A(n1147), .ZN(n3508) );
  AOI22_X1 U3178 ( .A1(DATAIN[26]), .A2(n867), .B1(n874), .B2(
        \registers[1][26] ), .ZN(n1147) );
  INV_X1 U3179 ( .A(n1148), .ZN(n3509) );
  AOI22_X1 U3180 ( .A1(DATAIN[27]), .A2(n867), .B1(n874), .B2(
        \registers[1][27] ), .ZN(n1148) );
  INV_X1 U3181 ( .A(n1149), .ZN(n3510) );
  AOI22_X1 U3182 ( .A1(DATAIN[28]), .A2(n867), .B1(n874), .B2(
        \registers[1][28] ), .ZN(n1149) );
  INV_X1 U3183 ( .A(n1150), .ZN(n3511) );
  AOI22_X1 U3184 ( .A1(DATAIN[29]), .A2(n867), .B1(n874), .B2(
        \registers[1][29] ), .ZN(n1150) );
  INV_X1 U3185 ( .A(n1151), .ZN(n3512) );
  AOI22_X1 U3186 ( .A1(DATAIN[30]), .A2(n867), .B1(n875), .B2(
        \registers[1][30] ), .ZN(n1151) );
  INV_X1 U3187 ( .A(n1152), .ZN(n3513) );
  AOI22_X1 U3188 ( .A1(DATAIN[31]), .A2(n867), .B1(n875), .B2(
        \registers[1][31] ), .ZN(n1152) );
  INV_X1 U3189 ( .A(n1077), .ZN(n3514) );
  AOI22_X1 U3190 ( .A1(n913), .A2(DATAIN[0]), .B1(n914), .B2(\registers[6][0] ), .ZN(n1077) );
  INV_X1 U3191 ( .A(n1079), .ZN(n3515) );
  AOI22_X1 U3192 ( .A1(n912), .A2(DATAIN[1]), .B1(n914), .B2(\registers[6][1] ), .ZN(n1079) );
  INV_X1 U3193 ( .A(n1080), .ZN(n3516) );
  AOI22_X1 U3194 ( .A1(n913), .A2(DATAIN[2]), .B1(n914), .B2(\registers[6][2] ), .ZN(n1080) );
  INV_X1 U3195 ( .A(n1081), .ZN(n3517) );
  AOI22_X1 U3196 ( .A1(n912), .A2(DATAIN[3]), .B1(n914), .B2(\registers[6][3] ), .ZN(n1081) );
  INV_X1 U3197 ( .A(n1082), .ZN(n3518) );
  AOI22_X1 U3198 ( .A1(n913), .A2(DATAIN[4]), .B1(n914), .B2(\registers[6][4] ), .ZN(n1082) );
  INV_X1 U3199 ( .A(n1083), .ZN(n3519) );
  AOI22_X1 U3200 ( .A1(n912), .A2(DATAIN[5]), .B1(n915), .B2(\registers[6][5] ), .ZN(n1083) );
  INV_X1 U3201 ( .A(n1084), .ZN(n3520) );
  AOI22_X1 U3202 ( .A1(n913), .A2(DATAIN[6]), .B1(n915), .B2(\registers[6][6] ), .ZN(n1084) );
  INV_X1 U3203 ( .A(n1085), .ZN(n3521) );
  AOI22_X1 U3204 ( .A1(n912), .A2(DATAIN[7]), .B1(n915), .B2(\registers[6][7] ), .ZN(n1085) );
  INV_X1 U3205 ( .A(n1098), .ZN(n3534) );
  AOI22_X1 U3206 ( .A1(n912), .A2(DATAIN[20]), .B1(n918), .B2(
        \registers[6][20] ), .ZN(n1098) );
  INV_X1 U3207 ( .A(n1099), .ZN(n3535) );
  AOI22_X1 U3208 ( .A1(n912), .A2(DATAIN[21]), .B1(n918), .B2(
        \registers[6][21] ), .ZN(n1099) );
  INV_X1 U3209 ( .A(n1100), .ZN(n3536) );
  AOI22_X1 U3210 ( .A1(n912), .A2(DATAIN[22]), .B1(n918), .B2(
        \registers[6][22] ), .ZN(n1100) );
  INV_X1 U3211 ( .A(n1086), .ZN(n3522) );
  AOI22_X1 U3212 ( .A1(n913), .A2(DATAIN[8]), .B1(n915), .B2(\registers[6][8] ), .ZN(n1086) );
  INV_X1 U3213 ( .A(n1087), .ZN(n3523) );
  AOI22_X1 U3214 ( .A1(n913), .A2(DATAIN[9]), .B1(n915), .B2(\registers[6][9] ), .ZN(n1087) );
  INV_X1 U3215 ( .A(n1088), .ZN(n3524) );
  AOI22_X1 U3216 ( .A1(n913), .A2(DATAIN[10]), .B1(n916), .B2(
        \registers[6][10] ), .ZN(n1088) );
  INV_X1 U3217 ( .A(n1089), .ZN(n3525) );
  AOI22_X1 U3218 ( .A1(n913), .A2(DATAIN[11]), .B1(n916), .B2(
        \registers[6][11] ), .ZN(n1089) );
  INV_X1 U3219 ( .A(n1090), .ZN(n3526) );
  AOI22_X1 U3220 ( .A1(n913), .A2(DATAIN[12]), .B1(n916), .B2(
        \registers[6][12] ), .ZN(n1090) );
  INV_X1 U3221 ( .A(n1091), .ZN(n3527) );
  AOI22_X1 U3222 ( .A1(n913), .A2(DATAIN[13]), .B1(n916), .B2(
        \registers[6][13] ), .ZN(n1091) );
  INV_X1 U3223 ( .A(n1092), .ZN(n3528) );
  AOI22_X1 U3224 ( .A1(n913), .A2(DATAIN[14]), .B1(n916), .B2(
        \registers[6][14] ), .ZN(n1092) );
  INV_X1 U3225 ( .A(n1093), .ZN(n3529) );
  AOI22_X1 U3226 ( .A1(n913), .A2(DATAIN[15]), .B1(n917), .B2(
        \registers[6][15] ), .ZN(n1093) );
  INV_X1 U3227 ( .A(n1094), .ZN(n3530) );
  AOI22_X1 U3228 ( .A1(n913), .A2(DATAIN[16]), .B1(n917), .B2(
        \registers[6][16] ), .ZN(n1094) );
  INV_X1 U3229 ( .A(n1095), .ZN(n3531) );
  AOI22_X1 U3230 ( .A1(n913), .A2(DATAIN[17]), .B1(n917), .B2(
        \registers[6][17] ), .ZN(n1095) );
  INV_X1 U3231 ( .A(n1096), .ZN(n3532) );
  AOI22_X1 U3232 ( .A1(n913), .A2(DATAIN[18]), .B1(n917), .B2(
        \registers[6][18] ), .ZN(n1096) );
  INV_X1 U3233 ( .A(n1097), .ZN(n3533) );
  AOI22_X1 U3234 ( .A1(n913), .A2(DATAIN[19]), .B1(n917), .B2(
        \registers[6][19] ), .ZN(n1097) );
  INV_X1 U3235 ( .A(n1569), .ZN(n3460) );
  AOI22_X1 U3236 ( .A1(n922), .A2(DATAIN[1]), .B1(n925), .B2(\registers[7][1] ), .ZN(n1569) );
  INV_X1 U3237 ( .A(n1570), .ZN(n3461) );
  AOI22_X1 U3238 ( .A1(n922), .A2(DATAIN[2]), .B1(n925), .B2(\registers[7][2] ), .ZN(n1570) );
  INV_X1 U3239 ( .A(n1571), .ZN(n3462) );
  AOI22_X1 U3240 ( .A1(n922), .A2(DATAIN[3]), .B1(n925), .B2(\registers[7][3] ), .ZN(n1571) );
  INV_X1 U3241 ( .A(n1572), .ZN(n3463) );
  AOI22_X1 U3242 ( .A1(n922), .A2(DATAIN[4]), .B1(n925), .B2(\registers[7][4] ), .ZN(n1572) );
  INV_X1 U3243 ( .A(n1573), .ZN(n3464) );
  AOI22_X1 U3244 ( .A1(n922), .A2(DATAIN[5]), .B1(n925), .B2(\registers[7][5] ), .ZN(n1573) );
  INV_X1 U3245 ( .A(n1574), .ZN(n3465) );
  AOI22_X1 U3246 ( .A1(n922), .A2(DATAIN[6]), .B1(n926), .B2(\registers[7][6] ), .ZN(n1574) );
  INV_X1 U3247 ( .A(n1575), .ZN(n3466) );
  AOI22_X1 U3248 ( .A1(n922), .A2(DATAIN[7]), .B1(n926), .B2(\registers[7][7] ), .ZN(n1575) );
  INV_X1 U3249 ( .A(n1576), .ZN(n3467) );
  AOI22_X1 U3250 ( .A1(n922), .A2(DATAIN[8]), .B1(n926), .B2(\registers[7][8] ), .ZN(n1576) );
  INV_X1 U3251 ( .A(n1577), .ZN(n3468) );
  AOI22_X1 U3252 ( .A1(n922), .A2(DATAIN[9]), .B1(n926), .B2(\registers[7][9] ), .ZN(n1577) );
  INV_X1 U3253 ( .A(n1578), .ZN(n3469) );
  AOI22_X1 U3254 ( .A1(n922), .A2(DATAIN[10]), .B1(n926), .B2(
        \registers[7][10] ), .ZN(n1578) );
  INV_X1 U3255 ( .A(n1579), .ZN(n3470) );
  AOI22_X1 U3256 ( .A1(n922), .A2(DATAIN[11]), .B1(n927), .B2(
        \registers[7][11] ), .ZN(n1579) );
  INV_X1 U3257 ( .A(n1580), .ZN(n3471) );
  AOI22_X1 U3258 ( .A1(n921), .A2(DATAIN[12]), .B1(n927), .B2(
        \registers[7][12] ), .ZN(n1580) );
  INV_X1 U3259 ( .A(n1581), .ZN(n3472) );
  AOI22_X1 U3260 ( .A1(n921), .A2(DATAIN[13]), .B1(n927), .B2(
        \registers[7][13] ), .ZN(n1581) );
  INV_X1 U3261 ( .A(n1582), .ZN(n3473) );
  AOI22_X1 U3262 ( .A1(n921), .A2(DATAIN[14]), .B1(n927), .B2(
        \registers[7][14] ), .ZN(n1582) );
  INV_X1 U3263 ( .A(n1583), .ZN(n3474) );
  AOI22_X1 U3264 ( .A1(n921), .A2(DATAIN[15]), .B1(n927), .B2(
        \registers[7][15] ), .ZN(n1583) );
  INV_X1 U3265 ( .A(n1584), .ZN(n3475) );
  AOI22_X1 U3266 ( .A1(n921), .A2(DATAIN[16]), .B1(n928), .B2(
        \registers[7][16] ), .ZN(n1584) );
  INV_X1 U3267 ( .A(n1585), .ZN(n3476) );
  AOI22_X1 U3268 ( .A1(n921), .A2(DATAIN[17]), .B1(n928), .B2(
        \registers[7][17] ), .ZN(n1585) );
  INV_X1 U3269 ( .A(n1586), .ZN(n3477) );
  AOI22_X1 U3270 ( .A1(n921), .A2(DATAIN[18]), .B1(n928), .B2(
        \registers[7][18] ), .ZN(n1586) );
  INV_X1 U3271 ( .A(n1587), .ZN(n3478) );
  AOI22_X1 U3272 ( .A1(n921), .A2(DATAIN[19]), .B1(n928), .B2(
        \registers[7][19] ), .ZN(n1587) );
  INV_X1 U3273 ( .A(n1588), .ZN(n3479) );
  AOI22_X1 U3274 ( .A1(n921), .A2(DATAIN[20]), .B1(n928), .B2(
        \registers[7][20] ), .ZN(n1588) );
  INV_X1 U3275 ( .A(n1589), .ZN(n3480) );
  AOI22_X1 U3276 ( .A1(n921), .A2(DATAIN[21]), .B1(n993), .B2(
        \registers[7][21] ), .ZN(n1589) );
  INV_X1 U3277 ( .A(n1590), .ZN(n3481) );
  AOI22_X1 U3278 ( .A1(n921), .A2(DATAIN[22]), .B1(n993), .B2(
        \registers[7][22] ), .ZN(n1590) );
  INV_X1 U3279 ( .A(n1568), .ZN(n3459) );
  AOI22_X1 U3280 ( .A1(n922), .A2(DATAIN[0]), .B1(n924), .B2(\registers[7][0] ), .ZN(n1568) );
  INV_X1 U3281 ( .A(n1067), .ZN(n3450) );
  AOI22_X1 U3282 ( .A1(n921), .A2(DATAIN[23]), .B1(n923), .B2(
        \registers[7][23] ), .ZN(n1067) );
  INV_X1 U3283 ( .A(n1069), .ZN(n3451) );
  AOI22_X1 U3284 ( .A1(n922), .A2(DATAIN[24]), .B1(n923), .B2(
        \registers[7][24] ), .ZN(n1069) );
  INV_X1 U3285 ( .A(n1070), .ZN(n3452) );
  AOI22_X1 U3286 ( .A1(n921), .A2(DATAIN[25]), .B1(n923), .B2(
        \registers[7][25] ), .ZN(n1070) );
  INV_X1 U3287 ( .A(n1071), .ZN(n3453) );
  AOI22_X1 U3288 ( .A1(n922), .A2(DATAIN[26]), .B1(n923), .B2(
        \registers[7][26] ), .ZN(n1071) );
  INV_X1 U3289 ( .A(n1072), .ZN(n3454) );
  AOI22_X1 U3290 ( .A1(n921), .A2(DATAIN[27]), .B1(n923), .B2(
        \registers[7][27] ), .ZN(n1072) );
  INV_X1 U3291 ( .A(n1073), .ZN(n3455) );
  AOI22_X1 U3292 ( .A1(n922), .A2(DATAIN[28]), .B1(n924), .B2(
        \registers[7][28] ), .ZN(n1073) );
  INV_X1 U3293 ( .A(n1074), .ZN(n3456) );
  AOI22_X1 U3294 ( .A1(n921), .A2(DATAIN[29]), .B1(n924), .B2(
        \registers[7][29] ), .ZN(n1074) );
  INV_X1 U3295 ( .A(n1075), .ZN(n3457) );
  AOI22_X1 U3296 ( .A1(n922), .A2(DATAIN[30]), .B1(n924), .B2(
        \registers[7][30] ), .ZN(n1075) );
  INV_X1 U3297 ( .A(n1076), .ZN(n3458) );
  AOI22_X1 U3298 ( .A1(n921), .A2(DATAIN[31]), .B1(n924), .B2(
        \registers[7][31] ), .ZN(n1076) );
  AND2_X1 U3299 ( .A1(RD2), .A2(ENABLE), .ZN(N217) );
  AND2_X1 U3300 ( .A1(RD1), .A2(ENABLE), .ZN(N82) );
  CLKBUF_X1 U3301 ( .A(N217), .Z(n994) );
  CLKBUF_X1 U3302 ( .A(N217), .Z(n995) );
  CLKBUF_X1 U3303 ( .A(N217), .Z(n996) );
  CLKBUF_X1 U3304 ( .A(N217), .Z(n997) );
  CLKBUF_X1 U3305 ( .A(N82), .Z(n998) );
  CLKBUF_X1 U3306 ( .A(N82), .Z(n999) );
  CLKBUF_X1 U3307 ( .A(N82), .Z(n1000) );
  CLKBUF_X1 U3308 ( .A(N82), .Z(n1001) );
  CLKBUF_X1 U3309 ( .A(n3321), .Z(n1013) );
  CLKBUF_X1 U3310 ( .A(n3320), .Z(n1014) );
  CLKBUF_X1 U3311 ( .A(n3320), .Z(n1015) );
  CLKBUF_X1 U3312 ( .A(n3320), .Z(n1016) );
  CLKBUF_X1 U3313 ( .A(n3320), .Z(n1017) );
  CLKBUF_X1 U3314 ( .A(n3320), .Z(n1018) );
  CLKBUF_X1 U3315 ( .A(n3320), .Z(n1019) );
  CLKBUF_X1 U3316 ( .A(n3319), .Z(n1020) );
  CLKBUF_X1 U3317 ( .A(n3319), .Z(n1021) );
  CLKBUF_X1 U3318 ( .A(n3319), .Z(n1022) );
  CLKBUF_X1 U3319 ( .A(n3319), .Z(n1023) );
  CLKBUF_X1 U3320 ( .A(n3319), .Z(n1024) );
  CLKBUF_X1 U3321 ( .A(n3319), .Z(n1025) );
  CLKBUF_X1 U3322 ( .A(n3318), .Z(n1026) );
  CLKBUF_X1 U3323 ( .A(n3318), .Z(n1027) );
  CLKBUF_X1 U3324 ( .A(n3318), .Z(n1028) );
  CLKBUF_X1 U3325 ( .A(n3318), .Z(n1029) );
  CLKBUF_X1 U3326 ( .A(n3318), .Z(n1030) );
  CLKBUF_X1 U3327 ( .A(n3318), .Z(n1031) );
  CLKBUF_X1 U3328 ( .A(n3317), .Z(n1032) );
  CLKBUF_X1 U3329 ( .A(n3317), .Z(n1033) );
  CLKBUF_X1 U3330 ( .A(n3317), .Z(n1034) );
  CLKBUF_X1 U3331 ( .A(n3317), .Z(n1035) );
  CLKBUF_X1 U3332 ( .A(n3317), .Z(n1036) );
  CLKBUF_X1 U3333 ( .A(n3317), .Z(n1037) );
  CLKBUF_X1 U3334 ( .A(n3316), .Z(n1038) );
  CLKBUF_X1 U3335 ( .A(n3316), .Z(n1039) );
  CLKBUF_X1 U3336 ( .A(n3316), .Z(n1040) );
  CLKBUF_X1 U3337 ( .A(n3316), .Z(n1041) );
  CLKBUF_X1 U3338 ( .A(n3316), .Z(n1042) );
  CLKBUF_X1 U3339 ( .A(n3316), .Z(n1043) );
  CLKBUF_X1 U3340 ( .A(n3315), .Z(n1044) );
  CLKBUF_X1 U3341 ( .A(n3315), .Z(n1045) );
  CLKBUF_X1 U3342 ( .A(n3315), .Z(n1046) );
  CLKBUF_X1 U3343 ( .A(n3315), .Z(n1047) );
  CLKBUF_X1 U3344 ( .A(n3315), .Z(n1048) );
  CLKBUF_X1 U3345 ( .A(n3315), .Z(n1049) );
  CLKBUF_X1 U3346 ( .A(n3314), .Z(n1050) );
  CLKBUF_X1 U3347 ( .A(n3314), .Z(n1051) );
  CLKBUF_X1 U3348 ( .A(n3314), .Z(n1052) );
  CLKBUF_X1 U3349 ( .A(n3314), .Z(n1053) );
  CLKBUF_X1 U3350 ( .A(n3314), .Z(n1054) );
  CLKBUF_X1 U3351 ( .A(n3314), .Z(n1055) );
  CLKBUF_X1 U3352 ( .A(n3313), .Z(n1056) );
  CLKBUF_X1 U3353 ( .A(n3313), .Z(n1057) );
  CLKBUF_X1 U3354 ( .A(n3313), .Z(n1058) );
  CLKBUF_X1 U3355 ( .A(n3313), .Z(n1059) );
  CLKBUF_X1 U3356 ( .A(n3313), .Z(n1060) );
  CLKBUF_X1 U3357 ( .A(n3313), .Z(n1061) );
  CLKBUF_X1 U3358 ( .A(n3312), .Z(n1062) );
  CLKBUF_X1 U3359 ( .A(n3312), .Z(n1063) );
  CLKBUF_X1 U3360 ( .A(n3312), .Z(n1064) );
  CLKBUF_X1 U3361 ( .A(n3312), .Z(n1065) );
  CLKBUF_X1 U3362 ( .A(n3312), .Z(n1066) );
  CLKBUF_X1 U3363 ( .A(n3312), .Z(n1112) );
  CLKBUF_X1 U3364 ( .A(n3311), .Z(n1114) );
  CLKBUF_X1 U3365 ( .A(n3311), .Z(n1116) );
  CLKBUF_X1 U3366 ( .A(n3311), .Z(n1118) );
  CLKBUF_X1 U3367 ( .A(n3311), .Z(n1155) );
  CLKBUF_X1 U3368 ( .A(n3311), .Z(n1158) );
  CLKBUF_X1 U3369 ( .A(n3311), .Z(n1225) );
  CLKBUF_X1 U3370 ( .A(n3310), .Z(n1226) );
  CLKBUF_X1 U3371 ( .A(n3310), .Z(n1361) );
  CLKBUF_X1 U3372 ( .A(n3310), .Z(n1362) );
  CLKBUF_X1 U3373 ( .A(n3310), .Z(n1429) );
  CLKBUF_X1 U3374 ( .A(n3310), .Z(n1430) );
  CLKBUF_X1 U3375 ( .A(n3310), .Z(n1431) );
  CLKBUF_X1 U3376 ( .A(n3309), .Z(n1433) );
  CLKBUF_X1 U3377 ( .A(n3309), .Z(n1500) );
  CLKBUF_X1 U3378 ( .A(n3309), .Z(n1501) );
  CLKBUF_X1 U3379 ( .A(n3309), .Z(n3285) );
  CLKBUF_X1 U3380 ( .A(n3309), .Z(n3286) );
  CLKBUF_X1 U3381 ( .A(n3309), .Z(n3287) );
  CLKBUF_X1 U3382 ( .A(n3308), .Z(n3288) );
  CLKBUF_X1 U3383 ( .A(n3308), .Z(n3289) );
  CLKBUF_X1 U3384 ( .A(n3308), .Z(n3290) );
  CLKBUF_X1 U3385 ( .A(n3308), .Z(n3291) );
  CLKBUF_X1 U3386 ( .A(n3308), .Z(n3292) );
  CLKBUF_X1 U3387 ( .A(n3308), .Z(n3293) );
  CLKBUF_X1 U3388 ( .A(n3307), .Z(n3294) );
  CLKBUF_X1 U3389 ( .A(n3307), .Z(n3295) );
  CLKBUF_X1 U3390 ( .A(n3307), .Z(n3296) );
  CLKBUF_X1 U3391 ( .A(n3307), .Z(n3297) );
  CLKBUF_X1 U3392 ( .A(n3307), .Z(n3298) );
  CLKBUF_X1 U3393 ( .A(n3307), .Z(n3299) );
  CLKBUF_X1 U3394 ( .A(n3306), .Z(n3300) );
  CLKBUF_X1 U3395 ( .A(n3306), .Z(n3301) );
  CLKBUF_X1 U3396 ( .A(n3306), .Z(n3302) );
  CLKBUF_X1 U3397 ( .A(n3306), .Z(n3303) );
  CLKBUF_X1 U3398 ( .A(n3306), .Z(n3304) );
  CLKBUF_X1 U3399 ( .A(n3306), .Z(n3305) );
endmodule


module REG_PIPO_6_00_00_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n27), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n26), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n25), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n24), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n22), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n28), .ZN(n20) );
  INV_X1 U3 ( .A(n21), .ZN(n22) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n20), .B1(n28), .B2(DOUT[0]), .ZN(n21) );
  INV_X1 U5 ( .A(n19), .ZN(n23) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n20), .B1(n28), .B2(DOUT[1]), .ZN(n19) );
  INV_X1 U7 ( .A(n18), .ZN(n24) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n20), .B1(n28), .B2(DOUT[2]), .ZN(n18) );
  INV_X1 U9 ( .A(n17), .ZN(n25) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n20), .B1(n28), .B2(DOUT[3]), .ZN(n17) );
  INV_X1 U11 ( .A(n16), .ZN(n26) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n20), .B1(n28), .B2(DOUT[4]), .ZN(n16) );
  INV_X1 U13 ( .A(n15), .ZN(n27) );
  AOI22_X1 U14 ( .A1(DIN[5]), .A2(n20), .B1(n28), .B2(DOUT[5]), .ZN(n15) );
  INV_X1 U15 ( .A(EN), .ZN(n28) );
endmodule


module REG_PIPO_32_00000000_00000000_21 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_32_00000000_00000000_20 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_32_00000000_00000000_19 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_32_00000000_00000000_18 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n177), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n177) );
  OAI22_X1 U60 ( .A1(n239), .A2(EN), .B1(n170), .B2(n181), .ZN(n271) );
  INV_X1 U61 ( .A(DIN[29]), .ZN(n181) );
  OAI22_X1 U62 ( .A1(n236), .A2(EN), .B1(n170), .B2(n178), .ZN(n268) );
  INV_X1 U63 ( .A(DIN[26]), .ZN(n178) );
  OAI22_X1 U64 ( .A1(n237), .A2(EN), .B1(n170), .B2(n179), .ZN(n269) );
  INV_X1 U65 ( .A(DIN[27]), .ZN(n179) );
  OAI22_X1 U66 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U67 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n182), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n182) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n183), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n183) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_5_00_00_7 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n22), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n21), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n20), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n19), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n24), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(n19) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n17), .B1(n24), .B2(DOUT[0]), .ZN(n18) );
  INV_X1 U5 ( .A(n16), .ZN(n20) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n17), .B1(n24), .B2(DOUT[1]), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(n21) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n17), .B1(n24), .B2(DOUT[2]), .ZN(n15) );
  INV_X1 U9 ( .A(n14), .ZN(n22) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n17), .B1(n24), .B2(DOUT[3]), .ZN(n14) );
  INV_X1 U11 ( .A(n13), .ZN(n23) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n17), .B1(n24), .B2(DOUT[4]), .ZN(n13) );
  INV_X1 U13 ( .A(EN), .ZN(n24) );
endmodule


module REG_PIPO_5_00_00_6 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n19), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n20), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n21), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n22), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n24), .ZN(n26) );
  INV_X1 U3 ( .A(n25), .ZN(n23) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n26), .B1(n24), .B2(DOUT[0]), .ZN(n25) );
  INV_X1 U5 ( .A(n27), .ZN(n22) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n26), .B1(n24), .B2(DOUT[1]), .ZN(n27) );
  INV_X1 U7 ( .A(n28), .ZN(n21) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n26), .B1(n24), .B2(DOUT[2]), .ZN(n28) );
  INV_X1 U9 ( .A(n29), .ZN(n20) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n26), .B1(n24), .B2(DOUT[3]), .ZN(n29) );
  INV_X1 U11 ( .A(n30), .ZN(n19) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n26), .B1(n24), .B2(DOUT[4]), .ZN(n30) );
  INV_X1 U13 ( .A(EN), .ZN(n24) );
endmodule


module PG_PRIM_32 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GG_37 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   net24009, n1, n2;
  assign G = net24009;

  NOR2_X1 U1 ( .A1(G_CURRENT), .A2(G_PREV), .ZN(n1) );
  NOR2_X1 U2 ( .A1(n2), .A2(n1), .ZN(net24009) );
  NOR2_X1 U3 ( .A1(P_CURRENT), .A2(G_CURRENT), .ZN(n2) );
endmodule


module PG_PRIM_63 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_62 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_61 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_60 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_59 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_58 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_57 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_56 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_55 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(G) );
endmodule


module PG_PRIM_54 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_53 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_52 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_51 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_50 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_49 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_48 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_47 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_46 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_45 ( A, B, G, P );
  input A, B;
  output G, P;
  wire   n1, n2, n3, n4, n5;

  BUF_X1 U1 ( .A(B), .Z(n1) );
  NAND2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n2), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n4), .A2(n5), .ZN(P) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
  INV_X1 U6 ( .A(A), .ZN(n3) );
  AND2_X1 U7 ( .A1(A), .A2(n1), .ZN(G) );
endmodule


module PG_PRIM_44 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_43 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_42 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_41 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_40 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_39 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_38 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_37 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_36 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_35 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_34 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_PRIM_33 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module GG_73 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   net24509, n1, n2;
  assign G = net24509;

  NOR2_X1 U1 ( .A1(P_CURRENT), .A2(G_CURRENT), .ZN(n1) );
  NOR2_X1 U2 ( .A1(n2), .A2(n1), .ZN(net24509) );
  NOR2_X1 U3 ( .A1(G_PREV), .A2(G_CURRENT), .ZN(n2) );
endmodule


module GG_72 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_27 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_71 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_53 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_70 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_52 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_69 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_51 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_68 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_50 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_67 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_49 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_66 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_48 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_65 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_47 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_64 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_46 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_63 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_45 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_62 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_44 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_61 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_43 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_60 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_42 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_59 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_41 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_58 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_40 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_57 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   net24493, n1;
  assign G = net24493;

  AOI21_X1 U1 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net24493) );
endmodule


module GG_56 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_39 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_55 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_38 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_54 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_37 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_53 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_36 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_52 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_35 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_51 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_34 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_50 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_33 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_49 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   net24485, n1;
  assign G = net24485;

  AOI21_X1 U1 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net24485) );
endmodule


module GG_48 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_32 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_47 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_31 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_46 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_30 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_45 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GG_44 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   net24480, n1;
  assign G = net24480;

  AOI21_X1 U1 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net24480) );
endmodule


module GG_43 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_29 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_42 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module GP_28 ( P_CURRENT, P_PREV, P );
  input P_CURRENT, P_PREV;
  output P;


  AND2_X1 U1 ( .A1(P_PREV), .A2(P_CURRENT), .ZN(P) );
endmodule


module GG_41 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   net24477, n1;
  assign G = net24477;

  AOI21_X1 U1 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(net24477) );
endmodule


module GG_40 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n3) );
endmodule


module GG_39 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(G_PREV), .B2(P_CURRENT), .A(G_CURRENT), .ZN(n3) );
endmodule


module GG_38 ( G_CURRENT, P_CURRENT, G_PREV, G );
  input G_CURRENT, P_CURRENT, G_PREV;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(P_CURRENT), .B2(G_PREV), .A(G_CURRENT), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 ( A, B, CIN, CO );
  input [31:0] A;
  input [31:0] B;
  output [7:0] CO;
  input CIN;
  wire   n7, n8, n9, p_0, g_0, \cg_xbars[4][31][1] , \cg_xbars[4][31][0] ,
         \cg_xbars[4][27][1] , \cg_xbars[4][27][0] , \cg_xbars[3][31][1] ,
         \cg_xbars[3][31][0] , \cg_xbars[3][23][1] , \cg_xbars[3][23][0] ,
         \cg_xbars[3][15][1] , \cg_xbars[3][15][0] , \cg_xbars[2][31][1] ,
         \cg_xbars[2][31][0] , \cg_xbars[2][27][1] , \cg_xbars[2][27][0] ,
         \cg_xbars[2][23][1] , \cg_xbars[2][23][0] , \cg_xbars[2][19][1] ,
         \cg_xbars[2][19][0] , \cg_xbars[2][15][1] , \cg_xbars[2][15][0] ,
         \cg_xbars[2][11][1] , \cg_xbars[2][11][0] , \cg_xbars[2][7][1] ,
         \cg_xbars[2][7][0] , \cg_xbars[1][31][1] , \cg_xbars[1][31][0] ,
         \cg_xbars[1][29][1] , \cg_xbars[1][29][0] , \cg_xbars[1][27][1] ,
         \cg_xbars[1][27][0] , \cg_xbars[1][25][1] , \cg_xbars[1][25][0] ,
         \cg_xbars[1][23][1] , \cg_xbars[1][23][0] , \cg_xbars[1][21][1] ,
         \cg_xbars[1][21][0] , \cg_xbars[1][19][1] , \cg_xbars[1][19][0] ,
         \cg_xbars[1][17][1] , \cg_xbars[1][17][0] , \cg_xbars[1][15][1] ,
         \cg_xbars[1][15][0] , \cg_xbars[1][13][1] , \cg_xbars[1][13][0] ,
         \cg_xbars[1][11][1] , \cg_xbars[1][11][0] , \cg_xbars[1][9][1] ,
         \cg_xbars[1][9][0] , \cg_xbars[1][7][1] , \cg_xbars[1][7][0] ,
         \cg_xbars[1][5][1] , \cg_xbars[1][5][0] , \cg_xbars[1][3][1] ,
         \cg_xbars[1][3][0] , \cg_xbars[1][1][0] , \cg_xbars[0][31][1] ,
         \cg_xbars[0][31][0] , \cg_xbars[0][30][1] , \cg_xbars[0][30][0] ,
         \cg_xbars[0][29][1] , \cg_xbars[0][29][0] , \cg_xbars[0][28][1] ,
         \cg_xbars[0][28][0] , \cg_xbars[0][27][1] , \cg_xbars[0][27][0] ,
         \cg_xbars[0][26][1] , \cg_xbars[0][26][0] , \cg_xbars[0][25][1] ,
         \cg_xbars[0][25][0] , \cg_xbars[0][24][1] , \cg_xbars[0][24][0] ,
         \cg_xbars[0][23][1] , \cg_xbars[0][23][0] , \cg_xbars[0][22][1] ,
         \cg_xbars[0][22][0] , \cg_xbars[0][21][1] , \cg_xbars[0][21][0] ,
         \cg_xbars[0][20][1] , \cg_xbars[0][20][0] , \cg_xbars[0][19][1] ,
         \cg_xbars[0][19][0] , \cg_xbars[0][18][1] , \cg_xbars[0][18][0] ,
         \cg_xbars[0][17][1] , \cg_xbars[0][17][0] , \cg_xbars[0][16][1] ,
         \cg_xbars[0][16][0] , \cg_xbars[0][15][1] , \cg_xbars[0][15][0] ,
         \cg_xbars[0][14][1] , \cg_xbars[0][14][0] , \cg_xbars[0][13][1] ,
         \cg_xbars[0][13][0] , \cg_xbars[0][12][1] , \cg_xbars[0][12][0] ,
         \cg_xbars[0][11][1] , \cg_xbars[0][11][0] , \cg_xbars[0][10][1] ,
         \cg_xbars[0][10][0] , \cg_xbars[0][9][1] , \cg_xbars[0][9][0] ,
         \cg_xbars[0][8][1] , \cg_xbars[0][8][0] , \cg_xbars[0][7][1] ,
         \cg_xbars[0][7][0] , \cg_xbars[0][6][1] , \cg_xbars[0][6][0] ,
         \cg_xbars[0][5][1] , \cg_xbars[0][5][0] , \cg_xbars[0][4][1] ,
         \cg_xbars[0][4][0] , \cg_xbars[0][3][1] , \cg_xbars[0][3][0] ,
         \cg_xbars[0][2][1] , \cg_xbars[0][2][0] , \cg_xbars[0][1][1] ,
         \cg_xbars[0][1][0] , \cg_xbars[0][0][0] , n2, n5, n6;

  PG_PRIM_32 U_PG_PRIM_0 ( .A(A[0]), .B(B[0]), .G(g_0), .P(p_0) );
  GG_37 U_RXMOST_PG_PRIM_IS_GG_UNIT_0 ( .G_CURRENT(g_0), .P_CURRENT(p_0), 
        .G_PREV(CIN), .G(\cg_xbars[0][0][0] ) );
  PG_PRIM_63 U_PG_PRIM_1 ( .A(A[1]), .B(B[1]), .G(\cg_xbars[0][1][0] ), .P(
        \cg_xbars[0][1][1] ) );
  PG_PRIM_62 U_PG_PRIM_2 ( .A(A[2]), .B(B[2]), .G(\cg_xbars[0][2][0] ), .P(
        \cg_xbars[0][2][1] ) );
  PG_PRIM_61 U_PG_PRIM_3 ( .A(A[3]), .B(B[3]), .G(\cg_xbars[0][3][0] ), .P(
        \cg_xbars[0][3][1] ) );
  PG_PRIM_60 U_PG_PRIM_4 ( .A(A[4]), .B(B[4]), .G(\cg_xbars[0][4][0] ), .P(
        \cg_xbars[0][4][1] ) );
  PG_PRIM_59 U_PG_PRIM_5 ( .A(A[5]), .B(B[5]), .G(\cg_xbars[0][5][0] ), .P(
        \cg_xbars[0][5][1] ) );
  PG_PRIM_58 U_PG_PRIM_6 ( .A(A[6]), .B(B[6]), .G(\cg_xbars[0][6][0] ), .P(
        \cg_xbars[0][6][1] ) );
  PG_PRIM_57 U_PG_PRIM_7 ( .A(A[7]), .B(B[7]), .G(\cg_xbars[0][7][0] ), .P(
        \cg_xbars[0][7][1] ) );
  PG_PRIM_56 U_PG_PRIM_8 ( .A(A[8]), .B(B[8]), .G(\cg_xbars[0][8][0] ), .P(
        \cg_xbars[0][8][1] ) );
  PG_PRIM_55 U_PG_PRIM_9 ( .A(A[9]), .B(B[9]), .G(\cg_xbars[0][9][0] ), .P(
        \cg_xbars[0][9][1] ) );
  PG_PRIM_54 U_PG_PRIM_10 ( .A(A[10]), .B(B[10]), .G(\cg_xbars[0][10][0] ), 
        .P(\cg_xbars[0][10][1] ) );
  PG_PRIM_53 U_PG_PRIM_11 ( .A(A[11]), .B(B[11]), .G(\cg_xbars[0][11][0] ), 
        .P(\cg_xbars[0][11][1] ) );
  PG_PRIM_52 U_PG_PRIM_12 ( .A(A[12]), .B(B[12]), .G(\cg_xbars[0][12][0] ), 
        .P(\cg_xbars[0][12][1] ) );
  PG_PRIM_51 U_PG_PRIM_13 ( .A(A[13]), .B(B[13]), .G(\cg_xbars[0][13][0] ), 
        .P(\cg_xbars[0][13][1] ) );
  PG_PRIM_50 U_PG_PRIM_14 ( .A(A[14]), .B(B[14]), .G(\cg_xbars[0][14][0] ), 
        .P(\cg_xbars[0][14][1] ) );
  PG_PRIM_49 U_PG_PRIM_15 ( .A(A[15]), .B(B[15]), .G(\cg_xbars[0][15][0] ), 
        .P(\cg_xbars[0][15][1] ) );
  PG_PRIM_48 U_PG_PRIM_16 ( .A(A[16]), .B(B[16]), .G(\cg_xbars[0][16][0] ), 
        .P(\cg_xbars[0][16][1] ) );
  PG_PRIM_47 U_PG_PRIM_17 ( .A(A[17]), .B(B[17]), .G(\cg_xbars[0][17][0] ), 
        .P(\cg_xbars[0][17][1] ) );
  PG_PRIM_46 U_PG_PRIM_18 ( .A(A[18]), .B(B[18]), .G(\cg_xbars[0][18][0] ), 
        .P(\cg_xbars[0][18][1] ) );
  PG_PRIM_45 U_PG_PRIM_19 ( .A(A[19]), .B(B[19]), .G(\cg_xbars[0][19][0] ), 
        .P(\cg_xbars[0][19][1] ) );
  PG_PRIM_44 U_PG_PRIM_20 ( .A(A[20]), .B(B[20]), .G(\cg_xbars[0][20][0] ), 
        .P(\cg_xbars[0][20][1] ) );
  PG_PRIM_43 U_PG_PRIM_21 ( .A(A[21]), .B(B[21]), .G(\cg_xbars[0][21][0] ), 
        .P(\cg_xbars[0][21][1] ) );
  PG_PRIM_42 U_PG_PRIM_22 ( .A(A[22]), .B(B[22]), .G(\cg_xbars[0][22][0] ), 
        .P(\cg_xbars[0][22][1] ) );
  PG_PRIM_41 U_PG_PRIM_23 ( .A(A[23]), .B(B[23]), .G(\cg_xbars[0][23][0] ), 
        .P(\cg_xbars[0][23][1] ) );
  PG_PRIM_40 U_PG_PRIM_24 ( .A(A[24]), .B(B[24]), .G(\cg_xbars[0][24][0] ), 
        .P(\cg_xbars[0][24][1] ) );
  PG_PRIM_39 U_PG_PRIM_25 ( .A(A[25]), .B(B[25]), .G(\cg_xbars[0][25][0] ), 
        .P(\cg_xbars[0][25][1] ) );
  PG_PRIM_38 U_PG_PRIM_26 ( .A(A[26]), .B(B[26]), .G(\cg_xbars[0][26][0] ), 
        .P(\cg_xbars[0][26][1] ) );
  PG_PRIM_37 U_PG_PRIM_27 ( .A(A[27]), .B(B[27]), .G(\cg_xbars[0][27][0] ), 
        .P(\cg_xbars[0][27][1] ) );
  PG_PRIM_36 U_PG_PRIM_28 ( .A(A[28]), .B(B[28]), .G(\cg_xbars[0][28][0] ), 
        .P(\cg_xbars[0][28][1] ) );
  PG_PRIM_35 U_PG_PRIM_29 ( .A(A[29]), .B(B[29]), .G(\cg_xbars[0][29][0] ), 
        .P(\cg_xbars[0][29][1] ) );
  PG_PRIM_34 U_PG_PRIM_30 ( .A(A[30]), .B(B[30]), .G(\cg_xbars[0][30][0] ), 
        .P(\cg_xbars[0][30][1] ) );
  PG_PRIM_33 U_PG_PRIM_31 ( .A(A[31]), .B(B[31]), .G(\cg_xbars[0][31][0] ), 
        .P(\cg_xbars[0][31][1] ) );
  GG_73 U_BKBONE_GG_UNIT_1_1 ( .G_CURRENT(\cg_xbars[0][1][0] ), .P_CURRENT(
        \cg_xbars[0][1][1] ), .G_PREV(\cg_xbars[0][0][0] ), .G(
        \cg_xbars[1][1][0] ) );
  GG_72 U_BKBONE_GG_UNIT_1_3 ( .G_CURRENT(\cg_xbars[0][3][0] ), .P_CURRENT(
        \cg_xbars[0][3][1] ), .G_PREV(\cg_xbars[0][2][0] ), .G(
        \cg_xbars[1][3][0] ) );
  GP_27 U_BKBONE_GP_UNIT_1_3 ( .P_CURRENT(\cg_xbars[0][3][1] ), .P_PREV(
        \cg_xbars[0][2][1] ), .P(\cg_xbars[1][3][1] ) );
  GG_71 U_BKBONE_GG_UNIT_1_5 ( .G_CURRENT(\cg_xbars[0][5][0] ), .P_CURRENT(
        \cg_xbars[0][5][1] ), .G_PREV(\cg_xbars[0][4][0] ), .G(
        \cg_xbars[1][5][0] ) );
  GP_53 U_BKBONE_GP_UNIT_1_5 ( .P_CURRENT(\cg_xbars[0][5][1] ), .P_PREV(
        \cg_xbars[0][4][1] ), .P(\cg_xbars[1][5][1] ) );
  GG_70 U_BKBONE_GG_UNIT_1_7 ( .G_CURRENT(\cg_xbars[0][7][0] ), .P_CURRENT(
        \cg_xbars[0][7][1] ), .G_PREV(\cg_xbars[0][6][0] ), .G(
        \cg_xbars[1][7][0] ) );
  GP_52 U_BKBONE_GP_UNIT_1_7 ( .P_CURRENT(\cg_xbars[0][7][1] ), .P_PREV(
        \cg_xbars[0][6][1] ), .P(\cg_xbars[1][7][1] ) );
  GG_69 U_BKBONE_GG_UNIT_1_9 ( .G_CURRENT(\cg_xbars[0][9][0] ), .P_CURRENT(
        \cg_xbars[0][9][1] ), .G_PREV(\cg_xbars[0][8][0] ), .G(
        \cg_xbars[1][9][0] ) );
  GP_51 U_BKBONE_GP_UNIT_1_9 ( .P_CURRENT(\cg_xbars[0][9][1] ), .P_PREV(
        \cg_xbars[0][8][1] ), .P(\cg_xbars[1][9][1] ) );
  GG_68 U_BKBONE_GG_UNIT_1_11 ( .G_CURRENT(\cg_xbars[0][11][0] ), .P_CURRENT(
        \cg_xbars[0][11][1] ), .G_PREV(\cg_xbars[0][10][0] ), .G(
        \cg_xbars[1][11][0] ) );
  GP_50 U_BKBONE_GP_UNIT_1_11 ( .P_CURRENT(\cg_xbars[0][11][1] ), .P_PREV(
        \cg_xbars[0][10][1] ), .P(\cg_xbars[1][11][1] ) );
  GG_67 U_BKBONE_GG_UNIT_1_13 ( .G_CURRENT(\cg_xbars[0][13][0] ), .P_CURRENT(
        \cg_xbars[0][13][1] ), .G_PREV(\cg_xbars[0][12][0] ), .G(
        \cg_xbars[1][13][0] ) );
  GP_49 U_BKBONE_GP_UNIT_1_13 ( .P_CURRENT(\cg_xbars[0][13][1] ), .P_PREV(
        \cg_xbars[0][12][1] ), .P(\cg_xbars[1][13][1] ) );
  GG_66 U_BKBONE_GG_UNIT_1_15 ( .G_CURRENT(\cg_xbars[0][15][0] ), .P_CURRENT(
        \cg_xbars[0][15][1] ), .G_PREV(\cg_xbars[0][14][0] ), .G(
        \cg_xbars[1][15][0] ) );
  GP_48 U_BKBONE_GP_UNIT_1_15 ( .P_CURRENT(\cg_xbars[0][15][1] ), .P_PREV(
        \cg_xbars[0][14][1] ), .P(\cg_xbars[1][15][1] ) );
  GG_65 U_BKBONE_GG_UNIT_1_17 ( .G_CURRENT(\cg_xbars[0][17][0] ), .P_CURRENT(
        \cg_xbars[0][17][1] ), .G_PREV(\cg_xbars[0][16][0] ), .G(
        \cg_xbars[1][17][0] ) );
  GP_47 U_BKBONE_GP_UNIT_1_17 ( .P_CURRENT(\cg_xbars[0][17][1] ), .P_PREV(
        \cg_xbars[0][16][1] ), .P(\cg_xbars[1][17][1] ) );
  GG_64 U_BKBONE_GG_UNIT_1_19 ( .G_CURRENT(\cg_xbars[0][19][0] ), .P_CURRENT(
        \cg_xbars[0][19][1] ), .G_PREV(\cg_xbars[0][18][0] ), .G(
        \cg_xbars[1][19][0] ) );
  GP_46 U_BKBONE_GP_UNIT_1_19 ( .P_CURRENT(\cg_xbars[0][19][1] ), .P_PREV(
        \cg_xbars[0][18][1] ), .P(\cg_xbars[1][19][1] ) );
  GG_63 U_BKBONE_GG_UNIT_1_21 ( .G_CURRENT(\cg_xbars[0][21][0] ), .P_CURRENT(
        \cg_xbars[0][21][1] ), .G_PREV(\cg_xbars[0][20][0] ), .G(
        \cg_xbars[1][21][0] ) );
  GP_45 U_BKBONE_GP_UNIT_1_21 ( .P_CURRENT(\cg_xbars[0][21][1] ), .P_PREV(
        \cg_xbars[0][20][1] ), .P(\cg_xbars[1][21][1] ) );
  GG_62 U_BKBONE_GG_UNIT_1_23 ( .G_CURRENT(\cg_xbars[0][23][0] ), .P_CURRENT(
        \cg_xbars[0][23][1] ), .G_PREV(\cg_xbars[0][22][0] ), .G(
        \cg_xbars[1][23][0] ) );
  GP_44 U_BKBONE_GP_UNIT_1_23 ( .P_CURRENT(\cg_xbars[0][23][1] ), .P_PREV(
        \cg_xbars[0][22][1] ), .P(\cg_xbars[1][23][1] ) );
  GG_61 U_BKBONE_GG_UNIT_1_25 ( .G_CURRENT(\cg_xbars[0][25][0] ), .P_CURRENT(
        \cg_xbars[0][25][1] ), .G_PREV(\cg_xbars[0][24][0] ), .G(
        \cg_xbars[1][25][0] ) );
  GP_43 U_BKBONE_GP_UNIT_1_25 ( .P_CURRENT(\cg_xbars[0][25][1] ), .P_PREV(
        \cg_xbars[0][24][1] ), .P(\cg_xbars[1][25][1] ) );
  GG_60 U_BKBONE_GG_UNIT_1_27 ( .G_CURRENT(\cg_xbars[0][27][0] ), .P_CURRENT(
        \cg_xbars[0][27][1] ), .G_PREV(\cg_xbars[0][26][0] ), .G(
        \cg_xbars[1][27][0] ) );
  GP_42 U_BKBONE_GP_UNIT_1_27 ( .P_CURRENT(\cg_xbars[0][27][1] ), .P_PREV(
        \cg_xbars[0][26][1] ), .P(\cg_xbars[1][27][1] ) );
  GG_59 U_BKBONE_GG_UNIT_1_29 ( .G_CURRENT(\cg_xbars[0][29][0] ), .P_CURRENT(
        \cg_xbars[0][29][1] ), .G_PREV(\cg_xbars[0][28][0] ), .G(
        \cg_xbars[1][29][0] ) );
  GP_41 U_BKBONE_GP_UNIT_1_29 ( .P_CURRENT(\cg_xbars[0][29][1] ), .P_PREV(
        \cg_xbars[0][28][1] ), .P(\cg_xbars[1][29][1] ) );
  GG_58 U_BKBONE_GG_UNIT_1_31 ( .G_CURRENT(\cg_xbars[0][31][0] ), .P_CURRENT(
        \cg_xbars[0][31][1] ), .G_PREV(\cg_xbars[0][30][0] ), .G(
        \cg_xbars[1][31][0] ) );
  GP_40 U_BKBONE_GP_UNIT_1_31 ( .P_CURRENT(\cg_xbars[0][31][1] ), .P_PREV(
        \cg_xbars[0][30][1] ), .P(\cg_xbars[1][31][1] ) );
  GG_57 U_BKBONE_GG_UNIT_2_3 ( .G_CURRENT(\cg_xbars[1][3][0] ), .P_CURRENT(
        \cg_xbars[1][3][1] ), .G_PREV(\cg_xbars[1][1][0] ), .G(n9) );
  GG_56 U_BKBONE_GG_UNIT_2_7 ( .G_CURRENT(\cg_xbars[1][7][0] ), .P_CURRENT(
        \cg_xbars[1][7][1] ), .G_PREV(\cg_xbars[1][5][0] ), .G(
        \cg_xbars[2][7][0] ) );
  GP_39 U_BKBONE_GP_UNIT_2_7 ( .P_CURRENT(\cg_xbars[1][7][1] ), .P_PREV(
        \cg_xbars[1][5][1] ), .P(\cg_xbars[2][7][1] ) );
  GG_55 U_BKBONE_GG_UNIT_2_11 ( .G_CURRENT(\cg_xbars[1][11][0] ), .P_CURRENT(
        \cg_xbars[1][11][1] ), .G_PREV(\cg_xbars[1][9][0] ), .G(
        \cg_xbars[2][11][0] ) );
  GP_38 U_BKBONE_GP_UNIT_2_11 ( .P_CURRENT(\cg_xbars[1][11][1] ), .P_PREV(
        \cg_xbars[1][9][1] ), .P(\cg_xbars[2][11][1] ) );
  GG_54 U_BKBONE_GG_UNIT_2_15 ( .G_CURRENT(\cg_xbars[1][15][0] ), .P_CURRENT(
        \cg_xbars[1][15][1] ), .G_PREV(\cg_xbars[1][13][0] ), .G(
        \cg_xbars[2][15][0] ) );
  GP_37 U_BKBONE_GP_UNIT_2_15 ( .P_CURRENT(\cg_xbars[1][15][1] ), .P_PREV(
        \cg_xbars[1][13][1] ), .P(\cg_xbars[2][15][1] ) );
  GG_53 U_BKBONE_GG_UNIT_2_19 ( .G_CURRENT(\cg_xbars[1][19][0] ), .P_CURRENT(
        \cg_xbars[1][19][1] ), .G_PREV(\cg_xbars[1][17][0] ), .G(
        \cg_xbars[2][19][0] ) );
  GP_36 U_BKBONE_GP_UNIT_2_19 ( .P_CURRENT(\cg_xbars[1][19][1] ), .P_PREV(
        \cg_xbars[1][17][1] ), .P(\cg_xbars[2][19][1] ) );
  GG_52 U_BKBONE_GG_UNIT_2_23 ( .G_CURRENT(\cg_xbars[1][23][0] ), .P_CURRENT(
        \cg_xbars[1][23][1] ), .G_PREV(\cg_xbars[1][21][0] ), .G(
        \cg_xbars[2][23][0] ) );
  GP_35 U_BKBONE_GP_UNIT_2_23 ( .P_CURRENT(\cg_xbars[1][23][1] ), .P_PREV(
        \cg_xbars[1][21][1] ), .P(\cg_xbars[2][23][1] ) );
  GG_51 U_BKBONE_GG_UNIT_2_27 ( .G_CURRENT(\cg_xbars[1][27][0] ), .P_CURRENT(
        \cg_xbars[1][27][1] ), .G_PREV(\cg_xbars[1][25][0] ), .G(
        \cg_xbars[2][27][0] ) );
  GP_34 U_BKBONE_GP_UNIT_2_27 ( .P_CURRENT(\cg_xbars[1][27][1] ), .P_PREV(
        \cg_xbars[1][25][1] ), .P(\cg_xbars[2][27][1] ) );
  GG_50 U_BKBONE_GG_UNIT_2_31 ( .G_CURRENT(\cg_xbars[1][31][0] ), .P_CURRENT(
        \cg_xbars[1][31][1] ), .G_PREV(\cg_xbars[1][29][0] ), .G(
        \cg_xbars[2][31][0] ) );
  GP_33 U_BKBONE_GP_UNIT_2_31 ( .P_CURRENT(\cg_xbars[1][31][1] ), .P_PREV(
        \cg_xbars[1][29][1] ), .P(\cg_xbars[2][31][1] ) );
  GG_49 U_LF_GG_UNIT_1_7 ( .G_CURRENT(\cg_xbars[2][7][0] ), .P_CURRENT(
        \cg_xbars[2][7][1] ), .G_PREV(n9), .G(n8) );
  GG_48 U_LF_GG_UNIT_1_15 ( .G_CURRENT(\cg_xbars[2][15][0] ), .P_CURRENT(
        \cg_xbars[2][15][1] ), .G_PREV(\cg_xbars[2][11][0] ), .G(
        \cg_xbars[3][15][0] ) );
  GP_32 U_LF_GP_UNIT_1_15 ( .P_CURRENT(\cg_xbars[2][15][1] ), .P_PREV(
        \cg_xbars[2][11][1] ), .P(\cg_xbars[3][15][1] ) );
  GG_47 U_LF_GG_UNIT_1_23 ( .G_CURRENT(\cg_xbars[2][23][0] ), .P_CURRENT(
        \cg_xbars[2][23][1] ), .G_PREV(\cg_xbars[2][19][0] ), .G(
        \cg_xbars[3][23][0] ) );
  GP_31 U_LF_GP_UNIT_1_23 ( .P_CURRENT(\cg_xbars[2][23][1] ), .P_PREV(
        \cg_xbars[2][19][1] ), .P(\cg_xbars[3][23][1] ) );
  GG_46 U_LF_GG_UNIT_1_31 ( .G_CURRENT(\cg_xbars[2][31][0] ), .P_CURRENT(
        \cg_xbars[2][31][1] ), .G_PREV(\cg_xbars[2][27][0] ), .G(
        \cg_xbars[3][31][0] ) );
  GP_30 U_LF_GP_UNIT_1_31 ( .P_CURRENT(\cg_xbars[2][31][1] ), .P_PREV(
        \cg_xbars[2][27][1] ), .P(\cg_xbars[3][31][1] ) );
  GG_45 U_LF_GG_UNIT_2_11 ( .G_CURRENT(n5), .P_CURRENT(\cg_xbars[2][11][1] ), 
        .G_PREV(n6), .G(CO[2]) );
  GG_44 U_LF_GG_UNIT_2_15 ( .G_CURRENT(\cg_xbars[3][15][0] ), .P_CURRENT(
        \cg_xbars[3][15][1] ), .G_PREV(n8), .G(n7) );
  GG_43 U_LF_GG_UNIT_2_27 ( .G_CURRENT(\cg_xbars[2][27][0] ), .P_CURRENT(
        \cg_xbars[2][27][1] ), .G_PREV(\cg_xbars[3][23][0] ), .G(
        \cg_xbars[4][27][0] ) );
  GP_29 U_LF_GP_UNIT_2_27 ( .P_CURRENT(\cg_xbars[2][27][1] ), .P_PREV(
        \cg_xbars[3][23][1] ), .P(\cg_xbars[4][27][1] ) );
  GG_42 U_LF_GG_UNIT_2_31 ( .G_CURRENT(\cg_xbars[3][31][0] ), .P_CURRENT(
        \cg_xbars[3][31][1] ), .G_PREV(n2), .G(\cg_xbars[4][31][0] ) );
  GP_28 U_LF_GP_UNIT_2_31 ( .P_CURRENT(\cg_xbars[3][31][1] ), .P_PREV(
        \cg_xbars[3][23][1] ), .P(\cg_xbars[4][31][1] ) );
  GG_41 U_LF_GG_UNIT_3_19 ( .G_CURRENT(\cg_xbars[2][19][0] ), .P_CURRENT(
        \cg_xbars[2][19][1] ), .G_PREV(n7), .G(CO[4]) );
  GG_40 U_LF_GG_UNIT_3_23 ( .G_CURRENT(n2), .P_CURRENT(\cg_xbars[3][23][1] ), 
        .G_PREV(n7), .G(CO[5]) );
  GG_39 U_LF_GG_UNIT_3_27 ( .G_CURRENT(\cg_xbars[4][27][0] ), .P_CURRENT(
        \cg_xbars[4][27][1] ), .G_PREV(n7), .G(CO[6]) );
  GG_38 U_LF_GG_UNIT_3_31 ( .G_CURRENT(\cg_xbars[4][31][0] ), .P_CURRENT(
        \cg_xbars[4][31][1] ), .G_PREV(CO[3]), .G(CO[7]) );
  CLKBUF_X1 U1 ( .A(n8), .Z(n6) );
  BUF_X1 U2 ( .A(n6), .Z(CO[1]) );
  BUF_X1 U3 ( .A(n7), .Z(CO[3]) );
  CLKBUF_X1 U4 ( .A(\cg_xbars[3][23][0] ), .Z(n2) );
  CLKBUF_X1 U5 ( .A(n9), .Z(CO[0]) );
  CLKBUF_X1 U6 ( .A(\cg_xbars[2][11][0] ), .Z(n5) );
endmodule


module RCA_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_7 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n7, n8, n9, n10, n11, n6;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_NBIT4_29 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_28 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  INV_X1 U3 ( .A(Cin), .ZN(n6) );
  INV_X1 U4 ( .A(n11), .ZN(Co) );
  INV_X1 U5 ( .A(n7), .ZN(S[3]) );
  AOI22_X1 U6 ( .A1(S0[3]), .A2(n6), .B1(S1[3]), .B2(Cin), .ZN(n7) );
  INV_X1 U7 ( .A(n9), .ZN(S[1]) );
  AOI22_X1 U8 ( .A1(S0[1]), .A2(n6), .B1(S1[1]), .B2(Cin), .ZN(n9) );
  INV_X1 U9 ( .A(n8), .ZN(S[2]) );
  AOI22_X1 U10 ( .A1(S0[2]), .A2(n6), .B1(S1[2]), .B2(Cin), .ZN(n8) );
  AOI22_X1 U11 ( .A1(Co0), .A2(n6), .B1(Co1), .B2(Cin), .ZN(n11) );
  INV_X1 U12 ( .A(n10), .ZN(S[0]) );
  AOI22_X1 U13 ( .A1(S0[0]), .A2(n6), .B1(S1[0]), .B2(Cin), .ZN(n10) );
endmodule


module RCA_NBIT4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_13 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n6, n12, n13, n14, n15, n16;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_NBIT4_27 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_26 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  INV_X1 U3 ( .A(Cin), .ZN(n6) );
  INV_X1 U4 ( .A(n12), .ZN(Co) );
  INV_X1 U5 ( .A(n14), .ZN(S[1]) );
  AOI22_X1 U6 ( .A1(S0[1]), .A2(n6), .B1(S1[1]), .B2(Cin), .ZN(n14) );
  INV_X1 U7 ( .A(n15), .ZN(S[2]) );
  AOI22_X1 U8 ( .A1(S0[2]), .A2(n6), .B1(S1[2]), .B2(Cin), .ZN(n15) );
  INV_X1 U9 ( .A(n16), .ZN(S[3]) );
  AOI22_X1 U10 ( .A1(S0[3]), .A2(n6), .B1(S1[3]), .B2(Cin), .ZN(n16) );
  AOI22_X1 U11 ( .A1(Co0), .A2(n6), .B1(Co1), .B2(Cin), .ZN(n12) );
  INV_X1 U12 ( .A(n13), .ZN(S[0]) );
  AOI22_X1 U13 ( .A1(S0[0]), .A2(n6), .B1(S1[0]), .B2(Cin), .ZN(n13) );
endmodule


module RCA_NBIT4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_12 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n1, n2, n3, n4, n15, n16, n17, n18, n19, n20;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_NBIT4_25 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_24 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  CLKBUF_X1 U3 ( .A(Cin), .Z(n1) );
  CLKBUF_X1 U4 ( .A(Cin), .Z(n2) );
  INV_X1 U5 ( .A(n4), .ZN(n3) );
  INV_X1 U6 ( .A(n1), .ZN(n4) );
  INV_X1 U7 ( .A(Cin), .ZN(n15) );
  INV_X1 U8 ( .A(n16), .ZN(Co) );
  INV_X1 U9 ( .A(n18), .ZN(S[1]) );
  AOI22_X1 U10 ( .A1(S0[1]), .A2(n15), .B1(S1[1]), .B2(Cin), .ZN(n18) );
  INV_X1 U11 ( .A(n19), .ZN(S[2]) );
  AOI22_X1 U12 ( .A1(S0[2]), .A2(n15), .B1(S1[2]), .B2(Cin), .ZN(n19) );
  INV_X1 U13 ( .A(n20), .ZN(S[3]) );
  AOI22_X1 U14 ( .A1(S0[3]), .A2(n4), .B1(S1[3]), .B2(n2), .ZN(n20) );
  AOI22_X1 U15 ( .A1(Co0), .A2(n4), .B1(Co1), .B2(n3), .ZN(n16) );
  INV_X1 U16 ( .A(n17), .ZN(S[0]) );
  AOI22_X1 U17 ( .A1(n15), .A2(S0[0]), .B1(S1[0]), .B2(Cin), .ZN(n17) );
endmodule


module RCA_NBIT4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_11 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n6, n12, n13, n14, n15, n16;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_NBIT4_23 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_22 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  INV_X1 U3 ( .A(n12), .ZN(Co) );
  INV_X1 U4 ( .A(n14), .ZN(S[1]) );
  INV_X1 U5 ( .A(n15), .ZN(S[2]) );
  INV_X1 U6 ( .A(n16), .ZN(S[3]) );
  INV_X1 U7 ( .A(n13), .ZN(S[0]) );
  AOI22_X1 U8 ( .A1(Co0), .A2(n6), .B1(Co1), .B2(Cin), .ZN(n12) );
  AOI22_X1 U9 ( .A1(S0[3]), .A2(n6), .B1(S1[3]), .B2(Cin), .ZN(n16) );
  AOI22_X1 U10 ( .A1(S0[2]), .A2(n6), .B1(S1[2]), .B2(Cin), .ZN(n15) );
  AOI22_X1 U11 ( .A1(S0[1]), .A2(n6), .B1(S1[1]), .B2(Cin), .ZN(n14) );
  AOI22_X1 U12 ( .A1(S0[0]), .A2(n6), .B1(S1[0]), .B2(Cin), .ZN(n13) );
  INV_X1 U13 ( .A(Cin), .ZN(n6) );
endmodule


module RCA_NBIT4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_10 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n9, n11, net24522, net24523, net24524, net24527, net34862,
         n1, n2, n3, n4, n5, n12, n13;
  wire   [3:0] S0;
  wire   [3:0] S1;
  assign S[0] = net24523;
  assign S[1] = net24524;
  assign Co = net24527;

  RCA_NBIT4_21 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_20 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  CLKBUF_X1 U3 ( .A(Cin), .Z(n1) );
  AOI22_X1 U4 ( .A1(S0[0]), .A2(n3), .B1(n5), .B2(S1[0]), .ZN(n2) );
  INV_X1 U5 ( .A(n2), .ZN(net24523) );
  CLKBUF_X1 U6 ( .A(Cin), .Z(n5) );
  INV_X1 U7 ( .A(Cin), .ZN(n3) );
  AOI22_X1 U8 ( .A1(S0[1]), .A2(n3), .B1(net34862), .B2(S1[1]), .ZN(n9) );
  INV_X1 U9 ( .A(n3), .ZN(n4) );
  AOI22_X1 U10 ( .A1(Co0), .A2(n3), .B1(Co1), .B2(n4), .ZN(n11) );
  CLKBUF_X1 U11 ( .A(Cin), .Z(net34862) );
  INV_X1 U12 ( .A(Cin), .ZN(net24522) );
  INV_X1 U13 ( .A(n11), .ZN(net24527) );
  AOI22_X1 U14 ( .A1(S0[2]), .A2(net24522), .B1(Cin), .B2(S1[2]), .ZN(n12) );
  AOI22_X1 U15 ( .A1(S0[3]), .A2(net24522), .B1(n1), .B2(S1[3]), .ZN(n13) );
  INV_X1 U16 ( .A(n13), .ZN(S[3]) );
  INV_X1 U17 ( .A(n12), .ZN(S[2]) );
  INV_X1 U18 ( .A(n9), .ZN(net24524) );
endmodule


module RCA_NBIT4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_9 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n1, n2, n3, n4, n6, n10, n12, n17, n18, n19, n20, n21;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_NBIT4_19 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_18 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  CLKBUF_X1 U3 ( .A(Cin), .Z(n1) );
  CLKBUF_X1 U4 ( .A(Cin), .Z(n2) );
  CLKBUF_X1 U5 ( .A(Cin), .Z(n3) );
  CLKBUF_X1 U6 ( .A(Cin), .Z(n12) );
  INV_X1 U7 ( .A(n3), .ZN(n4) );
  INV_X1 U8 ( .A(S0[0]), .ZN(n6) );
  INV_X1 U9 ( .A(S1[0]), .ZN(n10) );
  OAI22_X1 U10 ( .A1(n6), .A2(n12), .B1(n10), .B2(n4), .ZN(S[0]) );
  INV_X1 U11 ( .A(Cin), .ZN(n17) );
  INV_X1 U12 ( .A(n18), .ZN(Co) );
  AOI22_X1 U13 ( .A1(S0[1]), .A2(n17), .B1(n2), .B2(S1[1]), .ZN(n19) );
  AOI22_X1 U14 ( .A1(n17), .A2(S0[2]), .B1(Cin), .B2(S1[2]), .ZN(n20) );
  AOI22_X1 U15 ( .A1(S0[3]), .A2(n17), .B1(n1), .B2(S1[3]), .ZN(n21) );
  AOI22_X1 U16 ( .A1(Co0), .A2(n4), .B1(Co1), .B2(n12), .ZN(n18) );
  INV_X1 U17 ( .A(n19), .ZN(S[1]) );
  INV_X1 U18 ( .A(n21), .ZN(S[3]) );
  INV_X1 U19 ( .A(n20), .ZN(S[2]) );
endmodule


module RCA_NBIT4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_74_2/carry[3] , \add_1_root_add_74_2/carry[2] ,
         \add_1_root_add_74_2/carry[1] ;

  FA_X1 \add_1_root_add_74_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_74_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_74_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_74_2/carry[1] ), .CO(\add_1_root_add_74_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_74_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_74_2/carry[2] ), .CO(\add_1_root_add_74_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_74_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_74_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module CSB_NBIT4_8 ( A, B, Cin, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output Co;
  wire   Co0, Co1, n1, n2, n4, n5, n14, n15, n16, n17, n18;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_NBIT4_17 U_RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(S0), .Co(Co0) );
  RCA_NBIT4_16 U_RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(S1), .Co(Co1) );
  CLKBUF_X1 U3 ( .A(Cin), .Z(n1) );
  INV_X1 U4 ( .A(S0[0]), .ZN(n4) );
  INV_X1 U5 ( .A(Cin), .ZN(n2) );
  INV_X1 U6 ( .A(S1[0]), .ZN(n5) );
  OAI22_X1 U7 ( .A1(n1), .A2(n4), .B1(n5), .B2(n2), .ZN(S[0]) );
  INV_X1 U8 ( .A(Cin), .ZN(n14) );
  INV_X1 U9 ( .A(n15), .ZN(Co) );
  AOI22_X1 U10 ( .A1(n14), .A2(S0[2]), .B1(Cin), .B2(S1[2]), .ZN(n17) );
  AOI22_X1 U11 ( .A1(n14), .A2(S0[1]), .B1(Cin), .B2(S1[1]), .ZN(n16) );
  AOI22_X1 U12 ( .A1(S0[3]), .A2(n2), .B1(Cin), .B2(S1[3]), .ZN(n18) );
  AOI22_X1 U13 ( .A1(Co0), .A2(n14), .B1(Co1), .B2(n1), .ZN(n15) );
  INV_X1 U14 ( .A(n18), .ZN(S[3]) );
  INV_X1 U15 ( .A(n16), .ZN(S[1]) );
  INV_X1 U16 ( .A(n17), .ZN(S[2]) );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS7_1 ( A, B, Ci, S );
  input [27:0] A;
  input [27:0] B;
  input [6:0] Ci;
  output [27:0] S;


  CSB_NBIT4_7 U_CSB_1 ( .A(A[3:0]), .B(B[3:0]), .Cin(Ci[0]), .S(S[3:0]) );
  CSB_NBIT4_13 U_CSB_2 ( .A(A[7:4]), .B(B[7:4]), .Cin(Ci[1]), .S(S[7:4]) );
  CSB_NBIT4_12 U_CSB_3 ( .A(A[11:8]), .B(B[11:8]), .Cin(Ci[2]), .S(S[11:8]) );
  CSB_NBIT4_11 U_CSB_4 ( .A(A[15:12]), .B(B[15:12]), .Cin(Ci[3]), .S(S[15:12])
         );
  CSB_NBIT4_10 U_CSB_5 ( .A(A[19:16]), .B(B[19:16]), .Cin(Ci[4]), .S(S[19:16])
         );
  CSB_NBIT4_9 U_CSB_6 ( .A(A[23:20]), .B(B[23:20]), .Cin(Ci[5]), .S(S[23:20])
         );
  CSB_NBIT4_8 U_CSB_7 ( .A(A[27:24]), .B(B[27:24]), .Cin(Ci[6]), .S(S[27:24])
         );
endmodule


module P4_ADDER_NBIT32_1 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [6:0] carry_gen_Co;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 U_CARRY_GENERATOR ( .A(A), .B(B), 
        .CIN(Cin), .CO({Cout, carry_gen_Co}) );
  RCA_NBIT4_15 U_FIRST_RCA ( .A(A[3:0]), .B({B[3:1], n6}), .Ci(Cin), .S(S[3:0]) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS7_1 U_SUM_GENERATOR ( .A(A[31:4]), .B({
        B[31:20], n2, B[18:16], n5, B[14], n1, B[12], n4, B[10], n3, B[8:4]}), 
        .Ci(carry_gen_Co), .S(S[31:4]) );
  CLKBUF_X1 U1 ( .A(B[13]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[19]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(B[9]), .Z(n3) );
  CLKBUF_X1 U4 ( .A(B[11]), .Z(n4) );
  CLKBUF_X1 U5 ( .A(B[15]), .Z(n5) );
  CLKBUF_X1 U6 ( .A(B[0]), .Z(n6) );
endmodule


module T2_LOGIC_DATA_W32_1 ( OP, A, B, S );
  input [3:0] OP;
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n129, n130, n131, n132, n133,
         n134, n135, n136, n137;

  BUF_X1 U1 ( .A(OP[3]), .Z(n2) );
  BUF_X1 U2 ( .A(OP[3]), .Z(n3) );
  BUF_X1 U3 ( .A(OP[3]), .Z(n1) );
  INV_X1 U4 ( .A(A[2]), .ZN(n39) );
  INV_X1 U5 ( .A(A[3]), .ZN(n38) );
  BUF_X1 U6 ( .A(OP[2]), .Z(n8) );
  BUF_X1 U7 ( .A(OP[2]), .Z(n7) );
  BUF_X1 U8 ( .A(OP[1]), .Z(n5) );
  BUF_X1 U9 ( .A(OP[1]), .Z(n6) );
  BUF_X1 U10 ( .A(OP[1]), .Z(n4) );
  BUF_X1 U11 ( .A(OP[2]), .Z(n9) );
  INV_X1 U12 ( .A(A[31]), .ZN(n10) );
  INV_X1 U13 ( .A(A[30]), .ZN(n11) );
  INV_X1 U14 ( .A(A[7]), .ZN(n34) );
  INV_X1 U15 ( .A(A[16]), .ZN(n25) );
  INV_X1 U16 ( .A(A[17]), .ZN(n24) );
  INV_X1 U17 ( .A(A[18]), .ZN(n23) );
  INV_X1 U18 ( .A(A[19]), .ZN(n22) );
  INV_X1 U19 ( .A(A[20]), .ZN(n21) );
  INV_X1 U20 ( .A(A[21]), .ZN(n20) );
  INV_X1 U21 ( .A(A[22]), .ZN(n19) );
  INV_X1 U22 ( .A(A[23]), .ZN(n18) );
  INV_X1 U23 ( .A(A[8]), .ZN(n33) );
  INV_X1 U24 ( .A(A[6]), .ZN(n35) );
  INV_X1 U25 ( .A(A[9]), .ZN(n32) );
  INV_X1 U26 ( .A(A[24]), .ZN(n17) );
  INV_X1 U27 ( .A(A[26]), .ZN(n15) );
  INV_X1 U28 ( .A(A[27]), .ZN(n14) );
  INV_X1 U29 ( .A(A[29]), .ZN(n12) );
  INV_X1 U30 ( .A(A[10]), .ZN(n31) );
  INV_X1 U31 ( .A(A[11]), .ZN(n30) );
  INV_X1 U32 ( .A(A[12]), .ZN(n29) );
  INV_X1 U33 ( .A(A[13]), .ZN(n28) );
  INV_X1 U34 ( .A(A[14]), .ZN(n27) );
  INV_X1 U35 ( .A(A[15]), .ZN(n26) );
  INV_X1 U36 ( .A(A[25]), .ZN(n16) );
  INV_X1 U37 ( .A(A[28]), .ZN(n13) );
  AOI22_X1 U38 ( .A1(OP[0]), .A2(n39), .B1(A[2]), .B2(n7), .ZN(n124) );
  AOI22_X1 U39 ( .A1(n4), .A2(n39), .B1(A[2]), .B2(n1), .ZN(n123) );
  OAI22_X1 U40 ( .A1(n113), .A2(n130), .B1(B[7]), .B2(n114), .ZN(S[7]) );
  INV_X1 U41 ( .A(B[7]), .ZN(n130) );
  AOI22_X1 U42 ( .A1(n4), .A2(n34), .B1(A[7]), .B2(n1), .ZN(n113) );
  AOI22_X1 U43 ( .A1(OP[0]), .A2(n34), .B1(A[7]), .B2(n7), .ZN(n114) );
  OAI22_X1 U44 ( .A1(n95), .A2(n57), .B1(B[16]), .B2(n96), .ZN(S[16]) );
  INV_X1 U45 ( .A(B[16]), .ZN(n57) );
  AOI22_X1 U46 ( .A1(OP[0]), .A2(n25), .B1(A[16]), .B2(n8), .ZN(n96) );
  AOI22_X1 U47 ( .A1(n5), .A2(n25), .B1(A[16]), .B2(n2), .ZN(n95) );
  OAI22_X1 U48 ( .A1(n93), .A2(n56), .B1(B[17]), .B2(n94), .ZN(S[17]) );
  INV_X1 U49 ( .A(B[17]), .ZN(n56) );
  AOI22_X1 U50 ( .A1(OP[0]), .A2(n24), .B1(A[17]), .B2(n8), .ZN(n94) );
  AOI22_X1 U51 ( .A1(n5), .A2(n24), .B1(A[17]), .B2(n2), .ZN(n93) );
  OAI22_X1 U52 ( .A1(n91), .A2(n55), .B1(B[18]), .B2(n92), .ZN(S[18]) );
  INV_X1 U53 ( .A(B[18]), .ZN(n55) );
  AOI22_X1 U54 ( .A1(OP[0]), .A2(n23), .B1(A[18]), .B2(n8), .ZN(n92) );
  AOI22_X1 U55 ( .A1(n5), .A2(n23), .B1(A[18]), .B2(n2), .ZN(n91) );
  OAI22_X1 U56 ( .A1(n89), .A2(n54), .B1(B[19]), .B2(n90), .ZN(S[19]) );
  INV_X1 U57 ( .A(B[19]), .ZN(n54) );
  AOI22_X1 U58 ( .A1(OP[0]), .A2(n22), .B1(A[19]), .B2(n8), .ZN(n90) );
  AOI22_X1 U59 ( .A1(n5), .A2(n22), .B1(A[19]), .B2(n2), .ZN(n89) );
  OAI22_X1 U60 ( .A1(n111), .A2(n129), .B1(B[8]), .B2(n112), .ZN(S[8]) );
  INV_X1 U61 ( .A(B[8]), .ZN(n129) );
  AOI22_X1 U62 ( .A1(n4), .A2(n33), .B1(A[8]), .B2(n1), .ZN(n111) );
  AOI22_X1 U63 ( .A1(OP[0]), .A2(n33), .B1(A[8]), .B2(n7), .ZN(n112) );
  OAI22_X1 U64 ( .A1(n115), .A2(n131), .B1(B[6]), .B2(n116), .ZN(S[6]) );
  INV_X1 U65 ( .A(B[6]), .ZN(n131) );
  AOI22_X1 U66 ( .A1(n4), .A2(n35), .B1(A[6]), .B2(n1), .ZN(n115) );
  AOI22_X1 U67 ( .A1(OP[0]), .A2(n35), .B1(A[6]), .B2(n7), .ZN(n116) );
  OAI22_X1 U68 ( .A1(n117), .A2(n132), .B1(B[5]), .B2(n118), .ZN(S[5]) );
  INV_X1 U69 ( .A(B[5]), .ZN(n132) );
  OAI22_X1 U70 ( .A1(n109), .A2(n64), .B1(B[9]), .B2(n110), .ZN(S[9]) );
  INV_X1 U71 ( .A(B[9]), .ZN(n64) );
  AOI22_X1 U72 ( .A1(OP[0]), .A2(n32), .B1(A[9]), .B2(n7), .ZN(n110) );
  AOI22_X1 U73 ( .A1(n4), .A2(n32), .B1(A[9]), .B2(n1), .ZN(n109) );
  OAI22_X1 U74 ( .A1(n107), .A2(n63), .B1(B[10]), .B2(n108), .ZN(S[10]) );
  INV_X1 U75 ( .A(B[10]), .ZN(n63) );
  AOI22_X1 U76 ( .A1(n4), .A2(n31), .B1(A[10]), .B2(n1), .ZN(n107) );
  AOI22_X1 U77 ( .A1(OP[0]), .A2(n31), .B1(A[10]), .B2(n7), .ZN(n108) );
  OAI22_X1 U78 ( .A1(n105), .A2(n62), .B1(B[11]), .B2(n106), .ZN(S[11]) );
  INV_X1 U79 ( .A(B[11]), .ZN(n62) );
  AOI22_X1 U80 ( .A1(n5), .A2(n30), .B1(A[11]), .B2(n1), .ZN(n105) );
  AOI22_X1 U81 ( .A1(OP[0]), .A2(n30), .B1(A[11]), .B2(n7), .ZN(n106) );
  OAI22_X1 U82 ( .A1(n103), .A2(n61), .B1(B[12]), .B2(n104), .ZN(S[12]) );
  INV_X1 U83 ( .A(B[12]), .ZN(n61) );
  AOI22_X1 U84 ( .A1(n5), .A2(n29), .B1(A[12]), .B2(n2), .ZN(n103) );
  AOI22_X1 U85 ( .A1(OP[0]), .A2(n29), .B1(A[12]), .B2(n8), .ZN(n104) );
  OAI22_X1 U86 ( .A1(n101), .A2(n60), .B1(B[13]), .B2(n102), .ZN(S[13]) );
  INV_X1 U87 ( .A(B[13]), .ZN(n60) );
  AOI22_X1 U88 ( .A1(n5), .A2(n28), .B1(A[13]), .B2(n2), .ZN(n101) );
  AOI22_X1 U89 ( .A1(OP[0]), .A2(n28), .B1(A[13]), .B2(n8), .ZN(n102) );
  OAI22_X1 U90 ( .A1(n99), .A2(n59), .B1(B[14]), .B2(n100), .ZN(S[14]) );
  INV_X1 U91 ( .A(B[14]), .ZN(n59) );
  AOI22_X1 U92 ( .A1(n5), .A2(n27), .B1(A[14]), .B2(n2), .ZN(n99) );
  AOI22_X1 U93 ( .A1(OP[0]), .A2(n27), .B1(A[14]), .B2(n8), .ZN(n100) );
  OAI22_X1 U94 ( .A1(n97), .A2(n58), .B1(B[15]), .B2(n98), .ZN(S[15]) );
  INV_X1 U95 ( .A(B[15]), .ZN(n58) );
  AOI22_X1 U96 ( .A1(n5), .A2(n26), .B1(A[15]), .B2(n2), .ZN(n97) );
  AOI22_X1 U97 ( .A1(OP[0]), .A2(n26), .B1(A[15]), .B2(n8), .ZN(n98) );
  OAI22_X1 U98 ( .A1(n87), .A2(n53), .B1(B[20]), .B2(n88), .ZN(S[20]) );
  INV_X1 U99 ( .A(B[20]), .ZN(n53) );
  AOI22_X1 U100 ( .A1(OP[0]), .A2(n21), .B1(A[20]), .B2(n8), .ZN(n88) );
  AOI22_X1 U101 ( .A1(n5), .A2(n21), .B1(A[20]), .B2(n2), .ZN(n87) );
  OAI22_X1 U102 ( .A1(n85), .A2(n52), .B1(B[21]), .B2(n86), .ZN(S[21]) );
  INV_X1 U103 ( .A(B[21]), .ZN(n52) );
  AOI22_X1 U104 ( .A1(OP[0]), .A2(n20), .B1(A[21]), .B2(n8), .ZN(n86) );
  AOI22_X1 U105 ( .A1(n5), .A2(n20), .B1(A[21]), .B2(n2), .ZN(n85) );
  OAI22_X1 U106 ( .A1(n83), .A2(n51), .B1(B[22]), .B2(n84), .ZN(S[22]) );
  INV_X1 U107 ( .A(B[22]), .ZN(n51) );
  AOI22_X1 U108 ( .A1(OP[0]), .A2(n19), .B1(A[22]), .B2(n8), .ZN(n84) );
  AOI22_X1 U109 ( .A1(n6), .A2(n19), .B1(A[22]), .B2(n2), .ZN(n83) );
  OAI22_X1 U110 ( .A1(n81), .A2(n50), .B1(B[23]), .B2(n82), .ZN(S[23]) );
  INV_X1 U111 ( .A(B[23]), .ZN(n50) );
  AOI22_X1 U112 ( .A1(OP[0]), .A2(n18), .B1(A[23]), .B2(n8), .ZN(n82) );
  AOI22_X1 U113 ( .A1(n6), .A2(n18), .B1(A[23]), .B2(n2), .ZN(n81) );
  OAI22_X1 U114 ( .A1(n121), .A2(n134), .B1(B[3]), .B2(n122), .ZN(S[3]) );
  INV_X1 U115 ( .A(B[3]), .ZN(n134) );
  AOI22_X1 U116 ( .A1(OP[0]), .A2(n38), .B1(A[3]), .B2(n7), .ZN(n122) );
  AOI22_X1 U117 ( .A1(n4), .A2(n38), .B1(A[3]), .B2(n1), .ZN(n121) );
  OAI22_X1 U118 ( .A1(n67), .A2(n43), .B1(B[30]), .B2(n68), .ZN(S[30]) );
  INV_X1 U119 ( .A(B[30]), .ZN(n43) );
  AOI22_X1 U120 ( .A1(OP[0]), .A2(n11), .B1(A[30]), .B2(n9), .ZN(n68) );
  AOI22_X1 U121 ( .A1(n6), .A2(n11), .B1(A[30]), .B2(n3), .ZN(n67) );
  OAI22_X1 U122 ( .A1(n79), .A2(n49), .B1(B[24]), .B2(n80), .ZN(S[24]) );
  INV_X1 U123 ( .A(B[24]), .ZN(n49) );
  AOI22_X1 U124 ( .A1(OP[0]), .A2(n17), .B1(A[24]), .B2(n9), .ZN(n80) );
  AOI22_X1 U125 ( .A1(n6), .A2(n17), .B1(A[24]), .B2(n3), .ZN(n79) );
  OAI22_X1 U126 ( .A1(n75), .A2(n47), .B1(B[26]), .B2(n76), .ZN(S[26]) );
  INV_X1 U127 ( .A(B[26]), .ZN(n47) );
  AOI22_X1 U128 ( .A1(OP[0]), .A2(n15), .B1(A[26]), .B2(n9), .ZN(n76) );
  AOI22_X1 U129 ( .A1(n6), .A2(n15), .B1(A[26]), .B2(n3), .ZN(n75) );
  OAI22_X1 U130 ( .A1(n73), .A2(n46), .B1(B[27]), .B2(n74), .ZN(S[27]) );
  INV_X1 U131 ( .A(B[27]), .ZN(n46) );
  AOI22_X1 U132 ( .A1(OP[0]), .A2(n14), .B1(A[27]), .B2(n9), .ZN(n74) );
  AOI22_X1 U133 ( .A1(n6), .A2(n14), .B1(A[27]), .B2(n3), .ZN(n73) );
  OAI22_X1 U134 ( .A1(n69), .A2(n44), .B1(B[29]), .B2(n70), .ZN(S[29]) );
  INV_X1 U135 ( .A(B[29]), .ZN(n44) );
  AOI22_X1 U136 ( .A1(OP[0]), .A2(n12), .B1(A[29]), .B2(n9), .ZN(n70) );
  AOI22_X1 U137 ( .A1(n6), .A2(n12), .B1(A[29]), .B2(n3), .ZN(n69) );
  OAI22_X1 U138 ( .A1(n77), .A2(n48), .B1(B[25]), .B2(n78), .ZN(S[25]) );
  INV_X1 U139 ( .A(B[25]), .ZN(n48) );
  AOI22_X1 U140 ( .A1(OP[0]), .A2(n16), .B1(A[25]), .B2(n9), .ZN(n78) );
  AOI22_X1 U141 ( .A1(n6), .A2(n16), .B1(A[25]), .B2(n3), .ZN(n77) );
  OAI22_X1 U142 ( .A1(n71), .A2(n45), .B1(B[28]), .B2(n72), .ZN(S[28]) );
  INV_X1 U143 ( .A(B[28]), .ZN(n45) );
  AOI22_X1 U144 ( .A1(OP[0]), .A2(n13), .B1(A[28]), .B2(n9), .ZN(n72) );
  AOI22_X1 U145 ( .A1(n6), .A2(n13), .B1(A[28]), .B2(n3), .ZN(n71) );
  OAI22_X1 U146 ( .A1(n65), .A2(n42), .B1(B[31]), .B2(n66), .ZN(S[31]) );
  INV_X1 U147 ( .A(B[31]), .ZN(n42) );
  AOI22_X1 U148 ( .A1(OP[0]), .A2(n10), .B1(n9), .B2(A[31]), .ZN(n66) );
  AOI22_X1 U149 ( .A1(n6), .A2(n10), .B1(n3), .B2(A[31]), .ZN(n65) );
  AOI22_X1 U150 ( .A1(n4), .A2(n36), .B1(A[5]), .B2(n1), .ZN(n117) );
  AOI22_X1 U151 ( .A1(OP[0]), .A2(n36), .B1(A[5]), .B2(n7), .ZN(n118) );
  INV_X1 U152 ( .A(A[5]), .ZN(n36) );
  AOI22_X1 U153 ( .A1(n4), .A2(n40), .B1(A[1]), .B2(n1), .ZN(n125) );
  AOI22_X1 U154 ( .A1(OP[0]), .A2(n40), .B1(A[1]), .B2(n7), .ZN(n126) );
  INV_X1 U155 ( .A(A[1]), .ZN(n40) );
  OAI22_X1 U156 ( .A1(n123), .A2(n135), .B1(B[2]), .B2(n124), .ZN(S[2]) );
  INV_X1 U157 ( .A(B[2]), .ZN(n135) );
  AOI22_X1 U158 ( .A1(n4), .A2(n37), .B1(A[4]), .B2(n1), .ZN(n119) );
  AOI22_X1 U159 ( .A1(OP[0]), .A2(n37), .B1(A[4]), .B2(n7), .ZN(n120) );
  INV_X1 U160 ( .A(A[4]), .ZN(n37) );
  AOI22_X1 U161 ( .A1(OP[0]), .A2(n41), .B1(A[0]), .B2(n7), .ZN(n128) );
  AOI22_X1 U162 ( .A1(n4), .A2(n41), .B1(A[0]), .B2(n1), .ZN(n127) );
  INV_X1 U163 ( .A(A[0]), .ZN(n41) );
  OAI22_X1 U164 ( .A1(n127), .A2(n137), .B1(B[0]), .B2(n128), .ZN(S[0]) );
  INV_X1 U165 ( .A(B[0]), .ZN(n137) );
  OAI22_X1 U166 ( .A1(n119), .A2(n133), .B1(B[4]), .B2(n120), .ZN(S[4]) );
  INV_X1 U167 ( .A(B[4]), .ZN(n133) );
  OAI22_X1 U168 ( .A1(n125), .A2(n136), .B1(B[1]), .B2(n126), .ZN(S[1]) );
  INV_X1 U169 ( .A(B[1]), .ZN(n136) );
endmodule


module MASK_GEN_DATA_W32_MASK_SIZE41_1 ( OP, A, MASK0, MASK8, MASK16, MASK24, 
        MSB );
  input [1:0] OP;
  input [31:0] A;
  output [40:0] MASK0;
  output [40:0] MASK8;
  output [40:0] MASK16;
  output [40:0] MASK24;
  output MSB;
  wire   n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, \MASK16[40] , n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48,
         \MASK8[15] , n50, \MASK8[14] , n52, \MASK8[13] , n76, \MASK8[12] ,
         n78, \MASK8[11] , n80, \MASK8[10] , n82, \MASK8[9] , n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n99, n100,
         n101;
  assign MASK24[0] = 1'b0;
  assign MASK16[0] = 1'b0;
  assign MASK8[0] = 1'b0;
  assign MASK0[0] = 1'b0;
  assign MASK16[39] = MASK8[31];
  assign MASK16[38] = MASK8[30];
  assign MASK16[37] = MASK8[29];
  assign MASK16[36] = MASK8[28];
  assign MASK16[35] = MASK8[27];
  assign MASK16[34] = MASK8[26];
  assign MASK16[33] = MASK8[25];
  assign MASK24[39] = MASK16[31];
  assign MASK24[38] = MASK16[30];
  assign MASK24[37] = MASK16[29];
  assign MASK24[36] = MASK16[28];
  assign MASK24[35] = MASK16[27];
  assign MASK24[34] = MASK16[26];
  assign MASK24[33] = MASK16[25];
  assign MASK24[32] = MASK16[24];
  assign MASK24[8] = MASK16[16];
  assign MASK24[7] = MASK16[15];
  assign MASK24[6] = MASK16[14];
  assign MASK24[5] = MASK16[13];
  assign MASK24[4] = MASK16[12];
  assign MASK24[3] = MASK16[11];
  assign MASK24[2] = MASK16[10];
  assign MASK24[1] = MASK16[9];
  assign MASK24[15] = \MASK16[40] ;
  assign MASK24[13] = \MASK16[40] ;
  assign MASK24[29] = \MASK16[40] ;
  assign MASK24[30] = \MASK16[40] ;
  assign MASK24[14] = \MASK16[40] ;
  assign MASK24[11] = \MASK16[40] ;
  assign MASK24[31] = \MASK16[40] ;
  assign MASK16[17] = \MASK16[40] ;
  assign MASK16[18] = \MASK16[40] ;
  assign MASK24[19] = \MASK16[40] ;
  assign MASK24[20] = \MASK16[40] ;
  assign MASK24[21] = \MASK16[40] ;
  assign MASK24[22] = \MASK16[40] ;
  assign MASK24[24] = \MASK16[40] ;
  assign MASK24[16] = \MASK16[40] ;
  assign MASK24[26] = \MASK16[40] ;
  assign MASK0[40] = \MASK16[40] ;
  assign MASK24[10] = \MASK16[40] ;
  assign MASK24[18] = \MASK16[40] ;
  assign MASK24[28] = \MASK16[40] ;
  assign MASK24[23] = \MASK16[40] ;
  assign MASK24[12] = \MASK16[40] ;
  assign MASK8[40] = \MASK16[40] ;
  assign MASK24[17] = \MASK16[40] ;
  assign MASK24[9] = \MASK16[40] ;
  assign MASK24[25] = \MASK16[40] ;
  assign MASK24[27] = \MASK16[40] ;
  assign MASK24[40] = \MASK16[40] ;
  assign MASK16[19] = \MASK16[40] ;
  assign MASK16[20] = \MASK16[40] ;
  assign MASK16[21] = \MASK16[40] ;
  assign MASK16[22] = \MASK16[40] ;
  assign MASK16[23] = \MASK16[40] ;
  assign MASK16[40] = \MASK16[40] ;
  assign MASK16[7] = \MASK8[15] ;
  assign MASK8[15] = \MASK8[15] ;
  assign MASK16[6] = \MASK8[14] ;
  assign MASK8[14] = \MASK8[14] ;
  assign MASK16[5] = \MASK8[13] ;
  assign MASK8[13] = \MASK8[13] ;
  assign MASK16[4] = \MASK8[12] ;
  assign MASK8[12] = \MASK8[12] ;
  assign MASK16[3] = \MASK8[11] ;
  assign MASK8[11] = \MASK8[11] ;
  assign MASK16[2] = \MASK8[10] ;
  assign MASK8[10] = \MASK8[10] ;
  assign MASK16[1] = \MASK8[9] ;
  assign MASK8[9] = \MASK8[9] ;

  BUF_X1 U2 ( .A(n15), .Z(n29) );
  INV_X2 U3 ( .A(n1), .ZN(n2) );
  INV_X1 U4 ( .A(n29), .ZN(MSB) );
  AOI21_X1 U5 ( .B1(n100), .B2(OP[0]), .A(n74), .ZN(n73) );
  INV_X1 U6 ( .A(n73), .ZN(n1) );
  INV_X1 U7 ( .A(n1), .ZN(n3) );
  INV_X1 U8 ( .A(n2), .ZN(n4) );
  INV_X1 U9 ( .A(n2), .ZN(n5) );
  NOR2_X1 U10 ( .A1(n100), .A2(OP[0]), .ZN(n74) );
  BUF_X2 U11 ( .A(n6), .Z(n9) );
  INV_X2 U12 ( .A(n29), .ZN(\MASK16[40] ) );
  CLKBUF_X1 U13 ( .A(n15), .Z(n28) );
  CLKBUF_X1 U14 ( .A(n101), .Z(n7) );
  CLKBUF_X1 U15 ( .A(n16), .Z(n14) );
  CLKBUF_X1 U16 ( .A(n53), .Z(n16) );
  BUF_X1 U17 ( .A(n6), .Z(n8) );
  BUF_X1 U18 ( .A(n7), .Z(n10) );
  BUF_X1 U19 ( .A(n7), .Z(n11) );
  BUF_X1 U20 ( .A(n13), .Z(n22) );
  BUF_X1 U21 ( .A(n13), .Z(n23) );
  BUF_X1 U22 ( .A(n12), .Z(n21) );
  BUF_X1 U23 ( .A(n14), .Z(n25) );
  BUF_X1 U24 ( .A(n12), .Z(n19) );
  BUF_X1 U25 ( .A(n12), .Z(n20) );
  BUF_X1 U26 ( .A(n13), .Z(n24) );
  BUF_X1 U27 ( .A(n14), .Z(n26) );
  BUF_X1 U28 ( .A(n14), .Z(n27) );
  BUF_X1 U29 ( .A(n101), .Z(n6) );
  NAND2_X1 U30 ( .A1(n27), .A2(n64), .ZN(MASK16[24]) );
  NAND2_X1 U31 ( .A1(n29), .A2(n61), .ZN(MASK16[26]) );
  NAND2_X1 U32 ( .A1(n27), .A2(n60), .ZN(MASK16[27]) );
  INV_X1 U33 ( .A(MASK16[16]), .ZN(n30) );
  INV_X1 U34 ( .A(MASK16[15]), .ZN(n32) );
  INV_X1 U35 ( .A(MASK16[14]), .ZN(n34) );
  INV_X1 U36 ( .A(MASK16[13]), .ZN(n36) );
  INV_X1 U37 ( .A(MASK16[12]), .ZN(n38) );
  INV_X1 U38 ( .A(MASK16[11]), .ZN(n40) );
  INV_X1 U39 ( .A(MASK16[10]), .ZN(n42) );
  INV_X1 U40 ( .A(MASK16[9]), .ZN(n44) );
  NAND2_X1 U41 ( .A1(n42), .A2(n61), .ZN(MASK8[18]) );
  NAND2_X1 U42 ( .A1(n96), .A2(n61), .ZN(MASK0[10]) );
  INV_X1 U43 ( .A(MASK8[2]), .ZN(n96) );
  INV_X1 U44 ( .A(n72), .ZN(n101) );
  NAND2_X1 U45 ( .A1(n40), .A2(n60), .ZN(MASK8[19]) );
  NAND2_X1 U46 ( .A1(n94), .A2(n60), .ZN(MASK0[11]) );
  INV_X1 U47 ( .A(MASK8[3]), .ZN(n94) );
  BUF_X1 U48 ( .A(n16), .Z(n13) );
  BUF_X1 U49 ( .A(n16), .Z(n12) );
  BUF_X1 U50 ( .A(n53), .Z(n15) );
  NOR2_X1 U51 ( .A1(OP[0]), .A2(OP[1]), .ZN(n72) );
  OAI21_X1 U52 ( .B1(n10), .B2(n33), .A(n24), .ZN(MASK0[38]) );
  OAI21_X1 U53 ( .B1(n9), .B2(n50), .A(n19), .ZN(MASK8[37]) );
  OAI21_X1 U54 ( .B1(n9), .B2(n52), .A(n19), .ZN(MASK8[36]) );
  OAI21_X1 U55 ( .B1(n31), .B2(n8), .A(n24), .ZN(MASK0[39]) );
  NOR2_X1 U56 ( .A1(n41), .A2(n2), .ZN(MASK16[11]) );
  NOR2_X1 U57 ( .A1(n45), .A2(n2), .ZN(MASK16[9]) );
  NOR2_X1 U58 ( .A1(n31), .A2(n3), .ZN(MASK16[16]) );
  NOR2_X1 U59 ( .A1(n33), .A2(n3), .ZN(MASK16[15]) );
  NOR2_X1 U60 ( .A1(n35), .A2(n2), .ZN(MASK16[14]) );
  NOR2_X1 U61 ( .A1(n39), .A2(n2), .ZN(MASK16[12]) );
  NOR2_X1 U62 ( .A1(n43), .A2(n3), .ZN(MASK16[10]) );
  NOR2_X1 U63 ( .A1(n37), .A2(n3), .ZN(MASK16[13]) );
  NAND2_X1 U64 ( .A1(A[2]), .A2(n72), .ZN(n61) );
  OAI21_X1 U65 ( .B1(n95), .B2(n9), .A(n23), .ZN(MASK8[26]) );
  OAI21_X1 U66 ( .B1(n93), .B2(n9), .A(n22), .ZN(MASK8[27]) );
  OAI21_X1 U67 ( .B1(n89), .B2(n9), .A(n22), .ZN(MASK8[29]) );
  OAI21_X1 U68 ( .B1(n91), .B2(n8), .A(n22), .ZN(MASK8[28]) );
  OAI21_X1 U69 ( .B1(n87), .B2(n8), .A(n21), .ZN(MASK8[30]) );
  OAI21_X1 U70 ( .B1(n85), .B2(n8), .A(n21), .ZN(MASK8[31]) );
  OAI21_X1 U71 ( .B1(n9), .B2(n97), .A(n23), .ZN(MASK8[25]) );
  NOR2_X1 U72 ( .A1(n95), .A2(n3), .ZN(MASK8[3]) );
  NOR2_X1 U73 ( .A1(n89), .A2(n3), .ZN(MASK8[6]) );
  NOR2_X1 U74 ( .A1(n87), .A2(n3), .ZN(MASK8[7]) );
  NOR2_X1 U75 ( .A1(n97), .A2(n2), .ZN(MASK8[2]) );
  NOR2_X1 U76 ( .A1(n91), .A2(n3), .ZN(MASK8[5]) );
  NOR2_X1 U77 ( .A1(n93), .A2(n2), .ZN(MASK8[4]) );
  NOR2_X1 U78 ( .A1(n85), .A2(n2), .ZN(MASK8[8]) );
  OAI21_X1 U79 ( .B1(n82), .B2(n8), .A(n21), .ZN(MASK8[32]) );
  OAI21_X1 U80 ( .B1(n85), .B2(n8), .A(n65), .ZN(MASK0[23]) );
  OAI21_X1 U81 ( .B1(n87), .B2(n8), .A(n66), .ZN(MASK0[22]) );
  OAI21_X1 U82 ( .B1(n89), .B2(n8), .A(n67), .ZN(MASK0[21]) );
  OAI21_X1 U83 ( .B1(n93), .B2(n8), .A(n69), .ZN(MASK0[19]) );
  OAI21_X1 U84 ( .B1(n91), .B2(n8), .A(n68), .ZN(MASK0[20]) );
  OAI21_X1 U85 ( .B1(n95), .B2(n8), .A(n70), .ZN(MASK0[18]) );
  OAI21_X1 U86 ( .B1(n9), .B2(n80), .A(n20), .ZN(MASK8[33]) );
  OAI21_X1 U87 ( .B1(n9), .B2(n78), .A(n20), .ZN(MASK8[34]) );
  OAI21_X1 U88 ( .B1(n9), .B2(n76), .A(n20), .ZN(MASK8[35]) );
  OAI21_X1 U89 ( .B1(n9), .B2(n48), .A(n19), .ZN(MASK8[38]) );
  OAI21_X1 U90 ( .B1(n9), .B2(n46), .A(n23), .ZN(MASK8[39]) );
  OAI21_X1 U91 ( .B1(n82), .B2(n8), .A(n63), .ZN(MASK0[24]) );
  OAI21_X1 U92 ( .B1(n9), .B2(n97), .A(n71), .ZN(MASK0[17]) );
  NAND2_X1 U93 ( .A1(A[3]), .A2(n72), .ZN(n60) );
  OAI21_X1 U94 ( .B1(n10), .B2(n52), .A(n38), .ZN(MASK0[28]) );
  OAI21_X1 U95 ( .B1(n10), .B2(n46), .A(n32), .ZN(MASK0[31]) );
  OAI21_X1 U96 ( .B1(n10), .B2(n76), .A(n40), .ZN(MASK0[27]) );
  OAI21_X1 U97 ( .B1(n10), .B2(n48), .A(n34), .ZN(MASK0[30]) );
  OAI21_X1 U98 ( .B1(n10), .B2(n50), .A(n36), .ZN(MASK0[29]) );
  OAI21_X1 U99 ( .B1(n11), .B2(n78), .A(n42), .ZN(MASK0[26]) );
  OAI21_X1 U100 ( .B1(n11), .B2(n80), .A(n44), .ZN(MASK0[25]) );
  OAI21_X1 U101 ( .B1(n10), .B2(n45), .A(n30), .ZN(MASK0[32]) );
  OAI21_X1 U102 ( .B1(n10), .B2(n35), .A(n25), .ZN(MASK0[37]) );
  OAI21_X1 U103 ( .B1(n10), .B2(n41), .A(n26), .ZN(MASK0[34]) );
  OAI21_X1 U104 ( .B1(n10), .B2(n43), .A(n25), .ZN(MASK0[33]) );
  OAI21_X1 U105 ( .B1(n10), .B2(n37), .A(n24), .ZN(MASK0[36]) );
  NAND2_X1 U106 ( .A1(n26), .A2(n58), .ZN(MASK16[28]) );
  NAND2_X1 U107 ( .A1(n28), .A2(n57), .ZN(MASK16[29]) );
  NAND2_X1 U108 ( .A1(n27), .A2(n62), .ZN(MASK16[25]) );
  NAND2_X1 U109 ( .A1(n28), .A2(n55), .ZN(MASK16[31]) );
  NAND2_X1 U110 ( .A1(n26), .A2(n56), .ZN(MASK16[30]) );
  INV_X1 U111 ( .A(OP[1]), .ZN(n100) );
  NAND2_X1 U112 ( .A1(n36), .A2(n57), .ZN(MASK8[21]) );
  NAND2_X1 U113 ( .A1(n38), .A2(n58), .ZN(MASK8[20]) );
  NAND2_X1 U114 ( .A1(n92), .A2(n58), .ZN(MASK0[12]) );
  INV_X1 U115 ( .A(MASK8[4]), .ZN(n92) );
  NAND2_X1 U116 ( .A1(n90), .A2(n57), .ZN(MASK0[13]) );
  INV_X1 U117 ( .A(MASK8[5]), .ZN(n90) );
  NAND2_X1 U118 ( .A1(n44), .A2(n62), .ZN(MASK8[17]) );
  INV_X1 U119 ( .A(n71), .ZN(\MASK8[9] ) );
  INV_X1 U120 ( .A(n69), .ZN(\MASK8[11] ) );
  INV_X1 U121 ( .A(n66), .ZN(\MASK8[14] ) );
  INV_X1 U122 ( .A(n65), .ZN(\MASK8[15] ) );
  INV_X1 U123 ( .A(n70), .ZN(\MASK8[10] ) );
  INV_X1 U124 ( .A(n67), .ZN(\MASK8[13] ) );
  INV_X1 U125 ( .A(n68), .ZN(\MASK8[12] ) );
  NAND2_X1 U126 ( .A1(n59), .A2(n62), .ZN(MASK0[9]) );
  NAND2_X1 U127 ( .A1(n28), .A2(n54), .ZN(MASK16[32]) );
  NAND2_X1 U128 ( .A1(n32), .A2(n55), .ZN(MASK8[23]) );
  NAND2_X1 U129 ( .A1(n30), .A2(n54), .ZN(MASK8[24]) );
  NAND2_X1 U130 ( .A1(n34), .A2(n56), .ZN(MASK8[22]) );
  NAND2_X1 U131 ( .A1(n86), .A2(n55), .ZN(MASK0[15]) );
  INV_X1 U132 ( .A(MASK8[7]), .ZN(n86) );
  NAND2_X1 U133 ( .A1(n84), .A2(n54), .ZN(MASK0[16]) );
  INV_X1 U134 ( .A(MASK8[8]), .ZN(n84) );
  NAND2_X1 U135 ( .A1(n88), .A2(n56), .ZN(MASK0[14]) );
  INV_X1 U136 ( .A(MASK8[6]), .ZN(n88) );
  NAND2_X1 U137 ( .A1(n63), .A2(n64), .ZN(MASK8[16]) );
  OAI21_X1 U138 ( .B1(n10), .B2(n39), .A(n25), .ZN(MASK0[35]) );
  INV_X1 U139 ( .A(n63), .ZN(MASK16[8]) );
  INV_X1 U140 ( .A(n59), .ZN(MASK8[1]) );
  AND2_X1 U141 ( .A1(n5), .A2(A[2]), .ZN(MASK0[3]) );
  AND2_X1 U142 ( .A1(n4), .A2(A[3]), .ZN(MASK0[4]) );
  NAND2_X1 U143 ( .A1(A[7]), .A2(n72), .ZN(n55) );
  NAND2_X1 U144 ( .A1(A[8]), .A2(n72), .ZN(n54) );
  NAND2_X1 U145 ( .A1(A[6]), .A2(n72), .ZN(n56) );
  NAND2_X1 U146 ( .A1(A[23]), .A2(n1), .ZN(n63) );
  NAND2_X1 U147 ( .A1(A[16]), .A2(n4), .ZN(n71) );
  NAND2_X1 U148 ( .A1(A[18]), .A2(n1), .ZN(n69) );
  NAND2_X1 U149 ( .A1(A[21]), .A2(n5), .ZN(n66) );
  NAND2_X1 U150 ( .A1(A[22]), .A2(n1), .ZN(n65) );
  NAND2_X1 U151 ( .A1(A[17]), .A2(n5), .ZN(n70) );
  NAND2_X1 U152 ( .A1(A[20]), .A2(n4), .ZN(n67) );
  NAND2_X1 U153 ( .A1(A[19]), .A2(n1), .ZN(n68) );
  NAND2_X1 U154 ( .A1(A[8]), .A2(n5), .ZN(n59) );
  OAI21_X1 U155 ( .B1(n2), .B2(n99), .A(n64), .ZN(MASK0[8]) );
  INV_X1 U156 ( .A(A[7]), .ZN(n99) );
  NAND2_X1 U157 ( .A1(A[31]), .A2(n74), .ZN(n53) );
  INV_X1 U158 ( .A(A[9]), .ZN(n97) );
  INV_X1 U159 ( .A(A[10]), .ZN(n95) );
  INV_X1 U160 ( .A(A[13]), .ZN(n89) );
  INV_X1 U161 ( .A(A[14]), .ZN(n87) );
  INV_X1 U162 ( .A(A[11]), .ZN(n93) );
  INV_X1 U163 ( .A(A[12]), .ZN(n91) );
  INV_X1 U164 ( .A(A[15]), .ZN(n85) );
  INV_X1 U165 ( .A(A[31]), .ZN(n31) );
  INV_X1 U166 ( .A(A[30]), .ZN(n33) );
  INV_X1 U167 ( .A(A[21]), .ZN(n50) );
  INV_X1 U168 ( .A(A[20]), .ZN(n52) );
  INV_X1 U169 ( .A(A[18]), .ZN(n78) );
  INV_X1 U170 ( .A(A[17]), .ZN(n80) );
  INV_X1 U171 ( .A(A[19]), .ZN(n76) );
  INV_X1 U172 ( .A(A[23]), .ZN(n46) );
  INV_X1 U173 ( .A(A[22]), .ZN(n48) );
  INV_X1 U174 ( .A(A[16]), .ZN(n82) );
  INV_X1 U175 ( .A(A[27]), .ZN(n39) );
  INV_X1 U176 ( .A(A[29]), .ZN(n35) );
  INV_X1 U177 ( .A(A[24]), .ZN(n45) );
  INV_X1 U178 ( .A(A[26]), .ZN(n41) );
  INV_X1 U179 ( .A(A[25]), .ZN(n43) );
  INV_X1 U180 ( .A(A[28]), .ZN(n37) );
  AND2_X1 U181 ( .A1(n4), .A2(A[6]), .ZN(MASK0[7]) );
  AND2_X1 U182 ( .A1(n5), .A2(A[5]), .ZN(MASK0[6]) );
  NAND2_X1 U183 ( .A1(A[5]), .A2(n72), .ZN(n57) );
  AND2_X1 U184 ( .A1(n5), .A2(A[1]), .ZN(MASK0[2]) );
  NAND2_X1 U185 ( .A1(A[1]), .A2(n72), .ZN(n62) );
  AND2_X1 U186 ( .A1(n4), .A2(A[4]), .ZN(MASK0[5]) );
  NAND2_X1 U187 ( .A1(A[4]), .A2(n72), .ZN(n58) );
  NAND2_X1 U188 ( .A1(A[0]), .A2(n72), .ZN(n64) );
  AND2_X1 U189 ( .A1(n4), .A2(A[0]), .ZN(MASK0[1]) );
endmodule


module COARSE_SHIFT_DATA_W32_MASK_SIZE41_1 ( MASK0, MASK8, MASK16, MASK24, MSB, 
        AMOUNT, S );
  input [40:0] MASK0;
  input [40:0] MASK8;
  input [40:0] MASK16;
  input [40:0] MASK24;
  input [28:0] AMOUNT;
  output [40:0] S;
  input MSB;
  wire   n5, n6, n7, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, net27110, net27102,
         net27116, net27114, net27112, net27128, net27126, net27124, net27142,
         net27140, net27138, net27136, net27144, net27154, net27152, net27150,
         net27148, net27156, net34755, net34754, net35591, net35590, net40402,
         net40444, net40443, n91, net40386, net34894, net34892, net24005, n92,
         n90, net34840, net34565, n99, n98, n97, n96, n95, n93, n101, net34852,
         net34646, net27158, net27146, net27134, net24008, net24007, net24006,
         n9, n11, n10, n1, n2, n3, n4, n8, n43, n94, n100, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189;

  BUF_X2 U1 ( .A(net27146), .Z(n43) );
  BUF_X1 U2 ( .A(net27146), .Z(net27140) );
  BUF_X1 U3 ( .A(net24007), .Z(net27144) );
  AOI221_X1 U4 ( .B1(MASK16[0]), .B2(n2), .C1(MASK8[0]), .C2(n1), .A(net27102), 
        .ZN(n89) );
  INV_X1 U5 ( .A(net34892), .ZN(n1) );
  BUF_X1 U6 ( .A(net27144), .Z(net35591) );
  BUF_X2 U7 ( .A(net27158), .Z(net27154) );
  BUF_X1 U8 ( .A(net27156), .Z(n2) );
  CLKBUF_X3 U9 ( .A(net27134), .Z(net27128) );
  AND2_X1 U10 ( .A1(AMOUNT[1]), .A2(net24005), .ZN(n3) );
  AND2_X1 U11 ( .A1(net24006), .A2(AMOUNT[0]), .ZN(n4) );
  NAND2_X1 U12 ( .A1(MASK16[30]), .A2(net27152), .ZN(n8) );
  BUF_X1 U13 ( .A(net27144), .Z(net27136) );
  BUF_X1 U14 ( .A(net27158), .Z(net27152) );
  AOI221_X1 U15 ( .B1(MASK16[40]), .B2(net40402), .C1(MASK8[40]), .C2(net27142), .A(net27102), .ZN(n21) );
  CLKBUF_X1 U16 ( .A(n92), .Z(net34894) );
  AND4_X2 U17 ( .A1(n110), .A2(net34892), .A3(net34894), .A4(MSB), .ZN(n94) );
  AND4_X2 U18 ( .A1(n110), .A2(net34892), .A3(net34894), .A4(MSB), .ZN(n100)
         );
  BUF_X1 U19 ( .A(net27156), .Z(net40443) );
  AND2_X1 U20 ( .A1(net40386), .A2(n110), .ZN(n102) );
  CLKBUF_X1 U21 ( .A(net27146), .Z(net27138) );
  AND2_X1 U22 ( .A1(net40386), .A2(n110), .ZN(n7) );
  BUF_X2 U23 ( .A(net24008), .Z(net27156) );
  AND2_X1 U24 ( .A1(MASK16[39]), .A2(net40402), .ZN(n103) );
  AND2_X1 U25 ( .A1(MASK8[39]), .A2(net27142), .ZN(n104) );
  NOR3_X1 U26 ( .A1(n103), .A2(n104), .A3(net34754), .ZN(n25) );
  CLKBUF_X3 U27 ( .A(net27158), .Z(net40402) );
  CLKBUF_X3 U28 ( .A(net27144), .Z(net27142) );
  BUF_X1 U29 ( .A(net27156), .Z(net40444) );
  INV_X1 U30 ( .A(AMOUNT[11]), .ZN(n105) );
  NAND2_X1 U31 ( .A1(n107), .A2(n105), .ZN(n106) );
  NOR2_X1 U32 ( .A1(AMOUNT[12]), .A2(AMOUNT[10]), .ZN(n107) );
  NOR2_X1 U33 ( .A1(n101), .A2(n106), .ZN(n108) );
  CLKBUF_X3 U34 ( .A(net34646), .Z(net27112) );
  BUF_X2 U35 ( .A(net27156), .Z(net27150) );
  BUF_X1 U36 ( .A(n9), .Z(net27134) );
  CLKBUF_X3 U37 ( .A(net27134), .Z(n109) );
  NOR2_X1 U38 ( .A1(n9), .A2(net34565), .ZN(n110) );
  CLKBUF_X3 U39 ( .A(net34646), .Z(net27114) );
  BUF_X1 U40 ( .A(net34565), .Z(net34646) );
  CLKBUF_X3 U41 ( .A(net27134), .Z(net27126) );
  OR2_X1 U42 ( .A1(AMOUNT[18]), .A2(AMOUNT[16]), .ZN(n111) );
  AND2_X1 U43 ( .A1(n112), .A2(n113), .ZN(n95) );
  NOR4_X1 U44 ( .A1(AMOUNT[20]), .A2(AMOUNT[19]), .A3(AMOUNT[21]), .A4(
        AMOUNT[22]), .ZN(n112) );
  NOR2_X1 U45 ( .A1(n111), .A2(AMOUNT[17]), .ZN(n113) );
  OR2_X1 U46 ( .A1(AMOUNT[25]), .A2(AMOUNT[23]), .ZN(n114) );
  NAND4_X1 U47 ( .A1(n115), .A2(n8), .A3(n116), .A4(n42), .ZN(S[30]) );
  INV_X1 U48 ( .A(n145), .ZN(n115) );
  INV_X1 U49 ( .A(net34754), .ZN(n116) );
  NOR3_X1 U50 ( .A1(n138), .A2(n137), .A3(n102), .ZN(n59) );
  NAND4_X1 U51 ( .A1(n117), .A2(n118), .A3(n119), .A4(n120), .ZN(n98) );
  INV_X1 U52 ( .A(AMOUNT[7]), .ZN(n117) );
  INV_X1 U53 ( .A(AMOUNT[6]), .ZN(n118) );
  INV_X1 U54 ( .A(AMOUNT[8]), .ZN(n119) );
  INV_X1 U55 ( .A(AMOUNT[9]), .ZN(n120) );
  NAND3_X1 U56 ( .A1(n123), .A2(n122), .A3(n121), .ZN(n101) );
  INV_X1 U57 ( .A(AMOUNT[15]), .ZN(n121) );
  INV_X1 U58 ( .A(AMOUNT[14]), .ZN(n122) );
  INV_X1 U59 ( .A(AMOUNT[13]), .ZN(n123) );
  NAND4_X1 U60 ( .A1(n124), .A2(n125), .A3(n126), .A4(n127), .ZN(n99) );
  INV_X1 U61 ( .A(AMOUNT[27]), .ZN(n124) );
  INV_X1 U62 ( .A(AMOUNT[26]), .ZN(n125) );
  INV_X1 U63 ( .A(AMOUNT[2]), .ZN(n126) );
  INV_X1 U64 ( .A(AMOUNT[28]), .ZN(n127) );
  NAND2_X1 U65 ( .A1(n11), .A2(n10), .ZN(S[8]) );
  AOI22_X1 U66 ( .A1(MASK24[8]), .A2(net27112), .B1(MASK0[8]), .B2(net27128), 
        .ZN(n10) );
  CLKBUF_X1 U67 ( .A(net27134), .Z(net27124) );
  CLKBUF_X3 U68 ( .A(net34646), .Z(net27116) );
  NOR3_X1 U69 ( .A1(net34755), .A2(n129), .A3(n128), .ZN(n11) );
  AND2_X1 U70 ( .A1(MASK8[8]), .A2(net27140), .ZN(n129) );
  BUF_X1 U71 ( .A(net24007), .Z(net27146) );
  INV_X1 U72 ( .A(n90), .ZN(net24007) );
  AND2_X1 U73 ( .A1(MASK16[8]), .A2(net27154), .ZN(n128) );
  BUF_X1 U74 ( .A(net24008), .Z(net27158) );
  INV_X1 U75 ( .A(n92), .ZN(net24008) );
  AND2_X1 U76 ( .A1(n93), .A2(net34852), .ZN(n9) );
  NOR2_X1 U77 ( .A1(n9), .A2(net34565), .ZN(n91) );
  AND2_X1 U78 ( .A1(net24005), .A2(net24006), .ZN(net34852) );
  INV_X1 U79 ( .A(AMOUNT[1]), .ZN(net24006) );
  INV_X1 U80 ( .A(AMOUNT[0]), .ZN(net24005) );
  AND2_X1 U81 ( .A1(n93), .A2(net34840), .ZN(net34565) );
  AND2_X1 U82 ( .A1(AMOUNT[0]), .A2(AMOUNT[1]), .ZN(net34840) );
  AND4_X2 U83 ( .A1(n97), .A2(n96), .A3(n95), .A4(n108), .ZN(n93) );
  NAND2_X1 U84 ( .A1(n93), .A2(n4), .ZN(n90) );
  NAND2_X1 U85 ( .A1(n93), .A2(n3), .ZN(n92) );
  NOR3_X1 U86 ( .A1(n99), .A2(n114), .A3(AMOUNT[24]), .ZN(n96) );
  NOR3_X1 U87 ( .A1(n98), .A2(AMOUNT[3]), .A3(n130), .ZN(n97) );
  OR2_X1 U88 ( .A1(AMOUNT[4]), .A2(AMOUNT[5]), .ZN(n130) );
  AND4_X2 U89 ( .A1(n91), .A2(n92), .A3(n90), .A4(MSB), .ZN(net34755) );
  AND3_X1 U90 ( .A1(n92), .A2(n90), .A3(MSB), .ZN(net40386) );
  CLKBUF_X1 U91 ( .A(n90), .Z(net34892) );
  AND4_X2 U92 ( .A1(n110), .A2(net34892), .A3(net34894), .A4(MSB), .ZN(
        net34754) );
  AND2_X1 U93 ( .A1(MASK16[25]), .A2(n2), .ZN(n131) );
  AND2_X1 U94 ( .A1(MASK8[25]), .A2(net27138), .ZN(n132) );
  NOR3_X1 U95 ( .A1(n131), .A2(n132), .A3(n102), .ZN(n55) );
  BUF_X2 U96 ( .A(net27156), .Z(net27148) );
  AND2_X1 U97 ( .A1(MASK16[4]), .A2(net27152), .ZN(n133) );
  AND2_X1 U98 ( .A1(MASK8[4]), .A2(net27142), .ZN(n134) );
  NOR3_X1 U99 ( .A1(n134), .A2(n133), .A3(net34755), .ZN(n19) );
  AND2_X1 U100 ( .A1(MASK16[3]), .A2(net40402), .ZN(n135) );
  AND2_X1 U101 ( .A1(MASK8[3]), .A2(n43), .ZN(n136) );
  NOR3_X1 U102 ( .A1(n135), .A2(n136), .A3(net34755), .ZN(n23) );
  AND2_X1 U103 ( .A1(MASK16[23]), .A2(net40443), .ZN(n137) );
  AND2_X1 U104 ( .A1(MASK8[23]), .A2(net35591), .ZN(n138) );
  BUF_X1 U105 ( .A(net27144), .Z(net35590) );
  AND2_X1 U106 ( .A1(MASK16[22]), .A2(net27150), .ZN(n139) );
  AND2_X1 U107 ( .A1(MASK8[22]), .A2(net27136), .ZN(n140) );
  NOR3_X1 U108 ( .A1(n139), .A2(n140), .A3(n100), .ZN(n61) );
  AND2_X1 U109 ( .A1(MASK16[28]), .A2(net40443), .ZN(n141) );
  AND2_X1 U110 ( .A1(MASK8[28]), .A2(net35590), .ZN(n142) );
  NOR3_X1 U111 ( .A1(n141), .A2(n142), .A3(n94), .ZN(n49) );
  AND2_X1 U112 ( .A1(MASK16[27]), .A2(net40444), .ZN(n143) );
  AND2_X1 U113 ( .A1(MASK8[27]), .A2(net35591), .ZN(n144) );
  NOR3_X1 U114 ( .A1(n143), .A2(n144), .A3(net34755), .ZN(n51) );
  AND2_X1 U115 ( .A1(MASK8[30]), .A2(net35590), .ZN(n145) );
  AND2_X1 U116 ( .A1(MASK16[29]), .A2(net40443), .ZN(n146) );
  AND2_X1 U117 ( .A1(MASK8[29]), .A2(net27136), .ZN(n147) );
  NOR3_X1 U118 ( .A1(n146), .A2(net34755), .A3(n147), .ZN(n47) );
  AND2_X1 U119 ( .A1(MASK16[12]), .A2(net27150), .ZN(n148) );
  AND2_X1 U120 ( .A1(MASK8[12]), .A2(net27136), .ZN(n149) );
  NOR3_X1 U121 ( .A1(n148), .A2(n149), .A3(net34755), .ZN(n83) );
  AND2_X1 U122 ( .A1(MASK16[34]), .A2(net27154), .ZN(n150) );
  AND2_X1 U123 ( .A1(MASK8[34]), .A2(n43), .ZN(n151) );
  NOR3_X1 U124 ( .A1(n150), .A2(n151), .A3(net34754), .ZN(n35) );
  AND2_X1 U125 ( .A1(MASK16[17]), .A2(n2), .ZN(n152) );
  AND2_X1 U126 ( .A1(MASK8[17]), .A2(net35591), .ZN(n153) );
  NOR3_X1 U127 ( .A1(n152), .A2(n153), .A3(n94), .ZN(n73) );
  AND2_X1 U128 ( .A1(MASK16[21]), .A2(net40444), .ZN(n154) );
  AND2_X1 U129 ( .A1(MASK8[21]), .A2(n43), .ZN(n155) );
  NOR3_X1 U130 ( .A1(n154), .A2(n155), .A3(n94), .ZN(n63) );
  AND2_X1 U131 ( .A1(MASK16[20]), .A2(net27150), .ZN(n156) );
  AND2_X1 U132 ( .A1(MASK8[20]), .A2(n1), .ZN(n157) );
  NOR3_X1 U133 ( .A1(n156), .A2(n157), .A3(n102), .ZN(n65) );
  AND2_X1 U134 ( .A1(MASK16[19]), .A2(net27150), .ZN(n158) );
  AND2_X1 U135 ( .A1(MASK8[19]), .A2(n43), .ZN(n159) );
  NOR3_X1 U136 ( .A1(n158), .A2(n159), .A3(net34755), .ZN(n69) );
  AND2_X1 U137 ( .A1(MASK16[24]), .A2(net27148), .ZN(n160) );
  AND2_X1 U138 ( .A1(MASK8[24]), .A2(net27136), .ZN(n161) );
  NOR3_X1 U139 ( .A1(n160), .A2(n161), .A3(net34754), .ZN(n57) );
  AND2_X1 U140 ( .A1(MASK16[26]), .A2(net40443), .ZN(n162) );
  AND2_X1 U141 ( .A1(MASK8[26]), .A2(net35591), .ZN(n163) );
  NOR3_X1 U142 ( .A1(n162), .A2(n163), .A3(n100), .ZN(n53) );
  AND2_X1 U143 ( .A1(MASK16[16]), .A2(net27148), .ZN(n164) );
  AND2_X1 U144 ( .A1(MASK8[16]), .A2(n43), .ZN(n165) );
  NOR3_X1 U145 ( .A1(n164), .A2(n165), .A3(net34754), .ZN(n75) );
  AND2_X1 U146 ( .A1(MASK16[15]), .A2(net40444), .ZN(n166) );
  AND2_X1 U147 ( .A1(MASK8[15]), .A2(net27136), .ZN(n167) );
  NOR3_X1 U148 ( .A1(n166), .A2(n167), .A3(net34755), .ZN(n77) );
  AND2_X1 U149 ( .A1(MASK16[10]), .A2(n2), .ZN(n168) );
  AND2_X1 U150 ( .A1(MASK8[10]), .A2(net27138), .ZN(n169) );
  NOR3_X1 U151 ( .A1(n168), .A2(n169), .A3(net34755), .ZN(n87) );
  AND2_X1 U152 ( .A1(MASK16[14]), .A2(net27152), .ZN(n170) );
  AND2_X1 U153 ( .A1(MASK8[14]), .A2(net27140), .ZN(n171) );
  NOR3_X1 U154 ( .A1(n170), .A2(n171), .A3(net34755), .ZN(n79) );
  AND2_X1 U155 ( .A1(MASK16[11]), .A2(net27148), .ZN(n172) );
  AND2_X1 U156 ( .A1(MASK8[11]), .A2(net35590), .ZN(n173) );
  NOR3_X1 U157 ( .A1(n172), .A2(n173), .A3(net34755), .ZN(n85) );
  AND2_X1 U158 ( .A1(MASK16[9]), .A2(net27152), .ZN(n174) );
  AND2_X1 U159 ( .A1(MASK8[9]), .A2(net27138), .ZN(n175) );
  NOR3_X1 U160 ( .A1(n174), .A2(n175), .A3(n100), .ZN(n6) );
  AND2_X1 U161 ( .A1(MASK16[32]), .A2(net27152), .ZN(n176) );
  AND2_X1 U162 ( .A1(MASK8[32]), .A2(net27140), .ZN(n177) );
  NOR3_X1 U163 ( .A1(n176), .A2(n94), .A3(n177), .ZN(n39) );
  AND2_X1 U164 ( .A1(net27154), .A2(MASK16[35]), .ZN(n178) );
  AND2_X1 U165 ( .A1(MASK8[35]), .A2(net27138), .ZN(n179) );
  NOR3_X1 U166 ( .A1(n179), .A2(n178), .A3(net34755), .ZN(n33) );
  AND2_X1 U167 ( .A1(MASK16[31]), .A2(net27154), .ZN(n180) );
  AND2_X1 U168 ( .A1(MASK8[31]), .A2(net27140), .ZN(n181) );
  NOR3_X1 U169 ( .A1(n180), .A2(n181), .A3(net34755), .ZN(n41) );
  AND2_X1 U170 ( .A1(MASK16[13]), .A2(net27148), .ZN(n182) );
  AND2_X1 U171 ( .A1(MASK8[13]), .A2(net35590), .ZN(n183) );
  NOR3_X1 U172 ( .A1(n182), .A2(n183), .A3(n94), .ZN(n81) );
  AND2_X1 U173 ( .A1(MASK16[33]), .A2(net27154), .ZN(n184) );
  AND2_X1 U174 ( .A1(MASK8[33]), .A2(net27140), .ZN(n185) );
  NOR3_X1 U175 ( .A1(n100), .A2(n185), .A3(n184), .ZN(n37) );
  CLKBUF_X1 U176 ( .A(n7), .Z(net27110) );
  CLKBUF_X1 U177 ( .A(net27110), .Z(net27102) );
  AND2_X1 U178 ( .A1(MASK16[18]), .A2(net27150), .ZN(n186) );
  AND2_X1 U179 ( .A1(MASK8[18]), .A2(net35590), .ZN(n187) );
  NOR3_X1 U180 ( .A1(n186), .A2(n187), .A3(net34755), .ZN(n71) );
  AND2_X1 U181 ( .A1(MASK16[7]), .A2(net27154), .ZN(n188) );
  AND2_X1 U182 ( .A1(MASK8[7]), .A2(n43), .ZN(n189) );
  NOR3_X1 U183 ( .A1(n189), .A2(net34755), .A3(n188), .ZN(n13) );
  NAND2_X1 U184 ( .A1(n20), .A2(n21), .ZN(S[40]) );
  AOI22_X1 U185 ( .A1(MASK24[40]), .A2(net27112), .B1(MASK0[40]), .B2(net27124), .ZN(n20) );
  NAND2_X1 U186 ( .A1(n49), .A2(n48), .ZN(S[28]) );
  AOI22_X1 U187 ( .A1(MASK24[28]), .A2(net27114), .B1(MASK0[28]), .B2(net27126), .ZN(n48) );
  NAND2_X1 U188 ( .A1(n51), .A2(n50), .ZN(S[27]) );
  AOI22_X1 U189 ( .A1(MASK24[27]), .A2(net27114), .B1(MASK0[27]), .B2(net27126), .ZN(n50) );
  NAND2_X1 U190 ( .A1(n41), .A2(n40), .ZN(S[31]) );
  AOI22_X1 U191 ( .A1(MASK24[31]), .A2(net27114), .B1(MASK0[31]), .B2(net27128), .ZN(n40) );
  AOI22_X1 U192 ( .A1(MASK24[30]), .A2(net27114), .B1(MASK0[30]), .B2(net27128), .ZN(n42) );
  NAND2_X1 U193 ( .A1(n47), .A2(n46), .ZN(S[29]) );
  AOI22_X1 U194 ( .A1(MASK24[29]), .A2(net27114), .B1(MASK0[29]), .B2(net27128), .ZN(n46) );
  NAND2_X1 U195 ( .A1(n53), .A2(n52), .ZN(S[26]) );
  AOI22_X1 U196 ( .A1(MASK24[26]), .A2(net27114), .B1(MASK0[26]), .B2(n109), 
        .ZN(n52) );
  NAND2_X1 U197 ( .A1(n55), .A2(n54), .ZN(S[25]) );
  AOI22_X1 U198 ( .A1(MASK24[25]), .A2(net27116), .B1(MASK0[25]), .B2(n109), 
        .ZN(n54) );
  NAND2_X1 U199 ( .A1(n39), .A2(n38), .ZN(S[32]) );
  AOI22_X1 U200 ( .A1(MASK24[32]), .A2(net27114), .B1(MASK0[32]), .B2(net27126), .ZN(n38) );
  NAND2_X1 U201 ( .A1(n35), .A2(n34), .ZN(S[34]) );
  AOI22_X1 U202 ( .A1(MASK24[34]), .A2(net27114), .B1(MASK0[34]), .B2(net27128), .ZN(n34) );
  NAND2_X1 U203 ( .A1(n37), .A2(n36), .ZN(S[33]) );
  AOI22_X1 U204 ( .A1(MASK24[33]), .A2(net27114), .B1(MASK0[33]), .B2(net27128), .ZN(n36) );
  NAND2_X1 U205 ( .A1(n57), .A2(n56), .ZN(S[24]) );
  AOI22_X1 U206 ( .A1(MASK24[24]), .A2(net27116), .B1(MASK0[24]), .B2(n109), 
        .ZN(n56) );
  NAND2_X1 U207 ( .A1(n59), .A2(n58), .ZN(S[23]) );
  AOI22_X1 U208 ( .A1(MASK24[23]), .A2(net27116), .B1(MASK0[23]), .B2(net27126), .ZN(n58) );
  NAND2_X1 U209 ( .A1(n61), .A2(n60), .ZN(S[22]) );
  AOI22_X1 U210 ( .A1(MASK24[22]), .A2(net27116), .B1(MASK0[22]), .B2(net27124), .ZN(n60) );
  NAND2_X1 U211 ( .A1(n63), .A2(n62), .ZN(S[21]) );
  AOI22_X1 U212 ( .A1(MASK24[21]), .A2(net27116), .B1(MASK0[21]), .B2(n109), 
        .ZN(n62) );
  NAND2_X1 U213 ( .A1(n69), .A2(n68), .ZN(S[19]) );
  AOI22_X1 U214 ( .A1(MASK24[19]), .A2(net27116), .B1(MASK0[19]), .B2(net27124), .ZN(n68) );
  NAND2_X1 U215 ( .A1(n65), .A2(n64), .ZN(S[20]) );
  AOI22_X1 U216 ( .A1(MASK24[20]), .A2(net27116), .B1(MASK0[20]), .B2(net27126), .ZN(n64) );
  NAND2_X1 U217 ( .A1(n78), .A2(n79), .ZN(S[14]) );
  AOI22_X1 U218 ( .A1(MASK24[14]), .A2(net27116), .B1(MASK0[14]), .B2(net27126), .ZN(n78) );
  NAND2_X1 U219 ( .A1(n77), .A2(n76), .ZN(S[15]) );
  AOI22_X1 U220 ( .A1(MASK24[15]), .A2(net27116), .B1(MASK0[15]), .B2(n109), 
        .ZN(n76) );
  NAND2_X1 U221 ( .A1(n74), .A2(n75), .ZN(S[16]) );
  AOI22_X1 U222 ( .A1(MASK24[16]), .A2(net27116), .B1(MASK0[16]), .B2(n109), 
        .ZN(n74) );
  NAND2_X1 U223 ( .A1(n73), .A2(n72), .ZN(S[17]) );
  AOI22_X1 U224 ( .A1(MASK24[17]), .A2(net27116), .B1(MASK0[17]), .B2(net27126), .ZN(n72) );
  NAND2_X1 U225 ( .A1(n71), .A2(n70), .ZN(S[18]) );
  AOI22_X1 U226 ( .A1(MASK24[18]), .A2(net27116), .B1(MASK0[18]), .B2(net27126), .ZN(n70) );
  NAND2_X1 U227 ( .A1(n29), .A2(n28), .ZN(S[37]) );
  AOI22_X1 U228 ( .A1(MASK24[37]), .A2(net27112), .B1(MASK0[37]), .B2(net27128), .ZN(n28) );
  NAND2_X1 U229 ( .A1(n22), .A2(n23), .ZN(S[3]) );
  AOI22_X1 U230 ( .A1(MASK24[3]), .A2(net27112), .B1(MASK0[3]), .B2(net27126), 
        .ZN(n22) );
  NAND2_X1 U231 ( .A1(n19), .A2(n18), .ZN(S[4]) );
  AOI22_X1 U232 ( .A1(MASK24[4]), .A2(net27112), .B1(MASK0[4]), .B2(n109), 
        .ZN(n18) );
  NAND2_X1 U233 ( .A1(n30), .A2(n31), .ZN(S[36]) );
  AOI22_X1 U234 ( .A1(MASK24[36]), .A2(net27112), .B1(MASK0[36]), .B2(net27128), .ZN(n30) );
  NAND2_X1 U235 ( .A1(n5), .A2(n6), .ZN(S[9]) );
  AOI22_X1 U236 ( .A1(MASK24[9]), .A2(net27114), .B1(MASK0[9]), .B2(net27124), 
        .ZN(n5) );
  NAND2_X1 U237 ( .A1(n87), .A2(n86), .ZN(S[10]) );
  AOI22_X1 U238 ( .A1(MASK24[10]), .A2(net27116), .B1(MASK0[10]), .B2(n109), 
        .ZN(n86) );
  NAND2_X1 U239 ( .A1(n85), .A2(n84), .ZN(S[11]) );
  AOI22_X1 U240 ( .A1(MASK24[11]), .A2(net27116), .B1(MASK0[11]), .B2(net27126), .ZN(n84) );
  NAND2_X1 U241 ( .A1(n83), .A2(n82), .ZN(S[12]) );
  AOI22_X1 U242 ( .A1(MASK24[12]), .A2(net27116), .B1(MASK0[12]), .B2(net27128), .ZN(n82) );
  NAND2_X1 U243 ( .A1(n81), .A2(n80), .ZN(S[13]) );
  AOI22_X1 U244 ( .A1(MASK24[13]), .A2(net27116), .B1(MASK0[13]), .B2(net27124), .ZN(n80) );
  NAND2_X1 U245 ( .A1(n26), .A2(n27), .ZN(S[38]) );
  AOI22_X1 U246 ( .A1(MASK24[38]), .A2(net27112), .B1(MASK0[38]), .B2(n109), 
        .ZN(n26) );
  AOI221_X1 U247 ( .B1(MASK16[38]), .B2(net40402), .C1(MASK8[38]), .C2(
        net27142), .A(n7), .ZN(n27) );
  AOI221_X1 U248 ( .B1(MASK16[37]), .B2(net40402), .C1(MASK8[37]), .C2(
        net27142), .A(n7), .ZN(n29) );
  AOI221_X1 U249 ( .B1(net40402), .B2(MASK16[36]), .C1(MASK8[36]), .C2(
        net27142), .A(n7), .ZN(n31) );
  NAND2_X1 U250 ( .A1(n24), .A2(n25), .ZN(S[39]) );
  AOI22_X1 U251 ( .A1(MASK24[39]), .A2(net27112), .B1(MASK0[39]), .B2(n109), 
        .ZN(n24) );
  NAND2_X1 U252 ( .A1(n33), .A2(n32), .ZN(S[35]) );
  AOI22_X1 U253 ( .A1(MASK24[35]), .A2(net27114), .B1(MASK0[35]), .B2(net27124), .ZN(n32) );
  NAND2_X1 U254 ( .A1(n14), .A2(n15), .ZN(S[6]) );
  AOI22_X1 U255 ( .A1(MASK24[6]), .A2(net27112), .B1(MASK0[6]), .B2(net27126), 
        .ZN(n14) );
  AOI221_X1 U256 ( .B1(MASK16[6]), .B2(net27148), .C1(MASK8[6]), .C2(net27142), 
        .A(n102), .ZN(n15) );
  NAND2_X1 U257 ( .A1(n13), .A2(n12), .ZN(S[7]) );
  AOI22_X1 U258 ( .A1(MASK24[7]), .A2(net27112), .B1(MASK0[7]), .B2(net27128), 
        .ZN(n12) );
  NAND2_X1 U259 ( .A1(n66), .A2(n67), .ZN(S[1]) );
  AOI22_X1 U260 ( .A1(MASK24[1]), .A2(net27116), .B1(MASK0[1]), .B2(net27126), 
        .ZN(n66) );
  AOI221_X1 U261 ( .B1(MASK16[1]), .B2(net40444), .C1(MASK8[1]), .C2(net27142), 
        .A(net27110), .ZN(n67) );
  NAND2_X1 U262 ( .A1(n16), .A2(n17), .ZN(S[5]) );
  AOI22_X1 U263 ( .A1(MASK24[5]), .A2(net27112), .B1(MASK0[5]), .B2(net27126), 
        .ZN(n16) );
  AOI221_X1 U264 ( .B1(MASK16[5]), .B2(net40402), .C1(MASK8[5]), .C2(net27142), 
        .A(n102), .ZN(n17) );
  NAND2_X1 U265 ( .A1(n44), .A2(n45), .ZN(S[2]) );
  AOI22_X1 U266 ( .A1(MASK24[2]), .A2(net27114), .B1(MASK0[2]), .B2(n109), 
        .ZN(n44) );
  AOI221_X1 U267 ( .B1(MASK16[2]), .B2(net40402), .C1(MASK8[2]), .C2(net27142), 
        .A(n100), .ZN(n45) );
  NAND2_X1 U268 ( .A1(n88), .A2(n89), .ZN(S[0]) );
  AOI22_X1 U269 ( .A1(MASK24[0]), .A2(net27112), .B1(MASK0[0]), .B2(net27124), 
        .ZN(n88) );
endmodule


module FINE_SHIFT_DATA_W32_MASK_SIZE41_1 ( A, AMOUNT, S );
  input [40:0] A;
  input [2:0] AMOUNT;
  output [31:0] S;
  wire   \U1/net27040 , \U1/net27042 , \U1/net27044 , \U1/net27034 ,
         \U1/net27036 , \U1/net27038 , \U1/net27030 , \U1/net27022 ,
         \U1/net27024 , \U1/net27026 , \U1/net27028 , \U1/net24085 ,
         \U1/net24083 , \U1/net24076 , \U1/net24052 , \U1/net24040 ,
         \U1/net24039 , \U1/net24038 , \U1/net24034 , \U1/net24029 ,
         \U1/net5922 , \U1/net5920 , \U1/net5919 , \U1/net5917 , \U1/net5916 ,
         \U1/net5908 , \U1/net5905 , \U1/net5901 , \U1/net5898 , \U1/net5897 ,
         net34789, net34856, net34866, net34865, net40398, net40397,
         \U1/net5910 , \U1/net5904 , \U1/net5911 , \U1/net24082 , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141;

  BUF_X1 U1 ( .A(AMOUNT[1]), .Z(\U1/net27036 ) );
  BUF_X1 U2 ( .A(AMOUNT[1]), .Z(\U1/net27038 ) );
  BUF_X2 U3 ( .A(AMOUNT[1]), .Z(\U1/net27034 ) );
  BUF_X2 U4 ( .A(n16), .Z(\U1/net27026 ) );
  BUF_X1 U5 ( .A(AMOUNT[0]), .Z(\U1/net27040 ) );
  AND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(n1) );
  MUX2_X1 U7 ( .A(n75), .B(n71), .S(\U1/net27034 ), .Z(n2) );
  MUX2_X1 U8 ( .A(n75), .B(n71), .S(\U1/net27034 ), .Z(n76) );
  INV_X1 U9 ( .A(A[25]), .ZN(n3) );
  MUX2_X2 U10 ( .A(n116), .B(\U1/net24038 ), .S(\U1/net27024 ), .Z(n54) );
  MUX2_X1 U11 ( .A(n103), .B(n108), .S(\U1/net27024 ), .Z(n83) );
  MUX2_X2 U12 ( .A(n77), .B(n73), .S(\U1/net27034 ), .Z(n78) );
  NAND2_X1 U13 ( .A1(n58), .A2(n4), .ZN(n5) );
  NAND2_X1 U14 ( .A1(n54), .A2(\U1/net27036 ), .ZN(n6) );
  INV_X1 U15 ( .A(\U1/net27036 ), .ZN(n4) );
  MUX2_X1 U16 ( .A(n109), .B(n102), .S(net34865), .Z(n7) );
  NAND2_X1 U17 ( .A1(n12), .A2(\U1/net27028 ), .ZN(n8) );
  NAND2_X1 U18 ( .A1(n14), .A2(net34865), .ZN(n9) );
  NAND2_X1 U19 ( .A1(n8), .A2(n9), .ZN(n18) );
  MUX2_X1 U20 ( .A(n15), .B(\U1/net24083 ), .S(n22), .Z(S[6]) );
  MUX2_X1 U21 ( .A(n129), .B(n112), .S(n22), .Z(S[29]) );
  MUX2_X1 U22 ( .A(n103), .B(n99), .S(net40397), .Z(n44) );
  MUX2_X1 U23 ( .A(n109), .B(n102), .S(net34865), .Z(n85) );
  MUX2_X1 U24 ( .A(n135), .B(n113), .S(n22), .Z(S[23]) );
  MUX2_X1 U25 ( .A(n133), .B(n107), .S(net40397), .Z(n73) );
  MUX2_X1 U26 ( .A(n14), .B(\U1/net24052 ), .S(net34865), .Z(net34789) );
  OR2_X1 U27 ( .A1(n93), .A2(n22), .ZN(n43) );
  MUX2_X1 U28 ( .A(\U1/net24052 ), .B(n120), .S(net40397), .Z(n59) );
  MUX2_X1 U29 ( .A(n102), .B(n98), .S(net40397), .Z(n92) );
  BUF_X2 U30 ( .A(\U1/net27030 ), .Z(\U1/net27022 ) );
  MUX2_X1 U31 ( .A(A[12]), .B(A[8]), .S(AMOUNT[2]), .Z(n10) );
  INV_X1 U32 ( .A(n10), .ZN(\U1/net5910 ) );
  MUX2_X1 U33 ( .A(\U1/net24082 ), .B(n15), .S(n22), .Z(S[5]) );
  INV_X1 U34 ( .A(\U1/net27040 ), .ZN(n22) );
  INV_X1 U35 ( .A(n19), .ZN(n15) );
  MUX2_X1 U36 ( .A(n18), .B(n17), .S(\U1/net27038 ), .Z(n19) );
  INV_X1 U37 ( .A(\U1/net5911 ), .ZN(\U1/net24082 ) );
  MUX2_X1 U38 ( .A(\U1/net24082 ), .B(\U1/net24034 ), .S(\U1/net27044 ), .Z(
        S[4]) );
  MUX2_X1 U39 ( .A(\U1/net5910 ), .B(\U1/net5904 ), .S(\U1/net27038 ), .Z(
        \U1/net5911 ) );
  BUF_X1 U40 ( .A(AMOUNT[0]), .Z(\U1/net27042 ) );
  BUF_X1 U41 ( .A(AMOUNT[0]), .Z(\U1/net27044 ) );
  MUX2_X1 U42 ( .A(\U1/net5919 ), .B(n18), .S(\U1/net27038 ), .Z(\U1/net5920 )
         );
  BUF_X1 U43 ( .A(AMOUNT[2]), .Z(n16) );
  BUF_X1 U44 ( .A(n16), .Z(\U1/net27028 ) );
  INV_X1 U45 ( .A(A[9]), .ZN(n12) );
  NAND2_X1 U46 ( .A1(n12), .A2(net40397), .ZN(net40398) );
  INV_X1 U47 ( .A(A[13]), .ZN(n14) );
  NAND2_X1 U48 ( .A1(n21), .A2(n20), .ZN(n17) );
  MUX2_X1 U49 ( .A(n17), .B(\U1/net5901 ), .S(\U1/net27038 ), .Z(\U1/net5908 )
         );
  NAND2_X1 U50 ( .A1(n13), .A2(net34865), .ZN(n20) );
  INV_X1 U51 ( .A(A[11]), .ZN(n13) );
  MUX2_X1 U52 ( .A(\U1/net24039 ), .B(n13), .S(\U1/net27026 ), .Z(\U1/net5919 ) );
  NAND2_X1 U53 ( .A1(n11), .A2(\U1/net27026 ), .ZN(n21) );
  INV_X1 U54 ( .A(A[7]), .ZN(n11) );
  NAND2_X1 U55 ( .A1(n11), .A2(net34865), .ZN(net34856) );
  INV_X1 U56 ( .A(A[12]), .ZN(n25) );
  MUX2_X1 U57 ( .A(\U1/net24076 ), .B(n25), .S(\U1/net27026 ), .Z(\U1/net5922 ) );
  INV_X1 U58 ( .A(A[8]), .ZN(n26) );
  NAND2_X1 U59 ( .A1(n26), .A2(net34865), .ZN(net34866) );
  MUX2_X1 U60 ( .A(n24), .B(n23), .S(\U1/net27026 ), .Z(\U1/net5904 ) );
  MUX2_X1 U61 ( .A(\U1/net5904 ), .B(\U1/net5898 ), .S(\U1/net27038 ), .Z(
        \U1/net5905 ) );
  INV_X1 U62 ( .A(A[6]), .ZN(n23) );
  MUX2_X1 U63 ( .A(n23), .B(\U1/net24029 ), .S(\U1/net27026 ), .Z(\U1/net5897 ) );
  INV_X1 U64 ( .A(A[10]), .ZN(n24) );
  MUX2_X1 U65 ( .A(\U1/net24038 ), .B(n24), .S(\U1/net27026 ), .Z(\U1/net5916 ) );
  BUF_X1 U66 ( .A(AMOUNT[2]), .Z(\U1/net27030 ) );
  OR2_X1 U67 ( .A1(A[23]), .A2(\U1/net27024 ), .ZN(n37) );
  OR2_X1 U68 ( .A1(n78), .A2(\U1/net27040 ), .ZN(n30) );
  OR2_X1 U69 ( .A1(n76), .A2(n22), .ZN(n31) );
  NAND2_X1 U70 ( .A1(n106), .A2(net40397), .ZN(n27) );
  NAND2_X1 U71 ( .A1(n123), .A2(\U1/net27024 ), .ZN(n28) );
  NAND2_X1 U72 ( .A1(n27), .A2(n28), .ZN(n71) );
  BUF_X2 U73 ( .A(\U1/net27030 ), .Z(\U1/net27024 ) );
  NAND2_X1 U74 ( .A1(n94), .A2(\U1/net27026 ), .ZN(n29) );
  NAND2_X1 U75 ( .A1(net40398), .A2(n29), .ZN(\U1/net5901 ) );
  INV_X1 U76 ( .A(\U1/net27026 ), .ZN(net40397) );
  NAND2_X1 U77 ( .A1(n30), .A2(n31), .ZN(S[22]) );
  MUX2_X1 U78 ( .A(n108), .B(n3), .S(\U1/net27022 ), .Z(n32) );
  MUX2_X1 U79 ( .A(n100), .B(n128), .S(\U1/net27022 ), .Z(n33) );
  NAND2_X1 U80 ( .A1(n95), .A2(\U1/net27026 ), .ZN(n34) );
  NAND2_X1 U81 ( .A1(n34), .A2(net34866), .ZN(\U1/net5898 ) );
  INV_X1 U82 ( .A(\U1/net27026 ), .ZN(net34865) );
  NAND2_X1 U83 ( .A1(n96), .A2(\U1/net27026 ), .ZN(n35) );
  NAND2_X1 U84 ( .A1(net34856), .A2(n35), .ZN(n49) );
  MUX2_X1 U85 ( .A(n122), .B(n116), .S(\U1/net27024 ), .Z(n36) );
  NAND2_X1 U86 ( .A1(n117), .A2(\U1/net27024 ), .ZN(n38) );
  NAND2_X1 U87 ( .A1(n38), .A2(n37), .ZN(n63) );
  NAND2_X1 U88 ( .A1(n3), .A2(net40397), .ZN(n39) );
  NAND2_X1 U89 ( .A1(n120), .A2(\U1/net27024 ), .ZN(n40) );
  NAND2_X1 U90 ( .A1(n39), .A2(n40), .ZN(n67) );
  MUX2_X1 U91 ( .A(n126), .B(n136), .S(n22), .Z(S[16]) );
  MUX2_X1 U92 ( .A(A[37]), .B(A[33]), .S(\U1/net27022 ), .Z(n41) );
  NAND2_X1 U93 ( .A1(n48), .A2(n22), .ZN(n42) );
  NAND2_X1 U94 ( .A1(n43), .A2(n42), .ZN(S[31]) );
  INV_X1 U95 ( .A(n49), .ZN(n97) );
  INV_X1 U96 ( .A(A[28]), .ZN(n107) );
  INV_X1 U97 ( .A(A[27]), .ZN(n106) );
  INV_X1 U98 ( .A(A[31]), .ZN(n110) );
  INV_X1 U99 ( .A(A[30]), .ZN(n109) );
  INV_X1 U100 ( .A(A[29]), .ZN(n108) );
  INV_X1 U101 ( .A(A[26]), .ZN(n105) );
  INV_X1 U102 ( .A(A[32]), .ZN(n128) );
  INV_X1 U103 ( .A(A[34]), .ZN(n102) );
  INV_X1 U104 ( .A(A[33]), .ZN(n103) );
  INV_X1 U105 ( .A(A[24]), .ZN(n133) );
  INV_X1 U106 ( .A(A[23]), .ZN(n123) );
  INV_X1 U107 ( .A(A[22]), .ZN(n122) );
  INV_X1 U108 ( .A(A[21]), .ZN(n120) );
  INV_X1 U109 ( .A(A[19]), .ZN(n117) );
  INV_X1 U110 ( .A(A[20]), .ZN(n119) );
  INV_X1 U111 ( .A(A[14]), .ZN(\U1/net24038 ) );
  INV_X1 U112 ( .A(A[15]), .ZN(\U1/net24039 ) );
  INV_X1 U113 ( .A(A[16]), .ZN(\U1/net24076 ) );
  INV_X1 U114 ( .A(A[17]), .ZN(\U1/net24052 ) );
  INV_X1 U115 ( .A(A[18]), .ZN(n116) );
  INV_X1 U116 ( .A(A[37]), .ZN(n99) );
  INV_X1 U117 ( .A(A[3]), .ZN(n96) );
  INV_X1 U118 ( .A(n91), .ZN(n112) );
  INV_X1 U119 ( .A(n86), .ZN(n132) );
  INV_X1 U120 ( .A(n2), .ZN(n125) );
  INV_X1 U121 ( .A(n74), .ZN(n134) );
  INV_X1 U122 ( .A(n78), .ZN(n135) );
  INV_X1 U123 ( .A(n80), .ZN(n113) );
  INV_X1 U124 ( .A(n82), .ZN(n131) );
  INV_X1 U125 ( .A(n84), .ZN(n114) );
  INV_X1 U126 ( .A(n90), .ZN(n129) );
  INV_X1 U127 ( .A(n93), .ZN(n130) );
  INV_X1 U128 ( .A(A[38]), .ZN(n98) );
  INV_X1 U129 ( .A(n88), .ZN(n111) );
  INV_X1 U130 ( .A(n72), .ZN(n124) );
  INV_X1 U131 ( .A(n51), .ZN(n104) );
  INV_X1 U132 ( .A(n68), .ZN(n127) );
  INV_X1 U133 ( .A(n70), .ZN(n137) );
  INV_X1 U134 ( .A(\U1/net5908 ), .ZN(\U1/net24034 ) );
  INV_X1 U135 ( .A(\U1/net5905 ), .ZN(\U1/net24085 ) );
  INV_X1 U136 ( .A(\U1/net5917 ), .ZN(\U1/net24083 ) );
  INV_X1 U137 ( .A(\U1/net5920 ), .ZN(\U1/net24040 ) );
  INV_X1 U138 ( .A(n57), .ZN(n118) );
  INV_X1 U139 ( .A(n60), .ZN(n121) );
  INV_X1 U140 ( .A(n62), .ZN(n138) );
  INV_X1 U141 ( .A(n64), .ZN(n126) );
  INV_X1 U142 ( .A(n66), .ZN(n136) );
  INV_X1 U143 ( .A(n52), .ZN(n139) );
  INV_X1 U144 ( .A(n53), .ZN(n115) );
  INV_X1 U145 ( .A(n55), .ZN(n140) );
  INV_X1 U146 ( .A(A[35]), .ZN(n101) );
  INV_X1 U147 ( .A(A[4]), .ZN(n95) );
  INV_X1 U148 ( .A(A[36]), .ZN(n100) );
  INV_X1 U149 ( .A(n50), .ZN(n141) );
  INV_X1 U150 ( .A(A[2]), .ZN(\U1/net24029 ) );
  INV_X1 U151 ( .A(A[5]), .ZN(n94) );
  MUX2_X1 U152 ( .A(A[5]), .B(A[1]), .S(\U1/net27028 ), .Z(n45) );
  MUX2_X1 U153 ( .A(n97), .B(n45), .S(\U1/net27038 ), .Z(n46) );
  MUX2_X1 U154 ( .A(n141), .B(n46), .S(\U1/net27044 ), .Z(S[0]) );
  MUX2_X1 U155 ( .A(n104), .B(n141), .S(\U1/net27044 ), .Z(S[1]) );
  MUX2_X1 U156 ( .A(\U1/net24085 ), .B(n104), .S(\U1/net27044 ), .Z(S[2]) );
  MUX2_X1 U157 ( .A(\U1/net24034 ), .B(\U1/net24085 ), .S(\U1/net27044 ), .Z(
        S[3]) );
  MUX2_X1 U158 ( .A(\U1/net24040 ), .B(\U1/net24083 ), .S(\U1/net27044 ), .Z(
        S[7]) );
  MUX2_X1 U159 ( .A(n139), .B(\U1/net24040 ), .S(\U1/net27044 ), .Z(S[8]) );
  MUX2_X1 U160 ( .A(n115), .B(n139), .S(\U1/net27044 ), .Z(S[9]) );
  MUX2_X1 U161 ( .A(n140), .B(n115), .S(\U1/net27042 ), .Z(S[10]) );
  MUX2_X1 U162 ( .A(n118), .B(n140), .S(\U1/net27042 ), .Z(S[11]) );
  MUX2_X1 U163 ( .A(n1), .B(n118), .S(\U1/net27042 ), .Z(S[12]) );
  MUX2_X1 U164 ( .A(n121), .B(n1), .S(\U1/net27042 ), .Z(S[13]) );
  MUX2_X1 U165 ( .A(n138), .B(n121), .S(\U1/net27042 ), .Z(S[14]) );
  MUX2_X1 U166 ( .A(n126), .B(n138), .S(\U1/net27042 ), .Z(S[15]) );
  MUX2_X1 U167 ( .A(n127), .B(n136), .S(\U1/net27042 ), .Z(S[17]) );
  MUX2_X1 U168 ( .A(n137), .B(n127), .S(\U1/net27042 ), .Z(S[18]) );
  MUX2_X1 U169 ( .A(n124), .B(n137), .S(\U1/net27042 ), .Z(S[19]) );
  MUX2_X1 U170 ( .A(n134), .B(n124), .S(\U1/net27042 ), .Z(S[20]) );
  MUX2_X1 U171 ( .A(n125), .B(n134), .S(\U1/net27040 ), .Z(S[21]) );
  MUX2_X1 U172 ( .A(n131), .B(n113), .S(\U1/net27040 ), .Z(S[24]) );
  MUX2_X1 U173 ( .A(n114), .B(n131), .S(\U1/net27040 ), .Z(S[25]) );
  MUX2_X1 U174 ( .A(n132), .B(n114), .S(\U1/net27040 ), .Z(S[26]) );
  MUX2_X1 U175 ( .A(n111), .B(n132), .S(\U1/net27040 ), .Z(S[27]) );
  MUX2_X1 U176 ( .A(n129), .B(n111), .S(\U1/net27040 ), .Z(S[28]) );
  MUX2_X1 U177 ( .A(n130), .B(n112), .S(\U1/net27040 ), .Z(S[30]) );
  MUX2_X1 U178 ( .A(A[39]), .B(A[35]), .S(\U1/net27028 ), .Z(n47) );
  MUX2_X1 U179 ( .A(n47), .B(n41), .S(\U1/net27038 ), .Z(n48) );
  MUX2_X1 U180 ( .A(\U1/net5898 ), .B(\U1/net5897 ), .S(\U1/net27038 ), .Z(n50) );
  MUX2_X1 U181 ( .A(\U1/net5901 ), .B(n49), .S(\U1/net27038 ), .Z(n51) );
  MUX2_X1 U182 ( .A(\U1/net5916 ), .B(\U1/net5910 ), .S(\U1/net27038 ), .Z(
        \U1/net5917 ) );
  MUX2_X1 U183 ( .A(\U1/net5922 ), .B(\U1/net5916 ), .S(\U1/net27038 ), .Z(n52) );
  MUX2_X1 U184 ( .A(net34789), .B(\U1/net5919 ), .S(\U1/net27036 ), .Z(n53) );
  MUX2_X1 U185 ( .A(n54), .B(\U1/net5922 ), .S(\U1/net27036 ), .Z(n55) );
  MUX2_X1 U186 ( .A(n117), .B(\U1/net24039 ), .S(\U1/net27024 ), .Z(n56) );
  MUX2_X1 U187 ( .A(n56), .B(net34789), .S(\U1/net27036 ), .Z(n57) );
  MUX2_X1 U188 ( .A(n119), .B(\U1/net24076 ), .S(\U1/net27024 ), .Z(n58) );
  MUX2_X1 U189 ( .A(n59), .B(n56), .S(\U1/net27036 ), .Z(n60) );
  MUX2_X1 U190 ( .A(n122), .B(n116), .S(\U1/net27024 ), .Z(n61) );
  MUX2_X1 U191 ( .A(n61), .B(n58), .S(\U1/net27036 ), .Z(n62) );
  MUX2_X1 U192 ( .A(n63), .B(n59), .S(\U1/net27036 ), .Z(n64) );
  MUX2_X1 U193 ( .A(n133), .B(n119), .S(\U1/net27024 ), .Z(n65) );
  MUX2_X1 U194 ( .A(n65), .B(n36), .S(\U1/net27036 ), .Z(n66) );
  MUX2_X1 U195 ( .A(n67), .B(n63), .S(\U1/net27036 ), .Z(n68) );
  MUX2_X1 U196 ( .A(n105), .B(n122), .S(\U1/net27024 ), .Z(n69) );
  MUX2_X1 U197 ( .A(n69), .B(n65), .S(\U1/net27036 ), .Z(n70) );
  MUX2_X1 U198 ( .A(n71), .B(n67), .S(\U1/net27036 ), .Z(n72) );
  MUX2_X1 U199 ( .A(n73), .B(n69), .S(\U1/net27034 ), .Z(n74) );
  MUX2_X1 U200 ( .A(n108), .B(n3), .S(\U1/net27022 ), .Z(n75) );
  MUX2_X1 U201 ( .A(n109), .B(n105), .S(\U1/net27022 ), .Z(n77) );
  MUX2_X1 U202 ( .A(n110), .B(n106), .S(\U1/net27022 ), .Z(n79) );
  MUX2_X1 U203 ( .A(n79), .B(n32), .S(\U1/net27034 ), .Z(n80) );
  MUX2_X1 U204 ( .A(n128), .B(n107), .S(\U1/net27022 ), .Z(n81) );
  MUX2_X1 U205 ( .A(n81), .B(n77), .S(\U1/net27034 ), .Z(n82) );
  MUX2_X1 U206 ( .A(n83), .B(n79), .S(\U1/net27034 ), .Z(n84) );
  MUX2_X1 U207 ( .A(n7), .B(n81), .S(\U1/net27034 ), .Z(n86) );
  MUX2_X1 U208 ( .A(n101), .B(n110), .S(\U1/net27022 ), .Z(n87) );
  MUX2_X1 U209 ( .A(n87), .B(n83), .S(\U1/net27034 ), .Z(n88) );
  MUX2_X1 U210 ( .A(n100), .B(n128), .S(\U1/net27022 ), .Z(n89) );
  MUX2_X1 U211 ( .A(n89), .B(n85), .S(\U1/net27034 ), .Z(n90) );
  MUX2_X1 U212 ( .A(n44), .B(n87), .S(\U1/net27034 ), .Z(n91) );
  MUX2_X1 U213 ( .A(n92), .B(n33), .S(\U1/net27034 ), .Z(n93) );
endmodule


module T2_SHIFTER_DATA_W32_1 ( A, AMOUNT, OP, S );
  input [31:0] A;
  input [31:0] AMOUNT;
  input [1:0] OP;
  output [31:0] S;
  wire   msb, n1;
  wire   [40:0] m0;
  wire   [40:0] m8;
  wire   [40:0] m16;
  wire   [40:0] m24;
  wire   [40:0] m_selected;
  wire   [2:0] op_fine;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  XOR2_X1 U2 ( .A(n1), .B(AMOUNT[2]), .Z(op_fine[2]) );
  XOR2_X1 U3 ( .A(n1), .B(AMOUNT[1]), .Z(op_fine[1]) );
  XOR2_X1 U4 ( .A(n1), .B(AMOUNT[0]), .Z(op_fine[0]) );
  MASK_GEN_DATA_W32_MASK_SIZE41_1 MASKGEN ( .OP(OP), .A(A), .MASK0({m0[40:1], 
        SYNOPSYS_UNCONNECTED__0}), .MASK8({m8[40:1], SYNOPSYS_UNCONNECTED__1}), 
        .MASK16({m16[40:1], SYNOPSYS_UNCONNECTED__2}), .MASK24({m24[40:1], 
        SYNOPSYS_UNCONNECTED__3}), .MSB(msb) );
  COARSE_SHIFT_DATA_W32_MASK_SIZE41_1 COARSESHIFT ( .MASK0({m0[40:1], 1'b0}), 
        .MASK8({m8[40:1], 1'b0}), .MASK16({m16[40:1], 1'b0}), .MASK24({
        m24[40:1], 1'b0}), .MSB(msb), .AMOUNT(AMOUNT[31:3]), .S(m_selected) );
  FINE_SHIFT_DATA_W32_MASK_SIZE41_1 FINESHIFT ( .A(m_selected), .AMOUNT(
        op_fine), .S(S) );
  OR2_X1 U1 ( .A1(OP[0]), .A2(OP[1]), .ZN(n1) );
endmodule


module ALU_DATA_W32_1_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n222, net22948, net22867, net22866, net22865, net22864, net22863,
         net22862, net22861, net22860, net22859, net22858, net22857, net22856,
         net22847, net22845, net22843, net22842, net22841, net22840, net22837,
         net22836, net22833, net22832, net22831, net22830, net22823, net22822,
         net22821, net22820, net22817, net22816, net22813, net22812, net22811,
         net22810, net22802, net22801, net22800, net22796, net22793, net22792,
         net22791, net22790, net22781, net22780, net22777, net24555, net24561,
         net24563, net24573, net24575, net33867, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221;

  AND3_X1 U1 ( .A1(n103), .A2(n104), .A3(n105), .ZN(n102) );
  AND2_X1 U2 ( .A1(net22862), .A2(net22863), .ZN(n105) );
  INV_X1 U3 ( .A(net22802), .ZN(n117) );
  AND2_X1 U4 ( .A1(net22864), .A2(net22865), .ZN(n108) );
  AND2_X1 U5 ( .A1(n200), .A2(n192), .ZN(n56) );
  NAND2_X1 U6 ( .A1(net22867), .A2(net22866), .ZN(n85) );
  AND2_X1 U7 ( .A1(net22791), .A2(net22790), .ZN(n83) );
  INV_X1 U8 ( .A(net22812), .ZN(n115) );
  INV_X1 U9 ( .A(net22813), .ZN(n116) );
  OR2_X1 U10 ( .A1(n62), .A2(n9), .ZN(n151) );
  AND4_X1 U11 ( .A1(n2), .A2(n1), .A3(net22800), .A4(net22801), .ZN(n80) );
  NAND2_X1 U12 ( .A1(n110), .A2(n3), .ZN(n109) );
  AND2_X1 U13 ( .A1(net22793), .A2(net22792), .ZN(n111) );
  INV_X1 U14 ( .A(n124), .ZN(n47) );
  AND2_X1 U15 ( .A1(net22781), .A2(net22780), .ZN(n70) );
  XNOR2_X1 U16 ( .A(B[20]), .B(A[20]), .ZN(n1) );
  OR2_X1 U17 ( .A1(n169), .A2(A[19]), .ZN(n2) );
  OR2_X1 U18 ( .A1(n166), .A2(A[23]), .ZN(n3) );
  OR2_X1 U19 ( .A1(n162), .A2(A[27]), .ZN(n4) );
  OR2_X1 U20 ( .A1(n177), .A2(A[11]), .ZN(n5) );
  AND2_X1 U21 ( .A1(net24563), .A2(net22857), .ZN(n6) );
  AND2_X1 U22 ( .A1(n207), .A2(net24573), .ZN(n7) );
  AND2_X1 U23 ( .A1(net22843), .A2(net22948), .ZN(n8) );
  AND2_X1 U24 ( .A1(n202), .A2(net22790), .ZN(n9) );
  AND2_X1 U25 ( .A1(net22841), .A2(net22842), .ZN(n10) );
  AND2_X1 U26 ( .A1(net24555), .A2(n58), .ZN(n11) );
  AND2_X1 U27 ( .A1(n110), .A2(net22865), .ZN(n12) );
  AND2_X1 U28 ( .A1(n200), .A2(net22780), .ZN(n13) );
  NAND2_X1 U29 ( .A1(n197), .A2(n196), .ZN(n14) );
  AND2_X1 U30 ( .A1(net22800), .A2(n204), .ZN(n15) );
  AND2_X1 U31 ( .A1(net22801), .A2(net22802), .ZN(n16) );
  AND2_X1 U32 ( .A1(net22810), .A2(n206), .ZN(n17) );
  AND2_X1 U33 ( .A1(net22811), .A2(net22812), .ZN(n18) );
  AND2_X1 U34 ( .A1(A[20]), .A2(n59), .ZN(n19) );
  AND2_X1 U35 ( .A1(n191), .A2(n192), .ZN(n20) );
  AND2_X1 U36 ( .A1(net22820), .A2(n209), .ZN(n21) );
  AND2_X1 U37 ( .A1(net22821), .A2(net22822), .ZN(n22) );
  AND2_X1 U38 ( .A1(net22831), .A2(net22832), .ZN(n23) );
  AND2_X1 U39 ( .A1(n5), .A2(n210), .ZN(n24) );
  AND2_X1 U40 ( .A1(n3), .A2(n203), .ZN(n25) );
  AND2_X1 U41 ( .A1(net24561), .A2(n214), .ZN(n26) );
  NAND2_X1 U42 ( .A1(A[11]), .A2(n177), .ZN(n27) );
  AND2_X1 U43 ( .A1(n130), .A2(n66), .ZN(n28) );
  NAND2_X1 U44 ( .A1(n218), .A2(n11), .ZN(n217) );
  INV_X1 U45 ( .A(net22796), .ZN(n110) );
  NOR2_X1 U46 ( .A1(n92), .A2(n91), .ZN(n75) );
  NOR2_X1 U47 ( .A1(net22836), .A2(net22837), .ZN(n89) );
  NAND2_X1 U48 ( .A1(n29), .A2(B[8]), .ZN(n212) );
  INV_X1 U49 ( .A(A[8]), .ZN(n29) );
  OAI211_X1 U50 ( .C1(n30), .C2(n31), .A(net22856), .B(net22857), .ZN(n90) );
  INV_X1 U51 ( .A(net22840), .ZN(n30) );
  INV_X1 U52 ( .A(n214), .ZN(n31) );
  NAND3_X1 U53 ( .A1(n118), .A2(n88), .A3(n87), .ZN(n119) );
  OAI21_X1 U54 ( .B1(n165), .B2(A[24]), .A(net22793), .ZN(net22796) );
  INV_X1 U55 ( .A(n60), .ZN(n32) );
  OAI21_X1 U56 ( .B1(net22821), .B2(n96), .A(n98), .ZN(n99) );
  NAND2_X1 U57 ( .A1(n124), .A2(n37), .ZN(n46) );
  AND2_X1 U58 ( .A1(n209), .A2(net22823), .ZN(n33) );
  NAND2_X1 U59 ( .A1(n213), .A2(n36), .ZN(n34) );
  AND2_X1 U60 ( .A1(n34), .A2(n35), .ZN(n211) );
  OR2_X1 U61 ( .A1(n122), .A2(n6), .ZN(n35) );
  AND2_X1 U62 ( .A1(n26), .A2(n123), .ZN(n36) );
  AND2_X1 U63 ( .A1(n209), .A2(net22823), .ZN(net33867) );
  OAI21_X1 U64 ( .B1(net22831), .B2(n93), .A(n5), .ZN(n77) );
  NAND2_X1 U65 ( .A1(n13), .A2(n140), .ZN(n37) );
  NOR2_X1 U66 ( .A1(A[4]), .A2(n154), .ZN(n38) );
  OR2_X1 U67 ( .A1(A[4]), .A2(n154), .ZN(net22948) );
  INV_X1 U68 ( .A(net22843), .ZN(n72) );
  OR2_X1 U69 ( .A1(n48), .A2(n28), .ZN(n39) );
  NAND2_X1 U70 ( .A1(n39), .A2(n40), .ZN(n156) );
  AND2_X1 U71 ( .A1(n41), .A2(n46), .ZN(n40) );
  INV_X1 U72 ( .A(n157), .ZN(n41) );
  AND2_X1 U73 ( .A1(n151), .A2(n50), .ZN(n42) );
  AND2_X1 U74 ( .A1(net22777), .A2(n144), .ZN(n43) );
  AOI21_X1 U75 ( .B1(n86), .B2(n14), .A(n72), .ZN(n87) );
  AOI21_X1 U76 ( .B1(n43), .B2(n186), .A(B[31]), .ZN(n44) );
  NAND2_X1 U77 ( .A1(n27), .A2(net22858), .ZN(n93) );
  NAND2_X1 U78 ( .A1(net22858), .A2(net22859), .ZN(n92) );
  NAND2_X1 U79 ( .A1(net33867), .A2(n94), .ZN(n76) );
  OR2_X1 U80 ( .A1(n51), .A2(n48), .ZN(n45) );
  NAND2_X1 U81 ( .A1(n45), .A2(n46), .ZN(n199) );
  OR2_X1 U82 ( .A1(n52), .A2(n47), .ZN(n48) );
  CLKBUF_X1 U83 ( .A(n220), .Z(n49) );
  NOR2_X1 U84 ( .A1(n101), .A2(n99), .ZN(n100) );
  NAND2_X1 U85 ( .A1(n151), .A2(n50), .ZN(n145) );
  NAND2_X1 U86 ( .A1(n12), .A2(n153), .ZN(n50) );
  NAND2_X1 U87 ( .A1(n215), .A2(n10), .ZN(n213) );
  INV_X1 U88 ( .A(net22845), .ZN(n113) );
  NAND2_X1 U89 ( .A1(n57), .A2(n138), .ZN(n133) );
  AND2_X1 U90 ( .A1(n130), .A2(n66), .ZN(n51) );
  NAND2_X1 U91 ( .A1(n64), .A2(n142), .ZN(n52) );
  AND3_X1 U92 ( .A1(net22856), .A2(net22842), .A3(net22857), .ZN(n88) );
  NAND2_X1 U93 ( .A1(n56), .A2(n4), .ZN(n112) );
  NOR2_X1 U94 ( .A1(n143), .A2(n44), .ZN(LE) );
  AND2_X1 U95 ( .A1(n22), .A2(n137), .ZN(n132) );
  NOR2_X1 U96 ( .A1(net22816), .A2(net22817), .ZN(n98) );
  AND2_X1 U97 ( .A1(net22791), .A2(net22792), .ZN(n54) );
  NAND2_X1 U98 ( .A1(n147), .A2(n55), .ZN(n208) );
  AND2_X1 U99 ( .A1(n148), .A2(n21), .ZN(n55) );
  AND2_X1 U100 ( .A1(n1), .A2(net22863), .ZN(n57) );
  OR2_X1 U101 ( .A1(A[2]), .A2(n184), .ZN(n58) );
  OR2_X1 U102 ( .A1(n184), .A2(A[2]), .ZN(n219) );
  INV_X1 U103 ( .A(B[20]), .ZN(n59) );
  AND2_X1 U104 ( .A1(n69), .A2(n68), .ZN(n66) );
  INV_X1 U105 ( .A(n188), .ZN(n60) );
  NAND2_X1 U106 ( .A1(n71), .A2(n70), .ZN(net22777) );
  AOI211_X1 U107 ( .C1(n74), .C2(n75), .A(n76), .B(n77), .ZN(n73) );
  AND2_X1 U108 ( .A1(n18), .A2(n57), .ZN(n134) );
  NAND2_X1 U109 ( .A1(n61), .A2(n186), .ZN(n128) );
  OR2_X1 U110 ( .A1(n157), .A2(n199), .ZN(n61) );
  NOR2_X1 U111 ( .A1(n38), .A2(net22847), .ZN(n86) );
  OAI21_X1 U112 ( .B1(n82), .B2(n112), .A(n20), .ZN(n71) );
  OAI21_X1 U113 ( .B1(n73), .B2(n95), .A(n100), .ZN(n120) );
  NAND2_X1 U114 ( .A1(n54), .A2(n159), .ZN(n62) );
  NAND2_X1 U115 ( .A1(n56), .A2(net22867), .ZN(n63) );
  INV_X1 U116 ( .A(net22830), .ZN(n114) );
  NAND2_X1 U117 ( .A1(net22833), .A2(net22832), .ZN(n91) );
  OR2_X1 U118 ( .A1(n65), .A2(n134), .ZN(n64) );
  INV_X1 U119 ( .A(n68), .ZN(n65) );
  INV_X1 U120 ( .A(B[28]), .ZN(n67) );
  AND2_X1 U121 ( .A1(n16), .A2(n145), .ZN(n142) );
  AND2_X1 U122 ( .A1(n133), .A2(n15), .ZN(n68) );
  AOI21_X1 U123 ( .B1(n84), .B2(n83), .A(n85), .ZN(n82) );
  OAI21_X1 U124 ( .B1(n78), .B2(n109), .A(n111), .ZN(n84) );
  AOI21_X1 U125 ( .B1(n79), .B2(n80), .A(n81), .ZN(n78) );
  NAND2_X1 U126 ( .A1(n120), .A2(n102), .ZN(n79) );
  AND2_X1 U127 ( .A1(n131), .A2(n17), .ZN(n69) );
  NAND3_X1 U128 ( .A1(n106), .A2(n107), .A3(n108), .ZN(n81) );
  NAND3_X1 U129 ( .A1(n113), .A2(net22948), .A3(net24555), .ZN(n118) );
  NAND3_X1 U130 ( .A1(n119), .A2(n90), .A3(n89), .ZN(n74) );
  NAND3_X1 U131 ( .A1(net22858), .A2(n114), .A3(net22859), .ZN(n94) );
  NAND3_X1 U132 ( .A1(net22810), .A2(n116), .A3(net22811), .ZN(n103) );
  NAND3_X1 U133 ( .A1(net22810), .A2(n115), .A3(net22811), .ZN(n104) );
  NAND3_X1 U134 ( .A1(net22800), .A2(n19), .A3(net22801), .ZN(n106) );
  NAND3_X1 U135 ( .A1(net22800), .A2(n117), .A3(net22801), .ZN(n107) );
  OAI211_X1 U136 ( .C1(net22820), .C2(n97), .A(net22810), .B(net22811), .ZN(
        n101) );
  NAND2_X1 U137 ( .A1(net22861), .A2(net22860), .ZN(n97) );
  NAND2_X1 U138 ( .A1(net22861), .A2(net22860), .ZN(n96) );
  NAND4_X1 U139 ( .A1(net22823), .A2(net22822), .A3(net22860), .A4(net22861), 
        .ZN(n95) );
  INV_X1 U140 ( .A(B[7]), .ZN(n121) );
  NAND2_X1 U141 ( .A1(net22830), .A2(n212), .ZN(n122) );
  INV_X1 U142 ( .A(n122), .ZN(n123) );
  AND2_X1 U143 ( .A1(net22781), .A2(n191), .ZN(n124) );
  AND2_X1 U144 ( .A1(n219), .A2(n196), .ZN(n125) );
  AND2_X1 U145 ( .A1(A[0]), .A2(n160), .ZN(n126) );
  AND2_X1 U146 ( .A1(n198), .A2(n128), .ZN(n127) );
  AND2_X1 U147 ( .A1(n33), .A2(n27), .ZN(n129) );
  NAND2_X1 U148 ( .A1(n208), .A2(n132), .ZN(n130) );
  OR2_X1 U149 ( .A1(n136), .A2(n7), .ZN(n131) );
  AND2_X1 U150 ( .A1(net22948), .A2(net22840), .ZN(n135) );
  NAND2_X1 U151 ( .A1(net24575), .A2(net22861), .ZN(n136) );
  INV_X1 U152 ( .A(n136), .ZN(n137) );
  NAND2_X1 U153 ( .A1(n205), .A2(n2), .ZN(n138) );
  AND2_X1 U154 ( .A1(net22777), .A2(n144), .ZN(n139) );
  AND2_X1 U155 ( .A1(n25), .A2(n151), .ZN(n146) );
  AND2_X1 U156 ( .A1(n54), .A2(n159), .ZN(n153) );
  AND2_X1 U157 ( .A1(n141), .A2(n152), .ZN(n140) );
  OR2_X1 U158 ( .A1(n42), .A2(n146), .ZN(n141) );
  AND2_X1 U159 ( .A1(n189), .A2(A[31]), .ZN(n143) );
  NOR2_X1 U160 ( .A1(n190), .A2(n143), .ZN(n222) );
  OR2_X1 U161 ( .A1(B[30]), .A2(n187), .ZN(n144) );
  NAND2_X1 U162 ( .A1(net22777), .A2(n144), .ZN(n189) );
  AND2_X1 U163 ( .A1(n23), .A2(n129), .ZN(n150) );
  NAND2_X1 U164 ( .A1(n211), .A2(n150), .ZN(n147) );
  OR2_X1 U165 ( .A1(n149), .A2(n24), .ZN(n148) );
  INV_X1 U166 ( .A(n129), .ZN(n149) );
  OR2_X1 U167 ( .A1(n63), .A2(n158), .ZN(n152) );
  INV_X1 U168 ( .A(B[4]), .ZN(n154) );
  CLKBUF_X1 U169 ( .A(n127), .Z(GE) );
  AND2_X1 U170 ( .A1(n187), .A2(B[30]), .ZN(n157) );
  INV_X1 U171 ( .A(net22847), .ZN(net24555) );
  INV_X1 U172 ( .A(net22816), .ZN(net24575) );
  INV_X1 U173 ( .A(net22817), .ZN(net24573) );
  INV_X1 U174 ( .A(net22836), .ZN(net24563) );
  INV_X1 U175 ( .A(net22837), .ZN(net24561) );
  AND2_X1 U176 ( .A1(n4), .A2(n201), .ZN(n158) );
  AND2_X1 U177 ( .A1(n56), .A2(net22867), .ZN(n159) );
  INV_X1 U178 ( .A(B[19]), .ZN(n169) );
  INV_X1 U179 ( .A(B[23]), .ZN(n166) );
  INV_X1 U180 ( .A(B[22]), .ZN(n167) );
  INV_X1 U181 ( .A(B[16]), .ZN(n172) );
  INV_X1 U182 ( .A(B[18]), .ZN(n170) );
  INV_X1 U183 ( .A(B[21]), .ZN(n168) );
  INV_X1 U184 ( .A(B[17]), .ZN(n171) );
  INV_X1 U185 ( .A(B[8]), .ZN(n180) );
  INV_X1 U186 ( .A(B[6]), .ZN(n181) );
  INV_X1 U187 ( .A(B[27]), .ZN(n162) );
  INV_X1 U188 ( .A(B[11]), .ZN(n177) );
  INV_X1 U189 ( .A(B[15]), .ZN(n173) );
  INV_X1 U190 ( .A(B[29]), .ZN(n161) );
  INV_X1 U191 ( .A(B[24]), .ZN(n165) );
  INV_X1 U192 ( .A(B[26]), .ZN(n163) );
  INV_X1 U193 ( .A(B[9]), .ZN(n179) );
  INV_X1 U194 ( .A(B[12]), .ZN(n176) );
  INV_X1 U195 ( .A(B[10]), .ZN(n178) );
  INV_X1 U196 ( .A(B[14]), .ZN(n174) );
  INV_X1 U197 ( .A(B[13]), .ZN(n175) );
  INV_X1 U198 ( .A(B[25]), .ZN(n164) );
  INV_X1 U199 ( .A(A[30]), .ZN(n187) );
  INV_X1 U200 ( .A(B[3]), .ZN(n183) );
  INV_X1 U201 ( .A(A[31]), .ZN(n186) );
  INV_X1 U202 ( .A(B[5]), .ZN(n182) );
  INV_X1 U203 ( .A(B[0]), .ZN(n160) );
  INV_X1 U204 ( .A(B[2]), .ZN(n184) );
  NAND2_X1 U205 ( .A1(n216), .A2(n135), .ZN(n215) );
  INV_X1 U206 ( .A(A[1]), .ZN(n188) );
  INV_X1 U207 ( .A(n221), .ZN(n185) );
  NAND2_X1 U208 ( .A1(n222), .A2(n127), .ZN(NE) );
  AOI21_X1 U209 ( .B1(n139), .B2(n186), .A(B[31]), .ZN(n190) );
  OAI211_X1 U210 ( .C1(n60), .C2(n126), .A(n194), .B(n193), .ZN(net22845) );
  OAI21_X1 U211 ( .B1(n188), .B2(n195), .A(B[1]), .ZN(n193) );
  NAND2_X1 U212 ( .A1(A[0]), .A2(n160), .ZN(n195) );
  OAI21_X1 U213 ( .B1(n156), .B2(n186), .A(B[31]), .ZN(n198) );
  XOR2_X1 U214 ( .A(n187), .B(B[30]), .Z(net22781) );
  NAND2_X1 U215 ( .A1(A[29]), .A2(n161), .ZN(n191) );
  OR2_X1 U216 ( .A1(n161), .A2(A[29]), .ZN(net22780) );
  NAND2_X1 U217 ( .A1(A[28]), .A2(n67), .ZN(n192) );
  OR2_X1 U218 ( .A1(n67), .A2(A[28]), .ZN(n200) );
  NAND2_X1 U219 ( .A1(A[27]), .A2(n162), .ZN(net22867) );
  AND2_X1 U220 ( .A1(n201), .A2(net22866), .ZN(net22791) );
  NAND2_X1 U221 ( .A1(A[26]), .A2(n163), .ZN(net22866) );
  OR2_X1 U222 ( .A1(n163), .A2(A[26]), .ZN(n201) );
  NAND2_X1 U223 ( .A1(A[25]), .A2(n164), .ZN(net22792) );
  OR2_X1 U224 ( .A1(n164), .A2(A[25]), .ZN(net22790) );
  NAND2_X1 U225 ( .A1(A[24]), .A2(n165), .ZN(net22793) );
  OR2_X1 U226 ( .A1(n165), .A2(A[24]), .ZN(n202) );
  NAND2_X1 U227 ( .A1(A[23]), .A2(n166), .ZN(net22865) );
  AND2_X1 U228 ( .A1(n203), .A2(net22864), .ZN(net22801) );
  NAND2_X1 U229 ( .A1(A[22]), .A2(n167), .ZN(net22864) );
  OR2_X1 U230 ( .A1(n167), .A2(A[22]), .ZN(n203) );
  NAND2_X1 U231 ( .A1(A[21]), .A2(n168), .ZN(net22802) );
  OR2_X1 U232 ( .A1(n168), .A2(A[21]), .ZN(net22800) );
  OR2_X1 U233 ( .A1(n59), .A2(A[20]), .ZN(n204) );
  NAND2_X1 U234 ( .A1(A[19]), .A2(n169), .ZN(net22863) );
  AND2_X1 U235 ( .A1(n205), .A2(net22862), .ZN(net22811) );
  NAND2_X1 U236 ( .A1(A[18]), .A2(n170), .ZN(net22862) );
  OR2_X1 U237 ( .A1(n170), .A2(A[18]), .ZN(n205) );
  NAND2_X1 U238 ( .A1(A[17]), .A2(n171), .ZN(net22812) );
  OR2_X1 U239 ( .A1(n171), .A2(A[17]), .ZN(net22810) );
  NAND2_X1 U240 ( .A1(n206), .A2(net22813), .ZN(net22816) );
  NAND2_X1 U241 ( .A1(A[16]), .A2(n172), .ZN(net22813) );
  OR2_X1 U242 ( .A1(n172), .A2(A[16]), .ZN(n206) );
  NAND2_X1 U243 ( .A1(A[15]), .A2(n173), .ZN(net22861) );
  NOR2_X1 U244 ( .A1(n173), .A2(A[15]), .ZN(net22817) );
  AND2_X1 U245 ( .A1(n207), .A2(net22860), .ZN(net22821) );
  NAND2_X1 U246 ( .A1(A[14]), .A2(n174), .ZN(net22860) );
  OR2_X1 U247 ( .A1(n174), .A2(A[14]), .ZN(n207) );
  NAND2_X1 U248 ( .A1(A[13]), .A2(n175), .ZN(net22822) );
  OR2_X1 U249 ( .A1(n175), .A2(A[13]), .ZN(net22820) );
  NAND2_X1 U250 ( .A1(A[12]), .A2(n176), .ZN(net22823) );
  OR2_X1 U251 ( .A1(A[12]), .A2(n176), .ZN(n209) );
  NAND2_X1 U252 ( .A1(A[11]), .A2(n177), .ZN(net22859) );
  AND2_X1 U253 ( .A1(n210), .A2(net22858), .ZN(net22831) );
  NAND2_X1 U254 ( .A1(A[10]), .A2(n178), .ZN(net22858) );
  OR2_X1 U255 ( .A1(n178), .A2(A[10]), .ZN(n210) );
  NAND2_X1 U256 ( .A1(A[9]), .A2(n179), .ZN(net22832) );
  OR2_X1 U257 ( .A1(n179), .A2(A[9]), .ZN(net22830) );
  NAND2_X1 U258 ( .A1(n212), .A2(net22833), .ZN(net22836) );
  NAND2_X1 U259 ( .A1(A[8]), .A2(n180), .ZN(net22833) );
  NAND2_X1 U260 ( .A1(A[7]), .A2(n121), .ZN(net22857) );
  NOR2_X1 U261 ( .A1(n121), .A2(A[7]), .ZN(net22837) );
  AND2_X1 U262 ( .A1(n214), .A2(net22856), .ZN(net22841) );
  NAND2_X1 U263 ( .A1(A[6]), .A2(n181), .ZN(net22856) );
  OR2_X1 U264 ( .A1(n181), .A2(A[6]), .ZN(n214) );
  NAND2_X1 U265 ( .A1(A[5]), .A2(n182), .ZN(net22842) );
  OR2_X1 U266 ( .A1(n182), .A2(A[5]), .ZN(net22840) );
  NAND3_X1 U267 ( .A1(n217), .A2(n197), .A3(n8), .ZN(n216) );
  NAND2_X1 U268 ( .A1(A[4]), .A2(n154), .ZN(net22843) );
  NAND2_X1 U269 ( .A1(A[3]), .A2(n183), .ZN(n197) );
  NOR2_X1 U270 ( .A1(A[3]), .A2(n183), .ZN(net22847) );
  OAI211_X1 U271 ( .C1(n32), .C2(n49), .A(n125), .B(n185), .ZN(n218) );
  AND2_X1 U272 ( .A1(n58), .A2(n196), .ZN(n194) );
  NAND2_X1 U273 ( .A1(A[2]), .A2(n184), .ZN(n196) );
  AOI21_X1 U274 ( .B1(n188), .B2(n220), .A(B[1]), .ZN(n221) );
  NOR2_X1 U275 ( .A1(n160), .A2(A[0]), .ZN(n220) );
endmodule


module ALU_DATA_W32_1 ( .FUNC({\FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), A, 
        B, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   \t2_logic_op[2] , N80, N81, N82, n80, n81, n101, n105, n111, n125,
         n128, net23818, net23819, net23821, net23856, net26984, net26982,
         net26980, net26988, net26986, net26996, net26994, net27002, net27000,
         net26998, net27008, net27006, net27004, net33642, net33774, net33873,
         net34641, net34699, net34897, net35350, net35616, net34607, n89,
         net35375, net35257, net34615, net23817, n87, n86, net35261, net23816,
         net34671, net34670, net40015, net40353, net40321, net40071, net40038,
         net35407, net35365, net35271, net35241, n94, n93, n91, n90, n82, n130,
         n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n39, n40, n41, n43, n44, n45, n46, n48,
         n49, n50, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n72, n73, n76, n77, n78, n79, n83, n84,
         n85, n88, n92, n95, n96, n97, n99, n100, n102, n103, n104, n106, n108,
         n114, n116, n117, n118, n119, n120, n122, n123, n124, n126, n127,
         n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245;
  wire   [3:0] FUNC;
  wire   [31:0] p4_adder_b;
  wire   [31:0] p4_adder_s;
  wire   [31:0] t2_logic_s;
  wire   [31:0] t2_shifter_s;
  assign RES[5] = net23856;
  assign RES[20] = net34699;

  P4_ADDER_NBIT32_1 P4_ADDER_U ( .A({n185, A[30:28], n114, n116, A[25:22], n72, 
        A[20:19], n76, A[17], n133, A[15:11], n188, n135, A[8], n78, n198, 
        A[5], n200, n203, n205, n201, n204}), .B(p4_adder_b), .Cin(net26984), 
        .S(p4_adder_s) );
  T2_LOGIC_DATA_W32_1 T2_LOGIC_U ( .OP({net23821, \t2_logic_op[2] , 
        \t2_logic_op[2] , 1'b0}), .A({n185, A[30:28], n114, n116, A[25:22], 
        n72, A[20:19], n76, A[17], n133, A[15:11], n188, n135, A[8], n78, n198, 
        A[5], n200, n203, n205, n201, n204}), .B({n96, n97, n8, n70, B[27], 
        n131, n178, n186, n99, n102, n123, n20, n73, n122, B[17:16], n15, n16, 
        n69, n77, n9, n19, n68, n23, n18, n197, n190, n199, n194, n196, n195, 
        n22}), .S(t2_logic_s) );
  T2_SHIFTER_DATA_W32_1 T2_SHIFTER_U ( .A({A[31:28], n114, n116, A[25:22], n72, 
        A[20:19], n76, A[17], n133, A[15:11], n188, n135, A[8], n78, n198, 
        A[5], n200, n203, n205, A[1], n204}), .AMOUNT({B[31:7], n197, B[5:4], 
        n194, n196, n195, n22}), .OP({net35350, net23819}), .S(t2_shifter_s)
         );
  ALU_DATA_W32_1_DW01_cmp6_0 r53 ( .A({n96, B[30], n8, B[28:26], n178, n186, 
        n99, n102, n123, B[20], n73, B[18:16], n15, B[14], n69, n77, n120, n19, 
        n68, B[8:6], n124, B[4:0]}), .B(A), .TC(1'b0), .LE(N80), .GE(N81), 
        .NE(N82) );
  NAND3_X1 U160 ( .A1(net23817), .A2(net34615), .A3(net35257), .ZN(n86) );
  NAND3_X1 U155 ( .A1(n91), .A2(n87), .A3(n130), .ZN(n94) );
  BUF_X1 U3 ( .A(n93), .Z(net26998) );
  BUF_X1 U4 ( .A(n94), .Z(net27006) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(p4_adder_b[7]) );
  NOR2_X1 U6 ( .A1(net35407), .A2(n86), .ZN(net35365) );
  NAND2_X1 U7 ( .A1(t2_logic_s[15]), .A2(net26994), .ZN(n119) );
  NAND2_X1 U8 ( .A1(t2_logic_s[20]), .A2(net26994), .ZN(net34671) );
  NAND2_X1 U9 ( .A1(t2_logic_s[21]), .A2(net26994), .ZN(n129) );
  OR2_X1 U10 ( .A1(net35365), .A2(net26984), .ZN(n93) );
  AND4_X1 U11 ( .A1(FUNC[0]), .A2(net35271), .A3(net34615), .A4(net23817), 
        .ZN(n1) );
  BUF_X1 U12 ( .A(n93), .Z(net27000) );
  BUF_X1 U13 ( .A(n90), .Z(net26994) );
  BUF_X1 U14 ( .A(B[12]), .Z(n77) );
  NAND2_X1 U15 ( .A1(net23818), .A2(net33642), .ZN(n80) );
  BUF_X1 U16 ( .A(net35261), .Z(net23817) );
  NOR2_X1 U17 ( .A1(n36), .A2(n31), .ZN(n2) );
  NOR2_X1 U18 ( .A1(n36), .A2(n37), .ZN(n3) );
  NAND2_X1 U19 ( .A1(t2_logic_s[12]), .A2(net26996), .ZN(n4) );
  NAND2_X1 U20 ( .A1(t2_logic_s[14]), .A2(net26994), .ZN(n5) );
  NAND2_X1 U21 ( .A1(t2_logic_s[13]), .A2(net26996), .ZN(n6) );
  CLKBUF_X1 U22 ( .A(n94), .Z(net27008) );
  CLKBUF_X1 U23 ( .A(B[29]), .Z(n8) );
  CLKBUF_X1 U24 ( .A(n100), .Z(n9) );
  BUF_X1 U25 ( .A(B[11]), .Z(n100) );
  OR2_X1 U26 ( .A1(net26982), .A2(B[7]), .ZN(n10) );
  OR2_X1 U27 ( .A1(n239), .A2(n1), .ZN(n11) );
  AND4_X1 U28 ( .A1(n85), .A2(n26), .A3(n86), .A4(n88), .ZN(net26986) );
  AND2_X2 U29 ( .A1(FUNC[1]), .A2(net40353), .ZN(n12) );
  INV_X1 U30 ( .A(net34615), .ZN(n13) );
  AND4_X1 U31 ( .A1(n85), .A2(n26), .A3(n86), .A4(n17), .ZN(n14) );
  AND4_X1 U32 ( .A1(n85), .A2(n26), .A3(n86), .A4(n17), .ZN(n92) );
  BUF_X1 U33 ( .A(B[0]), .Z(net33774) );
  INV_X1 U34 ( .A(n231), .ZN(n15) );
  AOI21_X2 U35 ( .B1(n12), .B2(net34607), .A(net35407), .ZN(n85) );
  INV_X1 U36 ( .A(n232), .ZN(n16) );
  NAND2_X1 U37 ( .A1(net40038), .A2(FUNC[1]), .ZN(net35241) );
  AND2_X1 U38 ( .A1(net40321), .A2(n87), .ZN(n17) );
  AND2_X1 U39 ( .A1(net40321), .A2(n87), .ZN(n88) );
  INV_X1 U40 ( .A(n79), .ZN(net26984) );
  BUF_X1 U41 ( .A(B[9]), .Z(n68) );
  CLKBUF_X1 U42 ( .A(FUNC[3]), .Z(net40071) );
  INV_X1 U43 ( .A(n242), .ZN(n199) );
  INV_X1 U44 ( .A(n239), .ZN(n18) );
  BUF_X1 U45 ( .A(B[10]), .Z(n19) );
  INV_X1 U46 ( .A(n226), .ZN(n20) );
  CLKBUF_X1 U47 ( .A(B[19]), .Z(n21) );
  INV_X1 U48 ( .A(n87), .ZN(net23819) );
  CLKBUF_X1 U49 ( .A(net33774), .Z(n22) );
  INV_X1 U50 ( .A(n238), .ZN(n23) );
  OR2_X1 U51 ( .A1(n24), .A2(n25), .ZN(RES[12]) );
  AND2_X1 U52 ( .A1(t2_shifter_s[12]), .A2(net27004), .ZN(n24) );
  NAND2_X1 U53 ( .A1(n4), .A2(n50), .ZN(n25) );
  AND2_X2 U54 ( .A1(net35241), .A2(n82), .ZN(n26) );
  INV_X1 U55 ( .A(n26), .ZN(n90) );
  NOR2_X1 U56 ( .A1(FUNC[1]), .A2(net23816), .ZN(n89) );
  NAND2_X1 U57 ( .A1(net23817), .A2(N80), .ZN(n28) );
  NAND2_X1 U58 ( .A1(n29), .A2(n28), .ZN(n27) );
  NAND2_X1 U59 ( .A1(N82), .A2(FUNC[1]), .ZN(n29) );
  INV_X1 U60 ( .A(t2_logic_s[30]), .ZN(n31) );
  NAND2_X1 U61 ( .A1(n34), .A2(n33), .ZN(RES[30]) );
  NAND2_X1 U62 ( .A1(net27000), .A2(p4_adder_s[30]), .ZN(n33) );
  NOR2_X1 U63 ( .A1(n30), .A2(n2), .ZN(n34) );
  AND2_X1 U64 ( .A1(net27008), .A2(t2_shifter_s[30]), .ZN(n30) );
  INV_X1 U65 ( .A(net26996), .ZN(n36) );
  INV_X1 U66 ( .A(t2_logic_s[23]), .ZN(n37) );
  NAND2_X1 U67 ( .A1(n40), .A2(n39), .ZN(RES[23]) );
  NAND2_X1 U68 ( .A1(net27002), .A2(p4_adder_s[23]), .ZN(n39) );
  NOR2_X1 U69 ( .A1(n35), .A2(n3), .ZN(n40) );
  AND2_X1 U70 ( .A1(net27004), .A2(t2_shifter_s[23]), .ZN(n35) );
  NAND2_X1 U71 ( .A1(t2_shifter_s[29]), .A2(net27006), .ZN(n41) );
  NAND2_X1 U72 ( .A1(t2_logic_s[29]), .A2(net26994), .ZN(n43) );
  OR2_X1 U73 ( .A1(n45), .A2(n44), .ZN(RES[29]) );
  AND2_X1 U74 ( .A1(p4_adder_s[29]), .A2(net27000), .ZN(n44) );
  NAND2_X1 U75 ( .A1(n41), .A2(n43), .ZN(n45) );
  NAND2_X1 U76 ( .A1(p4_adder_s[13]), .A2(net26998), .ZN(n46) );
  NAND2_X1 U77 ( .A1(t2_shifter_s[13]), .A2(net27004), .ZN(n48) );
  NAND2_X1 U78 ( .A1(n48), .A2(n49), .ZN(RES[13]) );
  AND2_X1 U79 ( .A1(n6), .A2(n46), .ZN(n49) );
  NAND2_X1 U80 ( .A1(p4_adder_s[12]), .A2(net26998), .ZN(n50) );
  NAND2_X1 U81 ( .A1(p4_adder_s[14]), .A2(net26998), .ZN(n52) );
  NAND2_X1 U82 ( .A1(t2_shifter_s[14]), .A2(net27004), .ZN(n54) );
  NAND2_X1 U83 ( .A1(n54), .A2(n55), .ZN(RES[14]) );
  AND2_X1 U84 ( .A1(n5), .A2(n52), .ZN(n55) );
  OAI211_X1 U85 ( .C1(n128), .C2(net33873), .A(n202), .B(n125), .ZN(RES[0]) );
  AND4_X2 U86 ( .A1(n17), .A2(n86), .A3(n85), .A4(n26), .ZN(net26988) );
  OAI222_X1 U87 ( .A1(n56), .A2(n57), .B1(n58), .B2(n59), .C1(n60), .C2(n36), 
        .ZN(RES[16]) );
  INV_X1 U88 ( .A(p4_adder_s[16]), .ZN(n56) );
  INV_X1 U89 ( .A(n93), .ZN(n57) );
  INV_X1 U90 ( .A(t2_shifter_s[16]), .ZN(n58) );
  INV_X1 U91 ( .A(n94), .ZN(n59) );
  INV_X1 U92 ( .A(t2_logic_s[16]), .ZN(n60) );
  OAI222_X1 U93 ( .A1(n61), .A2(n57), .B1(n62), .B2(n59), .C1(n63), .C2(n36), 
        .ZN(RES[26]) );
  INV_X1 U94 ( .A(p4_adder_s[26]), .ZN(n61) );
  INV_X1 U95 ( .A(t2_shifter_s[26]), .ZN(n62) );
  INV_X1 U96 ( .A(t2_logic_s[26]), .ZN(n63) );
  OAI222_X1 U97 ( .A1(n64), .A2(n57), .B1(n65), .B2(n59), .C1(n66), .C2(n36), 
        .ZN(net23856) );
  INV_X1 U98 ( .A(p4_adder_s[5]), .ZN(n64) );
  INV_X1 U99 ( .A(t2_shifter_s[5]), .ZN(n65) );
  INV_X1 U100 ( .A(t2_logic_s[5]), .ZN(n66) );
  INV_X1 U101 ( .A(FUNC[2]), .ZN(net34615) );
  CLKBUF_X1 U102 ( .A(n90), .Z(net26996) );
  BUF_X1 U103 ( .A(n93), .Z(net27002) );
  NOR2_X1 U104 ( .A1(net40071), .A2(FUNC[2]), .ZN(net40038) );
  BUF_X1 U105 ( .A(n94), .Z(net27004) );
  NAND2_X1 U106 ( .A1(net35271), .A2(n67), .ZN(n130) );
  INV_X1 U107 ( .A(net40321), .ZN(n67) );
  INV_X1 U108 ( .A(FUNC[3]), .ZN(net35271) );
  INV_X1 U109 ( .A(net35271), .ZN(net35407) );
  NAND4_X1 U110 ( .A1(net35271), .A2(net23816), .A3(net35261), .A4(FUNC[2]), 
        .ZN(n82) );
  INV_X1 U111 ( .A(net35350), .ZN(n91) );
  INV_X1 U112 ( .A(FUNC[1]), .ZN(net35261) );
  INV_X1 U113 ( .A(n233), .ZN(n69) );
  INV_X1 U114 ( .A(n218), .ZN(n70) );
  NAND3_X1 U115 ( .A1(n164), .A2(n163), .A3(n165), .ZN(RES[1]) );
  BUF_X2 U116 ( .A(A[21]), .Z(n72) );
  INV_X1 U117 ( .A(n227), .ZN(n73) );
  CLKBUF_X1 U118 ( .A(A[6]), .Z(n198) );
  NAND3_X1 U119 ( .A1(n136), .A2(n137), .A3(n138), .ZN(RES[2]) );
  NAND3_X1 U120 ( .A1(n161), .A2(n160), .A3(n162), .ZN(RES[3]) );
  BUF_X2 U121 ( .A(A[18]), .Z(n76) );
  BUF_X2 U122 ( .A(A[7]), .Z(n78) );
  NAND3_X1 U123 ( .A1(net33642), .A2(net34615), .A3(net35616), .ZN(n81) );
  MUX2_X1 U124 ( .A(net26984), .B(n84), .S(net33774), .Z(p4_adder_b[0]) );
  NAND2_X1 U125 ( .A1(net34615), .A2(net35407), .ZN(net33873) );
  NAND4_X1 U126 ( .A1(n85), .A2(n88), .A3(n86), .A4(n26), .ZN(n84) );
  NAND2_X1 U127 ( .A1(n89), .A2(FUNC[2]), .ZN(net40321) );
  NAND2_X1 U128 ( .A1(net35261), .A2(FUNC[0]), .ZN(n83) );
  OR3_X1 U129 ( .A1(FUNC[2]), .A2(net35407), .A3(n83), .ZN(n79) );
  OR3_X2 U130 ( .A1(n13), .A2(net40071), .A3(n83), .ZN(net26982) );
  OR3_X2 U131 ( .A1(FUNC[2]), .A2(net40071), .A3(n83), .ZN(net26980) );
  INV_X1 U132 ( .A(FUNC[3]), .ZN(net40353) );
  BUF_X1 U133 ( .A(net34897), .Z(net34641) );
  CLKBUF_X1 U134 ( .A(net35257), .Z(net40015) );
  NAND2_X1 U135 ( .A1(p4_adder_s[20]), .A2(net27000), .ZN(n95) );
  NAND3_X1 U136 ( .A1(n95), .A2(net34670), .A3(net34671), .ZN(net34699) );
  AOI22_X1 U137 ( .A1(n27), .A2(net40015), .B1(N81), .B2(n89), .ZN(n128) );
  NAND2_X1 U138 ( .A1(t2_shifter_s[20]), .A2(net27006), .ZN(net34670) );
  INV_X1 U139 ( .A(FUNC[0]), .ZN(net23816) );
  CLKBUF_X1 U140 ( .A(net23816), .Z(net35257) );
  AND2_X1 U141 ( .A1(net23816), .A2(FUNC[2]), .ZN(net35375) );
  AND2_X1 U142 ( .A1(FUNC[2]), .A2(FUNC[0]), .ZN(net34607) );
  NAND2_X1 U143 ( .A1(net35375), .A2(n12), .ZN(n87) );
  INV_X1 U144 ( .A(net40015), .ZN(net35616) );
  CLKBUF_X1 U145 ( .A(n12), .Z(net33642) );
  AND2_X1 U146 ( .A1(n12), .A2(net34607), .ZN(net35350) );
  CLKBUF_X1 U147 ( .A(B[31]), .Z(n96) );
  INV_X1 U148 ( .A(n216), .ZN(n97) );
  NAND3_X1 U149 ( .A1(n169), .A2(n170), .A3(n171), .ZN(RES[4]) );
  CLKBUF_X1 U150 ( .A(n14), .Z(net34897) );
  INV_X1 U151 ( .A(n223), .ZN(n99) );
  BUF_X1 U152 ( .A(B[3]), .Z(n194) );
  INV_X1 U153 ( .A(n224), .ZN(n102) );
  AND2_X1 U154 ( .A1(n139), .A2(n141), .ZN(n103) );
  NAND2_X1 U156 ( .A1(n140), .A2(n103), .ZN(RES[6]) );
  AND2_X1 U157 ( .A1(n155), .A2(n157), .ZN(n104) );
  NAND2_X1 U158 ( .A1(n156), .A2(n104), .ZN(RES[8]) );
  AND2_X1 U159 ( .A1(n152), .A2(n154), .ZN(n106) );
  NAND2_X1 U161 ( .A1(n153), .A2(n106), .ZN(RES[9]) );
  NAND3_X1 U162 ( .A1(n192), .A2(n191), .A3(n193), .ZN(RES[11]) );
  AND2_X1 U163 ( .A1(n166), .A2(n168), .ZN(n108) );
  NAND2_X1 U164 ( .A1(n167), .A2(n108), .ZN(RES[7]) );
  NAND3_X1 U165 ( .A1(n147), .A2(n146), .A3(n148), .ZN(RES[17]) );
  NAND3_X1 U166 ( .A1(n144), .A2(n143), .A3(n145), .ZN(RES[18]) );
  NAND3_X1 U167 ( .A1(n176), .A2(n175), .A3(n177), .ZN(RES[10]) );
  NAND3_X1 U168 ( .A1(n149), .A2(n150), .A3(n151), .ZN(RES[19]) );
  CLKBUF_X3 U169 ( .A(A[27]), .Z(n114) );
  NAND3_X1 U170 ( .A1(n117), .A2(n118), .A3(n119), .ZN(RES[15]) );
  CLKBUF_X3 U171 ( .A(A[26]), .Z(n116) );
  NAND2_X1 U172 ( .A1(p4_adder_s[15]), .A2(net26998), .ZN(n117) );
  NAND2_X1 U173 ( .A1(t2_shifter_s[15]), .A2(net27004), .ZN(n118) );
  INV_X1 U174 ( .A(n235), .ZN(n120) );
  NAND3_X1 U175 ( .A1(n126), .A2(n127), .A3(n129), .ZN(RES[21]) );
  INV_X1 U176 ( .A(n228), .ZN(n122) );
  INV_X1 U177 ( .A(n225), .ZN(n123) );
  INV_X1 U178 ( .A(n241), .ZN(n124) );
  NAND2_X1 U179 ( .A1(p4_adder_s[21]), .A2(net27000), .ZN(n126) );
  NAND2_X1 U180 ( .A1(t2_shifter_s[21]), .A2(net27006), .ZN(n127) );
  INV_X1 U181 ( .A(n220), .ZN(n131) );
  INV_X1 U182 ( .A(A[16]), .ZN(n132) );
  INV_X1 U183 ( .A(n132), .ZN(n133) );
  INV_X1 U184 ( .A(A[9]), .ZN(n134) );
  INV_X1 U185 ( .A(n134), .ZN(n135) );
  NAND2_X1 U186 ( .A1(p4_adder_s[2]), .A2(net27000), .ZN(n136) );
  NAND2_X1 U187 ( .A1(t2_shifter_s[2]), .A2(net27006), .ZN(n137) );
  NAND2_X1 U188 ( .A1(t2_logic_s[2]), .A2(net26994), .ZN(n138) );
  NAND2_X1 U189 ( .A1(p4_adder_s[6]), .A2(net27002), .ZN(n139) );
  NAND2_X1 U190 ( .A1(t2_shifter_s[6]), .A2(net27008), .ZN(n140) );
  NAND2_X1 U191 ( .A1(t2_logic_s[6]), .A2(net26994), .ZN(n141) );
  NAND3_X1 U192 ( .A1(n182), .A2(n183), .A3(n184), .ZN(RES[24]) );
  NAND2_X1 U193 ( .A1(p4_adder_s[18]), .A2(net26998), .ZN(n143) );
  NAND2_X1 U194 ( .A1(t2_shifter_s[18]), .A2(net27004), .ZN(n144) );
  NAND2_X1 U195 ( .A1(t2_logic_s[18]), .A2(net26994), .ZN(n145) );
  NAND2_X1 U196 ( .A1(p4_adder_s[17]), .A2(net26998), .ZN(n146) );
  NAND2_X1 U197 ( .A1(t2_shifter_s[17]), .A2(net27004), .ZN(n147) );
  NAND2_X1 U198 ( .A1(t2_logic_s[17]), .A2(net26996), .ZN(n148) );
  NAND2_X1 U199 ( .A1(p4_adder_s[19]), .A2(net26998), .ZN(n149) );
  NAND2_X1 U200 ( .A1(t2_shifter_s[19]), .A2(net27004), .ZN(n150) );
  NAND2_X1 U201 ( .A1(t2_logic_s[19]), .A2(net26994), .ZN(n151) );
  NAND2_X1 U202 ( .A1(p4_adder_s[9]), .A2(net27002), .ZN(n152) );
  NAND2_X1 U203 ( .A1(t2_shifter_s[9]), .A2(net27008), .ZN(n153) );
  NAND2_X1 U204 ( .A1(t2_logic_s[9]), .A2(net26996), .ZN(n154) );
  NAND2_X1 U205 ( .A1(p4_adder_s[8]), .A2(net27002), .ZN(n155) );
  NAND2_X1 U206 ( .A1(t2_shifter_s[8]), .A2(net27008), .ZN(n156) );
  NAND2_X1 U207 ( .A1(t2_logic_s[8]), .A2(net26994), .ZN(n157) );
  NAND3_X1 U208 ( .A1(n179), .A2(n180), .A3(n181), .ZN(RES[27]) );
  NAND3_X1 U209 ( .A1(n172), .A2(n173), .A3(n174), .ZN(RES[25]) );
  NAND2_X1 U210 ( .A1(p4_adder_s[3]), .A2(net27002), .ZN(n160) );
  NAND2_X1 U211 ( .A1(t2_shifter_s[3]), .A2(net27008), .ZN(n161) );
  NAND2_X1 U212 ( .A1(t2_logic_s[3]), .A2(net26996), .ZN(n162) );
  NAND2_X1 U213 ( .A1(p4_adder_s[1]), .A2(net26998), .ZN(n163) );
  NAND2_X1 U214 ( .A1(t2_shifter_s[1]), .A2(net27004), .ZN(n164) );
  NAND2_X1 U215 ( .A1(t2_logic_s[1]), .A2(net26994), .ZN(n165) );
  NAND2_X1 U216 ( .A1(p4_adder_s[7]), .A2(net27002), .ZN(n166) );
  NAND2_X1 U217 ( .A1(t2_shifter_s[7]), .A2(net27008), .ZN(n167) );
  NAND2_X1 U218 ( .A1(t2_logic_s[7]), .A2(net26994), .ZN(n168) );
  NAND2_X1 U219 ( .A1(p4_adder_s[4]), .A2(net27002), .ZN(n169) );
  NAND2_X1 U220 ( .A1(t2_shifter_s[4]), .A2(net27008), .ZN(n170) );
  NAND2_X1 U221 ( .A1(t2_logic_s[4]), .A2(net26994), .ZN(n171) );
  NAND2_X1 U222 ( .A1(p4_adder_s[25]), .A2(net27000), .ZN(n172) );
  NAND2_X1 U223 ( .A1(t2_shifter_s[25]), .A2(net27006), .ZN(n173) );
  NAND2_X1 U224 ( .A1(t2_logic_s[25]), .A2(net26996), .ZN(n174) );
  NAND2_X1 U225 ( .A1(p4_adder_s[10]), .A2(net26998), .ZN(n175) );
  NAND2_X1 U226 ( .A1(t2_shifter_s[10]), .A2(net27004), .ZN(n176) );
  NAND2_X1 U227 ( .A1(t2_logic_s[10]), .A2(net26994), .ZN(n177) );
  INV_X1 U228 ( .A(n221), .ZN(n178) );
  NAND2_X1 U229 ( .A1(p4_adder_s[27]), .A2(net27000), .ZN(n179) );
  NAND2_X1 U230 ( .A1(t2_shifter_s[27]), .A2(net27006), .ZN(n180) );
  NAND2_X1 U231 ( .A1(t2_logic_s[27]), .A2(net26994), .ZN(n181) );
  NAND2_X1 U232 ( .A1(p4_adder_s[24]), .A2(net27000), .ZN(n182) );
  NAND2_X1 U233 ( .A1(t2_shifter_s[24]), .A2(net27006), .ZN(n183) );
  NAND2_X1 U234 ( .A1(t2_logic_s[24]), .A2(net26994), .ZN(n184) );
  CLKBUF_X1 U235 ( .A(A[31]), .Z(n185) );
  INV_X1 U236 ( .A(n222), .ZN(n186) );
  INV_X1 U237 ( .A(A[10]), .ZN(n187) );
  INV_X1 U238 ( .A(n187), .ZN(n188) );
  CLKBUF_X1 U239 ( .A(B[2]), .Z(n189) );
  INV_X1 U240 ( .A(n241), .ZN(n190) );
  NAND2_X1 U241 ( .A1(p4_adder_s[11]), .A2(net26998), .ZN(n191) );
  NAND2_X1 U242 ( .A1(t2_shifter_s[11]), .A2(net27004), .ZN(n192) );
  NAND2_X1 U243 ( .A1(t2_logic_s[11]), .A2(net26996), .ZN(n193) );
  BUF_X2 U244 ( .A(B[6]), .Z(n197) );
  CLKBUF_X1 U245 ( .A(B[1]), .Z(n195) );
  INV_X1 U246 ( .A(n244), .ZN(n196) );
  CLKBUF_X1 U247 ( .A(A[3]), .Z(n203) );
  CLKBUF_X1 U248 ( .A(A[4]), .Z(n200) );
  CLKBUF_X1 U249 ( .A(A[1]), .Z(n201) );
  NAND2_X1 U250 ( .A1(t2_shifter_s[0]), .A2(net27004), .ZN(n202) );
  INV_X1 U251 ( .A(n80), .ZN(net23821) );
  OAI22_X1 U252 ( .A1(n197), .A2(net26980), .B1(net26986), .B2(n240), .ZN(
        p4_adder_b[6]) );
  INV_X1 U253 ( .A(n197), .ZN(n240) );
  INV_X1 U254 ( .A(B[7]), .ZN(n239) );
  OAI22_X1 U255 ( .A1(B[16]), .A2(net26980), .B1(n14), .B2(n230), .ZN(
        p4_adder_b[16]) );
  INV_X1 U256 ( .A(B[16]), .ZN(n230) );
  OAI22_X1 U257 ( .A1(B[17]), .A2(net26980), .B1(n1), .B2(n229), .ZN(
        p4_adder_b[17]) );
  INV_X1 U258 ( .A(B[17]), .ZN(n229) );
  OAI22_X1 U259 ( .A1(n21), .A2(net26980), .B1(n1), .B2(n227), .ZN(
        p4_adder_b[19]) );
  INV_X1 U260 ( .A(n21), .ZN(n227) );
  OAI22_X1 U261 ( .A1(B[18]), .A2(net26982), .B1(n14), .B2(n228), .ZN(
        p4_adder_b[18]) );
  INV_X1 U262 ( .A(B[18]), .ZN(n228) );
  OAI22_X1 U263 ( .A1(B[21]), .A2(net26980), .B1(net26988), .B2(n225), .ZN(
        p4_adder_b[21]) );
  INV_X1 U264 ( .A(B[21]), .ZN(n225) );
  OAI22_X1 U265 ( .A1(B[23]), .A2(net26980), .B1(n223), .B2(n1), .ZN(
        p4_adder_b[23]) );
  INV_X1 U266 ( .A(B[23]), .ZN(n223) );
  OAI22_X1 U267 ( .A1(B[20]), .A2(net26982), .B1(net26988), .B2(n226), .ZN(
        p4_adder_b[20]) );
  INV_X1 U268 ( .A(B[20]), .ZN(n226) );
  OAI22_X1 U269 ( .A1(n102), .A2(net26980), .B1(n14), .B2(n224), .ZN(
        p4_adder_b[22]) );
  INV_X1 U270 ( .A(B[22]), .ZN(n224) );
  OAI22_X1 U271 ( .A1(n178), .A2(net26982), .B1(net26986), .B2(n221), .ZN(
        p4_adder_b[25]) );
  INV_X1 U272 ( .A(B[25]), .ZN(n221) );
  OAI22_X1 U273 ( .A1(n186), .A2(net26980), .B1(net34897), .B2(n222), .ZN(
        p4_adder_b[24]) );
  INV_X1 U274 ( .A(B[24]), .ZN(n222) );
  OAI22_X1 U275 ( .A1(B[27]), .A2(net26982), .B1(n14), .B2(n219), .ZN(
        p4_adder_b[27]) );
  INV_X1 U276 ( .A(B[27]), .ZN(n219) );
  OAI22_X1 U277 ( .A1(n131), .A2(net26982), .B1(net26986), .B2(n220), .ZN(
        p4_adder_b[26]) );
  INV_X1 U278 ( .A(B[26]), .ZN(n220) );
  OAI22_X1 U279 ( .A1(B[13]), .A2(net26982), .B1(n233), .B2(n1), .ZN(
        p4_adder_b[13]) );
  INV_X1 U280 ( .A(B[13]), .ZN(n233) );
  OAI22_X1 U281 ( .A1(n77), .A2(net26982), .B1(n92), .B2(n234), .ZN(
        p4_adder_b[12]) );
  INV_X1 U282 ( .A(n77), .ZN(n234) );
  OAI22_X1 U283 ( .A1(B[15]), .A2(net26980), .B1(net26988), .B2(n231), .ZN(
        p4_adder_b[15]) );
  INV_X1 U284 ( .A(B[15]), .ZN(n231) );
  OAI22_X1 U285 ( .A1(B[8]), .A2(net26982), .B1(n92), .B2(n238), .ZN(
        p4_adder_b[8]) );
  INV_X1 U286 ( .A(B[8]), .ZN(n238) );
  OAI22_X1 U287 ( .A1(n68), .A2(net26980), .B1(n92), .B2(n237), .ZN(
        p4_adder_b[9]) );
  INV_X1 U288 ( .A(n68), .ZN(n237) );
  OAI22_X1 U289 ( .A1(n9), .A2(net26980), .B1(net26986), .B2(n235), .ZN(
        p4_adder_b[11]) );
  INV_X1 U290 ( .A(n100), .ZN(n235) );
  OAI22_X1 U291 ( .A1(B[14]), .A2(net26982), .B1(net26988), .B2(n232), .ZN(
        p4_adder_b[14]) );
  INV_X1 U292 ( .A(B[14]), .ZN(n232) );
  OAI22_X1 U293 ( .A1(n19), .A2(net26982), .B1(n92), .B2(n236), .ZN(
        p4_adder_b[10]) );
  INV_X1 U294 ( .A(n19), .ZN(n236) );
  OAI22_X1 U295 ( .A1(n70), .A2(net26980), .B1(n14), .B2(n218), .ZN(
        p4_adder_b[28]) );
  INV_X1 U296 ( .A(B[28]), .ZN(n218) );
  OAI22_X1 U297 ( .A1(n8), .A2(net26980), .B1(net34641), .B2(n217), .ZN(
        p4_adder_b[29]) );
  INV_X1 U298 ( .A(n8), .ZN(n217) );
  OAI22_X1 U299 ( .A1(B[30]), .A2(net26982), .B1(net34641), .B2(n216), .ZN(
        p4_adder_b[30]) );
  INV_X1 U300 ( .A(B[30]), .ZN(n216) );
  OAI22_X1 U301 ( .A1(n96), .A2(net26982), .B1(net34641), .B2(n215), .ZN(
        p4_adder_b[31]) );
  INV_X1 U302 ( .A(n96), .ZN(n215) );
  OAI22_X1 U303 ( .A1(n190), .A2(net26982), .B1(n241), .B2(net26988), .ZN(
        p4_adder_b[5]) );
  INV_X1 U304 ( .A(B[5]), .ZN(n241) );
  OAI22_X1 U305 ( .A1(B[3]), .A2(net26982), .B1(n1), .B2(n243), .ZN(
        p4_adder_b[3]) );
  INV_X1 U306 ( .A(B[3]), .ZN(n243) );
  AOI22_X1 U307 ( .A1(t2_logic_s[0]), .A2(net26996), .B1(p4_adder_s[0]), .B2(
        net26998), .ZN(n125) );
  INV_X1 U308 ( .A(n111), .ZN(RES[22]) );
  INV_X1 U309 ( .A(n105), .ZN(RES[28]) );
  INV_X1 U310 ( .A(n101), .ZN(RES[31]) );
  NAND2_X1 U311 ( .A1(n81), .A2(n82), .ZN(\t2_logic_op[2] ) );
  INV_X1 U312 ( .A(n13), .ZN(net23818) );
  CLKBUF_X1 U313 ( .A(A[2]), .Z(n205) );
  AOI222_X1 U314 ( .A1(p4_adder_s[31]), .A2(net27002), .B1(t2_shifter_s[31]), 
        .B2(net27008), .C1(t2_logic_s[31]), .C2(net26994), .ZN(n101) );
  AOI222_X1 U315 ( .A1(p4_adder_s[28]), .A2(net27000), .B1(t2_shifter_s[28]), 
        .B2(net27006), .C1(t2_logic_s[28]), .C2(net26994), .ZN(n105) );
  AOI222_X1 U316 ( .A1(p4_adder_s[22]), .A2(net27000), .B1(t2_shifter_s[22]), 
        .B2(net27006), .C1(t2_logic_s[22]), .C2(net26994), .ZN(n111) );
  CLKBUF_X1 U317 ( .A(A[0]), .Z(n204) );
  OAI22_X1 U318 ( .A1(n196), .A2(net26980), .B1(net26986), .B2(n244), .ZN(
        p4_adder_b[2]) );
  INV_X1 U319 ( .A(n189), .ZN(n244) );
  OAI22_X1 U320 ( .A1(n199), .A2(net26982), .B1(n92), .B2(n242), .ZN(
        p4_adder_b[4]) );
  INV_X1 U321 ( .A(B[4]), .ZN(n242) );
  OAI22_X1 U322 ( .A1(n195), .A2(net26980), .B1(n245), .B2(net26986), .ZN(
        p4_adder_b[1]) );
  INV_X1 U323 ( .A(n195), .ZN(n245) );
endmodule


module REG_PIPO_6_00_00_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n27), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n26), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n25), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n24), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n22), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n28), .ZN(n30) );
  INV_X1 U3 ( .A(n29), .ZN(n22) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n30), .B1(n28), .B2(DOUT[0]), .ZN(n29) );
  INV_X1 U5 ( .A(n31), .ZN(n23) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n30), .B1(n28), .B2(DOUT[1]), .ZN(n31) );
  INV_X1 U7 ( .A(n32), .ZN(n24) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n30), .B1(n28), .B2(DOUT[2]), .ZN(n32) );
  INV_X1 U9 ( .A(n33), .ZN(n25) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n30), .B1(n28), .B2(DOUT[3]), .ZN(n33) );
  INV_X1 U11 ( .A(n34), .ZN(n26) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n30), .B1(n28), .B2(DOUT[4]), .ZN(n34) );
  INV_X1 U13 ( .A(n35), .ZN(n27) );
  AOI22_X1 U14 ( .A1(DIN[5]), .A2(n30), .B1(n28), .B2(DOUT[5]), .ZN(n35) );
  INV_X1 U15 ( .A(EN), .ZN(n28) );
endmodule


module REG_PIPO_32_00000000_00000000_17 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_32_00000000_00000000_16 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n116, n131, n148, n163, net27188, net27186, net27184, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268;

  DFFR_X1 \reg_mem_reg[21]  ( .D(n258), .CK(CLK), .RN(n189), .Q(DOUT[21]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n189), .Q(DOUT[20]), 
        .QN(n148) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n250), .CK(CLK), .RN(n189), .Q(DOUT[12]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n239), .CK(CLK), .RN(n188), .Q(DOUT[0]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n240), .CK(CLK), .RN(n188), .Q(DOUT[1]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n241), .CK(CLK), .RN(n188), .Q(DOUT[2]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n242), .CK(CLK), .RN(n188), .Q(DOUT[3]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n251), .CK(CLK), .RN(n189), .Q(DOUT[13]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n247), .CK(CLK), .RN(n188), .Q(DOUT[9]), .QN(
        n223) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n246), .CK(CLK), .RN(n188), .Q(DOUT[8]), .QN(
        n222) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n243), .CK(CLK), .RN(n188), .Q(DOUT[4]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n255), .CK(CLK), .RN(n189), .Q(DOUT[17]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n253), .CK(CLK), .RN(n189), .Q(DOUT[15]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n256), .CK(CLK), .RN(n189), .Q(DOUT[18]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n249), .CK(CLK), .RN(n189), .Q(DOUT[11]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n261), .CK(CLK), .RN(n190), .Q(DOUT[24]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n257), .CK(CLK), .RN(n189), .Q(DOUT[19]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n248), .CK(CLK), .RN(n188), .Q(DOUT[10]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[31]  ( .D(n268), .CK(CLK), .RN(n190), .Q(DOUT[31]) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n252), .CK(CLK), .RN(n189), .Q(DOUT[14]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n263), .CK(CLK), .RN(n190), .Q(DOUT[26]) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n266), .CK(CLK), .RN(n190), .Q(DOUT[29]) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n262), .CK(CLK), .RN(n190), .Q(DOUT[25]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n260), .CK(CLK), .RN(n190), .Q(DOUT[23]) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n259), .CK(CLK), .RN(n190), .Q(DOUT[22]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n264), .CK(CLK), .RN(n190), .Q(DOUT[27]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n244), .CK(CLK), .RN(n188), .Q(DOUT[6]), .QN(
        n220) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n254), .CK(CLK), .RN(n189), .Q(DOUT[16]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n265), .CK(CLK), .RN(n190), .Q(DOUT[28]) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n245), .CK(CLK), .RN(n188), .Q(DOUT[7]), .QN(
        n221) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n188), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n267), .CK(CLK), .RN(RST_AN), .Q(DOUT[30]) );
  NAND2_X1 U2 ( .A1(n170), .A2(n171), .ZN(n263) );
  INV_X1 U3 ( .A(EN), .ZN(n172) );
  NAND2_X1 U4 ( .A1(n172), .A2(DOUT[26]), .ZN(n170) );
  NAND2_X1 U5 ( .A1(n183), .A2(DIN[26]), .ZN(n171) );
  NAND2_X1 U6 ( .A1(n173), .A2(n174), .ZN(n265) );
  NAND2_X1 U7 ( .A1(n172), .A2(DOUT[28]), .ZN(n174) );
  NAND2_X1 U8 ( .A1(DIN[28]), .A2(n183), .ZN(n173) );
  NAND2_X1 U9 ( .A1(n176), .A2(n175), .ZN(n266) );
  NAND2_X1 U10 ( .A1(n172), .A2(DOUT[29]), .ZN(n175) );
  NAND2_X1 U11 ( .A1(n183), .A2(DIN[29]), .ZN(n176) );
  NAND2_X1 U12 ( .A1(n177), .A2(n178), .ZN(n267) );
  NAND2_X1 U13 ( .A1(n172), .A2(DOUT[30]), .ZN(n178) );
  NAND2_X1 U14 ( .A1(n183), .A2(DIN[30]), .ZN(n177) );
  NAND2_X1 U15 ( .A1(n179), .A2(n180), .ZN(n260) );
  NAND2_X1 U16 ( .A1(n172), .A2(DOUT[23]), .ZN(n180) );
  NAND2_X1 U17 ( .A1(n183), .A2(DIN[23]), .ZN(n179) );
  NAND2_X1 U18 ( .A1(n181), .A2(n182), .ZN(n268) );
  INV_X1 U19 ( .A(net27184), .ZN(n183) );
  NAND2_X1 U20 ( .A1(n172), .A2(DOUT[31]), .ZN(n182) );
  NAND2_X1 U21 ( .A1(DIN[31]), .A2(n183), .ZN(n181) );
  OAI22_X1 U22 ( .A1(n197), .A2(n184), .B1(n227), .B2(EN), .ZN(n251) );
  OAI22_X1 U23 ( .A1(n202), .A2(n184), .B1(n230), .B2(EN), .ZN(n254) );
  OAI22_X1 U24 ( .A1(n204), .A2(n184), .B1(n234), .B2(EN), .ZN(n258) );
  OAI22_X1 U25 ( .A1(n187), .A2(n184), .B1(n148), .B2(EN), .ZN(n116) );
  OAI22_X1 U26 ( .A1(n203), .A2(n184), .B1(n235), .B2(EN), .ZN(n259) );
  OAI22_X1 U27 ( .A1(n208), .A2(n184), .B1(n215), .B2(EN), .ZN(n239) );
  OAI22_X1 U28 ( .A1(n185), .A2(n184), .B1(n163), .B2(EN), .ZN(n131) );
  BUF_X1 U29 ( .A(n184), .Z(net27186) );
  INV_X1 U30 ( .A(DIN[5]), .ZN(n185) );
  NAND2_X1 U31 ( .A1(n186), .A2(EN), .ZN(n184) );
  BUF_X1 U32 ( .A(n184), .Z(net27188) );
  BUF_X1 U33 ( .A(n184), .Z(net27184) );
  INV_X1 U34 ( .A(INIT), .ZN(n186) );
  INV_X1 U35 ( .A(DIN[20]), .ZN(n187) );
  BUF_X1 U36 ( .A(RST_AN), .Z(n188) );
  BUF_X1 U37 ( .A(RST_AN), .Z(n189) );
  BUF_X1 U38 ( .A(RST_AN), .Z(n190) );
  INV_X1 U39 ( .A(DIN[21]), .ZN(n204) );
  INV_X1 U40 ( .A(DIN[22]), .ZN(n203) );
  OAI22_X1 U41 ( .A1(n236), .A2(EN), .B1(net27184), .B2(n207), .ZN(n261) );
  INV_X1 U42 ( .A(DIN[24]), .ZN(n207) );
  OAI22_X1 U43 ( .A1(n237), .A2(EN), .B1(net27184), .B2(n206), .ZN(n262) );
  INV_X1 U44 ( .A(DIN[25]), .ZN(n206) );
  OAI22_X1 U45 ( .A1(n238), .A2(EN), .B1(net27184), .B2(n205), .ZN(n264) );
  INV_X1 U46 ( .A(DIN[27]), .ZN(n205) );
  OAI22_X1 U47 ( .A1(n216), .A2(EN), .B1(net27186), .B2(n211), .ZN(n240) );
  INV_X1 U48 ( .A(DIN[1]), .ZN(n211) );
  OAI22_X1 U49 ( .A1(n219), .A2(EN), .B1(net27186), .B2(n214), .ZN(n243) );
  INV_X1 U50 ( .A(DIN[4]), .ZN(n214) );
  OAI22_X1 U51 ( .A1(n218), .A2(EN), .B1(net27186), .B2(n210), .ZN(n242) );
  INV_X1 U52 ( .A(DIN[3]), .ZN(n210) );
  OAI22_X1 U53 ( .A1(n220), .A2(EN), .B1(net27186), .B2(n212), .ZN(n244) );
  INV_X1 U54 ( .A(DIN[6]), .ZN(n212) );
  OAI22_X1 U55 ( .A1(n221), .A2(EN), .B1(net27186), .B2(n213), .ZN(n245) );
  INV_X1 U56 ( .A(DIN[7]), .ZN(n213) );
  OAI22_X1 U57 ( .A1(n222), .A2(EN), .B1(net27186), .B2(n194), .ZN(n246) );
  INV_X1 U58 ( .A(DIN[8]), .ZN(n194) );
  OAI22_X1 U59 ( .A1(n223), .A2(EN), .B1(net27186), .B2(n193), .ZN(n247) );
  INV_X1 U60 ( .A(DIN[9]), .ZN(n193) );
  OAI22_X1 U61 ( .A1(n224), .A2(EN), .B1(net27186), .B2(n192), .ZN(n248) );
  INV_X1 U62 ( .A(DIN[10]), .ZN(n192) );
  OAI22_X1 U63 ( .A1(n225), .A2(EN), .B1(net27186), .B2(n191), .ZN(n249) );
  INV_X1 U64 ( .A(DIN[11]), .ZN(n191) );
  OAI22_X1 U65 ( .A1(n232), .A2(EN), .B1(net27188), .B2(n200), .ZN(n256) );
  INV_X1 U66 ( .A(DIN[18]), .ZN(n200) );
  OAI22_X1 U67 ( .A1(n233), .A2(EN), .B1(net27188), .B2(n199), .ZN(n257) );
  INV_X1 U68 ( .A(DIN[19]), .ZN(n199) );
  OAI22_X1 U69 ( .A1(n231), .A2(EN), .B1(net27188), .B2(n201), .ZN(n255) );
  INV_X1 U70 ( .A(DIN[17]), .ZN(n201) );
  OAI22_X1 U71 ( .A1(n226), .A2(EN), .B1(net27188), .B2(n198), .ZN(n250) );
  INV_X1 U72 ( .A(DIN[12]), .ZN(n198) );
  INV_X1 U73 ( .A(DIN[13]), .ZN(n197) );
  OAI22_X1 U74 ( .A1(n228), .A2(EN), .B1(n196), .B2(net27188), .ZN(n252) );
  INV_X1 U75 ( .A(DIN[14]), .ZN(n196) );
  OAI22_X1 U76 ( .A1(n229), .A2(EN), .B1(n195), .B2(net27188), .ZN(n253) );
  INV_X1 U77 ( .A(DIN[15]), .ZN(n195) );
  INV_X1 U78 ( .A(DIN[16]), .ZN(n202) );
  OAI22_X1 U79 ( .A1(n217), .A2(EN), .B1(n209), .B2(net27186), .ZN(n241) );
  INV_X1 U80 ( .A(DIN[2]), .ZN(n209) );
  INV_X1 U81 ( .A(DIN[0]), .ZN(n208) );
endmodule


module REG_PIPO_32_00000000_00000000_15 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U9 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U10 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U11 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U12 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U13 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U14 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U15 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U16 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U17 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U18 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U19 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U20 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U21 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U22 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U23 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U25 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U26 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U27 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U28 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U30 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U32 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U34 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U36 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U40 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U42 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U44 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U46 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U48 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U50 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_5_00_00_5 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n19), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n20), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n21), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n22), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n24), .ZN(n26) );
  INV_X1 U3 ( .A(n25), .ZN(n23) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n26), .B1(n24), .B2(DOUT[0]), .ZN(n25) );
  INV_X1 U5 ( .A(n27), .ZN(n22) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n26), .B1(n24), .B2(DOUT[1]), .ZN(n27) );
  INV_X1 U7 ( .A(n28), .ZN(n21) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n26), .B1(n24), .B2(DOUT[2]), .ZN(n28) );
  INV_X1 U9 ( .A(n29), .ZN(n20) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n26), .B1(n24), .B2(DOUT[3]), .ZN(n29) );
  INV_X1 U11 ( .A(n30), .ZN(n19) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n26), .B1(n24), .B2(DOUT[4]), .ZN(n30) );
  INV_X1 U13 ( .A(EN), .ZN(n24) );
endmodule


module REG_PIPO_1_0_0_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [0:0] DIN;
  output [0:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n3, n4, n2;

  DFFR_X1 \reg_mem_reg[0]  ( .D(n4), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]), .QN(
        n3) );
  NAND3_X1 U3 ( .A1(DIN[0]), .A2(n2), .A3(EN), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n4) );
  INV_X1 U4 ( .A(INIT), .ZN(n2) );
endmodule


module REG_PIPO_32_00000000_00000000_14 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n210), .A2(EN), .B1(n170), .B2(n207), .ZN(n242) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n207) );
  OAI22_X1 U10 ( .A1(n211), .A2(EN), .B1(n171), .B2(n206), .ZN(n243) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n206) );
  OAI22_X1 U12 ( .A1(n212), .A2(EN), .B1(n171), .B2(n205), .ZN(n244) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n205) );
  OAI22_X1 U14 ( .A1(n213), .A2(EN), .B1(n171), .B2(n204), .ZN(n245) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n204) );
  OAI22_X1 U16 ( .A1(n214), .A2(EN), .B1(n171), .B2(n203), .ZN(n246) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n203) );
  OAI22_X1 U18 ( .A1(n215), .A2(EN), .B1(n171), .B2(n202), .ZN(n247) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n202) );
  OAI22_X1 U20 ( .A1(n216), .A2(EN), .B1(n171), .B2(n201), .ZN(n248) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n201) );
  OAI22_X1 U22 ( .A1(n217), .A2(EN), .B1(n171), .B2(n200), .ZN(n249) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n200) );
  OAI22_X1 U24 ( .A1(n218), .A2(EN), .B1(n171), .B2(n199), .ZN(n250) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n199) );
  OAI22_X1 U26 ( .A1(n219), .A2(EN), .B1(n171), .B2(n198), .ZN(n251) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n198) );
  OAI22_X1 U28 ( .A1(n220), .A2(EN), .B1(n171), .B2(n197), .ZN(n252) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n197) );
  OAI22_X1 U30 ( .A1(n221), .A2(EN), .B1(n171), .B2(n196), .ZN(n253) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n196) );
  OAI22_X1 U32 ( .A1(n222), .A2(EN), .B1(n172), .B2(n195), .ZN(n254) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n195) );
  OAI22_X1 U34 ( .A1(n223), .A2(EN), .B1(n172), .B2(n194), .ZN(n255) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n194) );
  OAI22_X1 U36 ( .A1(n224), .A2(EN), .B1(n172), .B2(n193), .ZN(n256) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n193) );
  OAI22_X1 U38 ( .A1(n225), .A2(EN), .B1(n172), .B2(n192), .ZN(n257) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n192) );
  OAI22_X1 U40 ( .A1(n226), .A2(EN), .B1(n172), .B2(n191), .ZN(n258) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n191) );
  OAI22_X1 U42 ( .A1(n227), .A2(EN), .B1(n172), .B2(n190), .ZN(n259) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n190) );
  OAI22_X1 U44 ( .A1(n228), .A2(EN), .B1(n172), .B2(n189), .ZN(n260) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n189) );
  OAI22_X1 U46 ( .A1(n229), .A2(EN), .B1(n172), .B2(n188), .ZN(n261) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n188) );
  OAI22_X1 U48 ( .A1(n230), .A2(EN), .B1(n172), .B2(n187), .ZN(n262) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n187) );
  OAI22_X1 U50 ( .A1(n231), .A2(EN), .B1(n172), .B2(n186), .ZN(n263) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n186) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n185), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n185) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n184), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n184) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n183), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n183) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n182), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n182) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n181), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n181) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n180), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n180) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n179), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n179) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n178), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n178) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n177), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n177) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n176), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n176) );
  NAND2_X1 U72 ( .A1(n208), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n208) );
endmodule


module REG_PIPO_32_00000000_00000000_13 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n210), .A2(EN), .B1(n170), .B2(n207), .ZN(n242) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n207) );
  OAI22_X1 U10 ( .A1(n211), .A2(EN), .B1(n171), .B2(n206), .ZN(n243) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n206) );
  OAI22_X1 U12 ( .A1(n212), .A2(EN), .B1(n171), .B2(n205), .ZN(n244) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n205) );
  OAI22_X1 U14 ( .A1(n213), .A2(EN), .B1(n171), .B2(n204), .ZN(n245) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n204) );
  OAI22_X1 U16 ( .A1(n214), .A2(EN), .B1(n171), .B2(n203), .ZN(n246) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n203) );
  OAI22_X1 U18 ( .A1(n215), .A2(EN), .B1(n171), .B2(n202), .ZN(n247) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n202) );
  OAI22_X1 U20 ( .A1(n216), .A2(EN), .B1(n171), .B2(n201), .ZN(n248) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n201) );
  OAI22_X1 U22 ( .A1(n217), .A2(EN), .B1(n171), .B2(n200), .ZN(n249) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n200) );
  OAI22_X1 U24 ( .A1(n218), .A2(EN), .B1(n171), .B2(n199), .ZN(n250) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n199) );
  OAI22_X1 U26 ( .A1(n219), .A2(EN), .B1(n171), .B2(n198), .ZN(n251) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n198) );
  OAI22_X1 U28 ( .A1(n220), .A2(EN), .B1(n171), .B2(n197), .ZN(n252) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n197) );
  OAI22_X1 U30 ( .A1(n221), .A2(EN), .B1(n171), .B2(n196), .ZN(n253) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n196) );
  OAI22_X1 U32 ( .A1(n222), .A2(EN), .B1(n172), .B2(n195), .ZN(n254) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n195) );
  OAI22_X1 U34 ( .A1(n223), .A2(EN), .B1(n172), .B2(n194), .ZN(n255) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n194) );
  OAI22_X1 U36 ( .A1(n224), .A2(EN), .B1(n172), .B2(n193), .ZN(n256) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n193) );
  OAI22_X1 U38 ( .A1(n225), .A2(EN), .B1(n172), .B2(n192), .ZN(n257) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n192) );
  OAI22_X1 U40 ( .A1(n226), .A2(EN), .B1(n172), .B2(n191), .ZN(n258) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n191) );
  OAI22_X1 U42 ( .A1(n227), .A2(EN), .B1(n172), .B2(n190), .ZN(n259) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n190) );
  OAI22_X1 U44 ( .A1(n228), .A2(EN), .B1(n172), .B2(n189), .ZN(n260) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n189) );
  OAI22_X1 U46 ( .A1(n229), .A2(EN), .B1(n172), .B2(n188), .ZN(n261) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n188) );
  OAI22_X1 U48 ( .A1(n230), .A2(EN), .B1(n172), .B2(n187), .ZN(n262) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n187) );
  OAI22_X1 U50 ( .A1(n231), .A2(EN), .B1(n172), .B2(n186), .ZN(n263) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n186) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n185), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n185) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n184), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n184) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n183), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n183) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n182), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n182) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n181), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n181) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n180), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n180) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n179), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n179) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n178), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n178) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n177), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n177) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n176), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n176) );
  NAND2_X1 U72 ( .A1(n208), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n208) );
endmodule


module REG_PIPO_32_00000000_00000000_12 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n273), .CK(CLK), .RN(n175), .Q(DOUT[31]), 
        .QN(n241) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n272), .CK(CLK), .RN(n175), .Q(DOUT[30]), 
        .QN(n240) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n271), .CK(CLK), .RN(n175), .Q(DOUT[29]), 
        .QN(n239) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n270), .CK(CLK), .RN(n175), .Q(DOUT[28]), 
        .QN(n238) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n269), .CK(CLK), .RN(n175), .Q(DOUT[27]), 
        .QN(n237) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n268), .CK(CLK), .RN(n175), .Q(DOUT[26]), 
        .QN(n236) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n267), .CK(CLK), .RN(n175), .Q(DOUT[25]), 
        .QN(n235) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n266), .CK(CLK), .RN(n175), .Q(DOUT[24]), 
        .QN(n234) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n265), .CK(CLK), .RN(n175), .Q(DOUT[23]), 
        .QN(n233) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n264), .CK(CLK), .RN(n175), .Q(DOUT[22]), 
        .QN(n232) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n263), .CK(CLK), .RN(n174), .Q(DOUT[21]), 
        .QN(n231) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n262), .CK(CLK), .RN(n174), .Q(DOUT[20]), 
        .QN(n230) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n261), .CK(CLK), .RN(n174), .Q(DOUT[19]), 
        .QN(n229) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n260), .CK(CLK), .RN(n174), .Q(DOUT[18]), 
        .QN(n228) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n259), .CK(CLK), .RN(n174), .Q(DOUT[17]), 
        .QN(n227) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n258), .CK(CLK), .RN(n174), .Q(DOUT[16]), 
        .QN(n226) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n257), .CK(CLK), .RN(n174), .Q(DOUT[15]), 
        .QN(n225) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n256), .CK(CLK), .RN(n174), .Q(DOUT[14]), 
        .QN(n224) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n255), .CK(CLK), .RN(n174), .Q(DOUT[13]), 
        .QN(n223) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n254), .CK(CLK), .RN(n174), .Q(DOUT[12]), 
        .QN(n222) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n253), .CK(CLK), .RN(n174), .Q(DOUT[11]), 
        .QN(n221) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n252), .CK(CLK), .RN(n173), .Q(DOUT[10]), 
        .QN(n220) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n251), .CK(CLK), .RN(n173), .Q(DOUT[9]), .QN(
        n219) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n250), .CK(CLK), .RN(n173), .Q(DOUT[8]), .QN(
        n218) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n249), .CK(CLK), .RN(n173), .Q(DOUT[7]), .QN(
        n217) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n248), .CK(CLK), .RN(n173), .Q(DOUT[6]), .QN(
        n216) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n247), .CK(CLK), .RN(n173), .Q(DOUT[5]), .QN(
        n215) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n246), .CK(CLK), .RN(n173), .Q(DOUT[4]), .QN(
        n214) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n245), .CK(CLK), .RN(n173), .Q(DOUT[3]), .QN(
        n213) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n244), .CK(CLK), .RN(n173), .Q(DOUT[2]), .QN(
        n212) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n243), .CK(CLK), .RN(n173), .Q(DOUT[1]), .QN(
        n211) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n242), .CK(CLK), .RN(n173), .Q(DOUT[0]), .QN(
        n210) );
  BUF_X1 U2 ( .A(n209), .Z(n172) );
  BUF_X1 U3 ( .A(n209), .Z(n171) );
  BUF_X1 U4 ( .A(n209), .Z(n170) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n173) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n174) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n175) );
  OAI22_X1 U8 ( .A1(n210), .A2(EN), .B1(n170), .B2(n208), .ZN(n242) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n208) );
  OAI22_X1 U10 ( .A1(n211), .A2(EN), .B1(n171), .B2(n207), .ZN(n243) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n207) );
  OAI22_X1 U12 ( .A1(n212), .A2(EN), .B1(n171), .B2(n206), .ZN(n244) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n206) );
  OAI22_X1 U14 ( .A1(n213), .A2(EN), .B1(n171), .B2(n205), .ZN(n245) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n205) );
  OAI22_X1 U16 ( .A1(n214), .A2(EN), .B1(n171), .B2(n204), .ZN(n246) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n204) );
  OAI22_X1 U18 ( .A1(n215), .A2(EN), .B1(n171), .B2(n203), .ZN(n247) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n203) );
  OAI22_X1 U20 ( .A1(n216), .A2(EN), .B1(n171), .B2(n202), .ZN(n248) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n202) );
  OAI22_X1 U22 ( .A1(n217), .A2(EN), .B1(n171), .B2(n201), .ZN(n249) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n201) );
  OAI22_X1 U24 ( .A1(n218), .A2(EN), .B1(n171), .B2(n200), .ZN(n250) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n200) );
  OAI22_X1 U26 ( .A1(n219), .A2(EN), .B1(n171), .B2(n199), .ZN(n251) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n199) );
  OAI22_X1 U28 ( .A1(n220), .A2(EN), .B1(n171), .B2(n198), .ZN(n252) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n198) );
  OAI22_X1 U30 ( .A1(n221), .A2(EN), .B1(n171), .B2(n197), .ZN(n253) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n197) );
  OAI22_X1 U32 ( .A1(n222), .A2(EN), .B1(n172), .B2(n196), .ZN(n254) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n196) );
  OAI22_X1 U34 ( .A1(n223), .A2(EN), .B1(n172), .B2(n195), .ZN(n255) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n195) );
  OAI22_X1 U36 ( .A1(n224), .A2(EN), .B1(n172), .B2(n194), .ZN(n256) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n194) );
  OAI22_X1 U38 ( .A1(n225), .A2(EN), .B1(n172), .B2(n193), .ZN(n257) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n193) );
  OAI22_X1 U40 ( .A1(n226), .A2(EN), .B1(n172), .B2(n192), .ZN(n258) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n192) );
  OAI22_X1 U42 ( .A1(n227), .A2(EN), .B1(n172), .B2(n191), .ZN(n259) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n191) );
  OAI22_X1 U44 ( .A1(n228), .A2(EN), .B1(n172), .B2(n190), .ZN(n260) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n190) );
  OAI22_X1 U46 ( .A1(n229), .A2(EN), .B1(n172), .B2(n189), .ZN(n261) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n189) );
  OAI22_X1 U48 ( .A1(n230), .A2(EN), .B1(n172), .B2(n188), .ZN(n262) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n188) );
  OAI22_X1 U50 ( .A1(n231), .A2(EN), .B1(n172), .B2(n187), .ZN(n263) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n187) );
  OAI22_X1 U52 ( .A1(n232), .A2(EN), .B1(n170), .B2(n186), .ZN(n264) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n186) );
  OAI22_X1 U54 ( .A1(n233), .A2(EN), .B1(n170), .B2(n185), .ZN(n265) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n185) );
  OAI22_X1 U56 ( .A1(n234), .A2(EN), .B1(n170), .B2(n184), .ZN(n266) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n184) );
  OAI22_X1 U58 ( .A1(n235), .A2(EN), .B1(n170), .B2(n183), .ZN(n267) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n183) );
  OAI22_X1 U60 ( .A1(n236), .A2(EN), .B1(n170), .B2(n182), .ZN(n268) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n182) );
  OAI22_X1 U62 ( .A1(n237), .A2(EN), .B1(n170), .B2(n181), .ZN(n269) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n181) );
  OAI22_X1 U64 ( .A1(n238), .A2(EN), .B1(n170), .B2(n180), .ZN(n270) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n180) );
  OAI22_X1 U66 ( .A1(n239), .A2(EN), .B1(n170), .B2(n179), .ZN(n271) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n179) );
  OAI22_X1 U68 ( .A1(n240), .A2(EN), .B1(n170), .B2(n178), .ZN(n272) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n178) );
  OAI22_X1 U70 ( .A1(n241), .A2(EN), .B1(n170), .B2(n177), .ZN(n273) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n177) );
  NAND2_X1 U72 ( .A1(n176), .A2(EN), .ZN(n209) );
  INV_X1 U73 ( .A(INIT), .ZN(n176) );
endmodule


module REG_PIPO_5_00_00_4 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n19), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n20), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n21), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n22), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  INV_X1 U2 ( .A(n25), .ZN(n23) );
  AOI22_X1 U3 ( .A1(DIN[0]), .A2(n26), .B1(n24), .B2(DOUT[0]), .ZN(n25) );
  INV_X1 U4 ( .A(n27), .ZN(n22) );
  AOI22_X1 U5 ( .A1(DIN[1]), .A2(n26), .B1(n24), .B2(DOUT[1]), .ZN(n27) );
  INV_X1 U6 ( .A(n28), .ZN(n21) );
  AOI22_X1 U7 ( .A1(DIN[2]), .A2(n26), .B1(n24), .B2(DOUT[2]), .ZN(n28) );
  INV_X1 U8 ( .A(n29), .ZN(n20) );
  AOI22_X1 U9 ( .A1(DIN[3]), .A2(n26), .B1(n24), .B2(DOUT[3]), .ZN(n29) );
  INV_X1 U10 ( .A(n30), .ZN(n19) );
  AOI22_X1 U11 ( .A1(DIN[4]), .A2(n26), .B1(n24), .B2(DOUT[4]), .ZN(n30) );
  INV_X1 U12 ( .A(EN), .ZN(n24) );
  NOR2_X1 U13 ( .A1(INIT), .A2(n24), .ZN(n26) );
endmodule


module DATAPATH_1_DW01_add_2 ( A, B, CI, SUM, CO );
  input [30:0] A;
  input [30:0] B;
  output [30:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X1 U2 ( .A1(n1), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n34), .A2(n35), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n32), .A2(n33), .ZN(n2) );
  XOR2_X1 U5 ( .A(A[11]), .B(n3), .Z(SUM[11]) );
  NOR2_X1 U6 ( .A1(n7), .A2(n44), .ZN(n3) );
  XNOR2_X1 U7 ( .A(n4), .B(A[23]), .ZN(SUM[23]) );
  NAND2_X1 U8 ( .A1(A[22]), .A2(n11), .ZN(n4) );
  XNOR2_X1 U9 ( .A(n5), .B(A[27]), .ZN(SUM[27]) );
  NAND2_X1 U10 ( .A1(A[26]), .A2(n10), .ZN(n5) );
  XNOR2_X1 U11 ( .A(n6), .B(A[30]), .ZN(SUM[30]) );
  NAND2_X1 U12 ( .A1(n12), .A2(A[29]), .ZN(n6) );
  XOR2_X1 U13 ( .A(n13), .B(n48), .Z(SUM[9]) );
  XOR2_X1 U14 ( .A(n7), .B(n44), .Z(SUM[10]) );
  NOR2_X1 U15 ( .A1(n46), .A2(n38), .ZN(n14) );
  NOR2_X1 U16 ( .A1(n43), .A2(n35), .ZN(n42) );
  OR2_X1 U17 ( .A1(n48), .A2(n13), .ZN(n7) );
  INV_X1 U18 ( .A(n20), .ZN(n22) );
  INV_X1 U19 ( .A(n24), .ZN(n26) );
  INV_X1 U20 ( .A(n28), .ZN(n31) );
  NAND2_X1 U21 ( .A1(n36), .A2(n37), .ZN(n34) );
  XOR2_X1 U22 ( .A(A[5]), .B(n17), .Z(SUM[5]) );
  XOR2_X1 U23 ( .A(A[13]), .B(n41), .Z(SUM[13]) );
  XOR2_X1 U24 ( .A(A[8]), .B(n14), .Z(SUM[8]) );
  AND2_X1 U25 ( .A1(n41), .A2(A[13]), .ZN(n40) );
  AND2_X1 U26 ( .A1(n17), .A2(A[5]), .ZN(n16) );
  XOR2_X1 U27 ( .A(A[20]), .B(n27), .Z(SUM[20]) );
  NOR2_X1 U28 ( .A1(n24), .A2(n25), .ZN(n23) );
  NAND4_X1 U29 ( .A1(A[11]), .A2(A[10]), .A3(A[9]), .A4(A[8]), .ZN(n35) );
  NOR2_X1 U30 ( .A1(n28), .A2(n29), .ZN(n27) );
  NOR2_X1 U31 ( .A1(n20), .A2(n21), .ZN(n19) );
  XNOR2_X1 U32 ( .A(n39), .B(A[15]), .ZN(SUM[15]) );
  NAND2_X1 U33 ( .A1(n40), .A2(A[14]), .ZN(n39) );
  XNOR2_X1 U34 ( .A(A[3]), .B(SUM[2]), .ZN(SUM[3]) );
  XNOR2_X1 U35 ( .A(n15), .B(A[7]), .ZN(SUM[7]) );
  NAND2_X1 U36 ( .A1(n16), .A2(A[6]), .ZN(n15) );
  XNOR2_X1 U37 ( .A(n30), .B(A[19]), .ZN(SUM[19]) );
  NAND2_X1 U38 ( .A1(n9), .A2(A[18]), .ZN(n30) );
  XOR2_X1 U39 ( .A(A[6]), .B(n16), .Z(SUM[6]) );
  XOR2_X1 U40 ( .A(A[12]), .B(n42), .Z(SUM[12]) );
  XOR2_X1 U41 ( .A(A[14]), .B(n40), .Z(SUM[14]) );
  XOR2_X1 U42 ( .A(A[16]), .B(n8), .Z(SUM[16]) );
  XOR2_X1 U43 ( .A(A[17]), .B(n31), .Z(SUM[17]) );
  XOR2_X1 U44 ( .A(A[4]), .B(n37), .Z(SUM[4]) );
  XOR2_X1 U45 ( .A(A[18]), .B(n9), .Z(SUM[18]) );
  NAND4_X1 U46 ( .A1(A[4]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n38) );
  AND2_X1 U47 ( .A1(A[12]), .A2(n42), .ZN(n41) );
  NOR2_X1 U48 ( .A1(n45), .A2(n46), .ZN(n17) );
  XOR2_X1 U49 ( .A(A[21]), .B(n26), .Z(SUM[21]) );
  XOR2_X1 U50 ( .A(A[25]), .B(n22), .Z(SUM[25]) );
  XOR2_X1 U51 ( .A(n10), .B(A[26]), .Z(SUM[26]) );
  XOR2_X1 U52 ( .A(n12), .B(A[29]), .Z(SUM[29]) );
  XOR2_X1 U53 ( .A(n11), .B(A[22]), .Z(SUM[22]) );
  XOR2_X1 U54 ( .A(n23), .B(A[24]), .Z(SUM[24]) );
  XOR2_X1 U55 ( .A(n19), .B(A[28]), .Z(SUM[28]) );
  NAND2_X1 U56 ( .A1(n8), .A2(A[16]), .ZN(n28) );
  NAND2_X1 U57 ( .A1(n27), .A2(A[20]), .ZN(n24) );
  NAND2_X1 U58 ( .A1(n23), .A2(A[24]), .ZN(n20) );
  NAND2_X1 U59 ( .A1(n14), .A2(A[8]), .ZN(n13) );
  AND2_X1 U60 ( .A1(A[17]), .A2(n31), .ZN(n9) );
  AND2_X1 U61 ( .A1(A[25]), .A2(n22), .ZN(n10) );
  AND2_X1 U62 ( .A1(A[21]), .A2(n26), .ZN(n11) );
  AND2_X1 U63 ( .A1(n19), .A2(A[28]), .ZN(n12) );
  NOR2_X1 U64 ( .A1(SUM[2]), .A2(n47), .ZN(n37) );
  NAND2_X1 U65 ( .A1(A[12]), .A2(A[13]), .ZN(n33) );
  NAND2_X1 U66 ( .A1(A[14]), .A2(A[15]), .ZN(n32) );
  INV_X1 U67 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U68 ( .A(A[4]), .ZN(n45) );
  INV_X1 U69 ( .A(A[9]), .ZN(n48) );
  INV_X1 U70 ( .A(A[3]), .ZN(n47) );
  NAND3_X1 U71 ( .A1(A[26]), .A2(A[27]), .A3(A[25]), .ZN(n21) );
  NAND3_X1 U72 ( .A1(A[22]), .A2(A[23]), .A3(A[21]), .ZN(n25) );
  NAND3_X1 U73 ( .A1(A[18]), .A2(A[19]), .A3(A[17]), .ZN(n29) );
  INV_X1 U74 ( .A(n38), .ZN(n36) );
  INV_X1 U75 ( .A(n14), .ZN(n43) );
  INV_X1 U76 ( .A(A[10]), .ZN(n44) );
  INV_X1 U77 ( .A(n37), .ZN(n46) );
endmodule


module DATAPATH_1 ( CLK, RST_AN, .CTRL_WORD({\CTRL_WORD[J_TYPE_IMM_SEL] , 
        \CTRL_WORD[R_TYPE_SEL] , \CTRL_WORD[IMM_SEL] , 
        \CTRL_WORD[PC_PLS_4_SEL] , \CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] , \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }), INSTR_CU, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .DP_SIG({
        \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] , 
        \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] , 
        \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] , 
        \DP_SIG[INSTR_OPCODE_M][0] }), IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] INSTR_CU;
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN, \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] , \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  wire   \npc_f[31] , n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n184, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n246, n247, n248, n249, n250, n251, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, net23121, net23132, net23138, net23147,
         net25878, net25874, net25872, net25868, net25862, net25860, net25888,
         net27502, net33900, net34379, net34378, net34429, net34728, net34727,
         net34734, net34744, net40517, net40540, n245, n1, n2, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n183, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n252, n303, n304, n305, n306, n307,
         n308, n309;
  wire   [30:0] pc_pls_4_f;
  wire   [31:0] pc_pls_4_d;
  wire   [31:0] instr_d;
  wire   [4:0] rf_waddr_d;
  wire   [31:0] rf_dout1_d;
  wire   [31:0] rf_dout2_d;
  wire   [4:0] rf_waddr_wb;
  wire   [31:16] imm_d;
  wire   [5:0] instr_opcode_e;
  wire   [31:0] pc_pls_4_e;
  wire   [31:0] rf_dout1_e;
  wire   [31:0] rf_dout2_e;
  wire   [31:0] imm_e;
  wire   [4:0] rs2_e;
  wire   [4:0] rs3_e;
  wire   [31:0] alu_a_e;
  wire   [31:0] alu_out_e;
  wire   [31:0] pc_pls_4_m;
  wire   [4:0] rf_waddr_m;
  wire   [31:0] pc_pls_4_wb;
  wire   [31:0] alu_out_wb;
  wire   [31:0] dmem_dout_wb;
  assign INSTR_CU[31] = IMEM_DOUT[31];
  assign INSTR_CU[30] = IMEM_DOUT[30];
  assign INSTR_CU[29] = IMEM_DOUT[29];
  assign INSTR_CU[28] = IMEM_DOUT[28];
  assign INSTR_CU[27] = IMEM_DOUT[27];
  assign INSTR_CU[26] = IMEM_DOUT[26];
  assign INSTR_CU[25] = IMEM_DOUT[25];
  assign INSTR_CU[24] = IMEM_DOUT[24];
  assign INSTR_CU[23] = IMEM_DOUT[23];
  assign INSTR_CU[22] = IMEM_DOUT[22];
  assign INSTR_CU[21] = IMEM_DOUT[21];
  assign INSTR_CU[20] = IMEM_DOUT[20];
  assign INSTR_CU[19] = IMEM_DOUT[19];
  assign INSTR_CU[18] = IMEM_DOUT[18];
  assign INSTR_CU[17] = IMEM_DOUT[17];
  assign INSTR_CU[16] = IMEM_DOUT[16];
  assign INSTR_CU[15] = IMEM_DOUT[15];
  assign INSTR_CU[14] = IMEM_DOUT[14];
  assign INSTR_CU[13] = IMEM_DOUT[13];
  assign INSTR_CU[12] = IMEM_DOUT[12];
  assign INSTR_CU[11] = IMEM_DOUT[11];
  assign INSTR_CU[10] = IMEM_DOUT[10];
  assign INSTR_CU[9] = IMEM_DOUT[9];
  assign INSTR_CU[8] = IMEM_DOUT[8];
  assign INSTR_CU[7] = IMEM_DOUT[7];
  assign INSTR_CU[6] = IMEM_DOUT[6];
  assign INSTR_CU[5] = IMEM_DOUT[5];
  assign INSTR_CU[4] = IMEM_DOUT[4];
  assign INSTR_CU[3] = IMEM_DOUT[3];
  assign INSTR_CU[2] = IMEM_DOUT[2];
  assign INSTR_CU[1] = IMEM_DOUT[1];
  assign INSTR_CU[0] = IMEM_DOUT[0];

  OAI21_X2 U192 ( .B1(n34), .B2(n102), .A(n291), .ZN(alu_a_e[19]) );
  OAI21_X2 U200 ( .B1(n23), .B2(n106), .A(n295), .ZN(alu_a_e[15]) );
  REG_PIPO_32_fffffffc_fffffffc_1 U_PC_REG ( .CLK(CLK), .RST_AN(n52), .EN(1'b1), .INIT(1'b0), .DIN({\npc_f[31] , n55, n56, n57, n58, n59, n60, n61, n62, n63, 
        n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
        n78, n79, n80, n81, n82, n83, n84, n189}), .DOUT(IMEM_ADDR) );
  REG_PIPO_32_00000000_00000000_23 U_PC_PLS_4_REG_FD ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN({1'b0, pc_pls_4_f}), 
        .DOUT(pc_pls_4_d) );
  REG_PIPO_32_00000000_00000000_22 U_INSTR_REG_FD ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN(IMEM_DOUT), .DOUT(instr_d) );
  RF_ADDR_W5_DATA_W32_1 U_RF ( .CLK(CLK), .RST_AN(n51), .ENABLE(1'b1), .RD1(
        1'b1), .RD2(1'b1), .WR(\CTRL_WORD[RF_WEN] ), .ADD_WR(rf_waddr_d), 
        .ADD_RD1(instr_d[25:21]), .ADD_RD2(instr_d[20:16]), .DATAIN({n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216, n252, n303, n304, n305, n306}), .OUT1(rf_dout1_d), .OUT2(
        rf_dout2_d) );
  REG_PIPO_6_00_00_3 U_INSTR_OPCODE_REG_DE ( .CLK(CLK), .RST_AN(n51), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[31:26]), .DOUT(instr_opcode_e) );
  REG_PIPO_32_00000000_00000000_21 U_PC_PLS_4_REG_DE ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(pc_pls_4_d), .DOUT(
        pc_pls_4_e) );
  REG_PIPO_32_00000000_00000000_20 U_RF_DOUT1_REG_DE ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout1_d), .DOUT(
        rf_dout1_e) );
  REG_PIPO_32_00000000_00000000_19 U_RF_DOUT2_REG_DE ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout2_d), .DOUT(
        rf_dout2_e) );
  REG_PIPO_32_00000000_00000000_18 U_IMM_REG_DE ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN({imm_d[31], imm_d[31], 
        imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[24:16], 
        instr_d[15:0]}), .DOUT(imm_e) );
  REG_PIPO_5_00_00_7 U_RS2_REG_DE ( .CLK(CLK), .RST_AN(n51), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[20:16]), .DOUT(rs2_e) );
  REG_PIPO_5_00_00_6 U_RS3_REG_DE ( .CLK(CLK), .RST_AN(n51), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[15:11]), .DOUT(rs3_e) );
  ALU_DATA_W32_1 U_ALU ( .FUNC({\CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] }), .A({alu_a_e[31:25], n20, alu_a_e[23], n6, 
        alu_a_e[21], n21, alu_a_e[19:18], n2, alu_a_e[16:13], n30, 
        alu_a_e[11:9], n18, alu_a_e[7:0]}), .B({net23147, n122, n123, n124, 
        n125, n126, n22, n127, n128, net23138, n129, n130, n131, n132, n133, 
        net23132, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
        net23121, n183, n185, n186, n187, n188}), .RES(alu_out_e) );
  REG_PIPO_6_00_00_2 U_INSTR_OPCODE_REG_EM ( .CLK(CLK), .RST_AN(n51), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(instr_opcode_e), .DOUT({
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }) );
  REG_PIPO_32_00000000_00000000_17 U_PC_PLS_4_REG_EM ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(pc_pls_4_e), .DOUT(
        pc_pls_4_m) );
  REG_PIPO_32_00000000_00000000_16 U_ALU_OUT_REG_EM ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(alu_out_e), .DOUT(
        DMEM_RWADDR) );
  REG_PIPO_32_00000000_00000000_15 U_DMEM_DOUT_REG_EM ( .CLK(CLK), .RST_AN(n52), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(rf_dout2_e), .DOUT(DMEM_DIN) );
  REG_PIPO_5_00_00_5 U_RF_WADDR_REG_EM ( .CLK(CLK), .RST_AN(n51), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN({n85, n86, n87, n88, n89}), .DOUT(
        rf_waddr_m) );
  REG_PIPO_1_0_0_1 U_IS_0_REG_EM ( .CLK(CLK), .RST_AN(n52), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_EM] ), .DIN(n302), .DOUT(\DP_SIG[CMPR_0_IS_0_M] ) );
  REG_PIPO_32_00000000_00000000_14 U_PC_PLS_4_REG_MWB ( .CLK(CLK), .RST_AN(n52), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(pc_pls_4_m), .DOUT(pc_pls_4_wb) );
  REG_PIPO_32_00000000_00000000_13 U_ALU_OUT_REG_MWB ( .CLK(CLK), .RST_AN(n52), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_RWADDR), .DOUT(
        alu_out_wb) );
  REG_PIPO_32_00000000_00000000_12 U_DMEM_DOUT_REG_MWB ( .CLK(CLK), .RST_AN(
        n52), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_DOUT), .DOUT(
        dmem_dout_wb) );
  REG_PIPO_5_00_00_4 U_RF_WADDR_REG_MWB ( .CLK(CLK), .RST_AN(n51), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(rf_waddr_m), .DOUT(rf_waddr_wb) );
  DATAPATH_1_DW01_add_2 add_242 ( .A(IMEM_ADDR[30:0]), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_pls_4_f) );
  CLKBUF_X3 U5 ( .A(alu_a_e[8]), .Z(n18) );
  BUF_X1 U7 ( .A(n8), .Z(net40540) );
  BUF_X2 U8 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n49) );
  OAI21_X1 U9 ( .B1(n33), .B2(n120), .A(n290), .ZN(alu_a_e[1]) );
  INV_X1 U10 ( .A(n257), .ZN(n130) );
  INV_X1 U11 ( .A(n250), .ZN(n125) );
  BUF_X2 U12 ( .A(alu_a_e[22]), .Z(n6) );
  BUF_X1 U13 ( .A(alu_a_e[24]), .Z(n20) );
  OAI21_X1 U14 ( .B1(n50), .B2(n110), .A(n299), .ZN(alu_a_e[11]) );
  BUF_X2 U15 ( .A(alu_a_e[17]), .Z(n2) );
  BUF_X1 U16 ( .A(alu_a_e[20]), .Z(n21) );
  BUF_X1 U17 ( .A(n49), .Z(n33) );
  BUF_X2 U18 ( .A(n17), .Z(n16) );
  BUF_X1 U19 ( .A(n15), .Z(n1) );
  BUF_X1 U20 ( .A(n17), .Z(net27502) );
  CLKBUF_X1 U21 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n11) );
  OAI21_X2 U22 ( .B1(n36), .B2(n98), .A(n286), .ZN(alu_a_e[23]) );
  OAI21_X2 U23 ( .B1(n33), .B2(n91), .A(n278), .ZN(alu_a_e[30]) );
  BUF_X1 U24 ( .A(n8), .Z(n7) );
  INV_X1 U25 ( .A(\CTRL_WORD[IMM_SEL] ), .ZN(n8) );
  INV_X1 U26 ( .A(n8), .ZN(n9) );
  CLKBUF_X1 U27 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n10) );
  CLKBUF_X1 U28 ( .A(n10), .Z(net25868) );
  CLKBUF_X1 U29 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net25874) );
  BUF_X1 U30 ( .A(net34429), .Z(n12) );
  INV_X1 U31 ( .A(net25888), .ZN(n13) );
  INV_X1 U32 ( .A(net25874), .ZN(n14) );
  CLKBUF_X1 U33 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net25888) );
  BUF_X1 U34 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n15) );
  BUF_X1 U35 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net34429) );
  AOI22_X1 U36 ( .A1(rf_dout2_e[31]), .A2(n16), .B1(net34378), .B2(imm_e[31]), 
        .ZN(n245) );
  INV_X1 U37 ( .A(n245), .ZN(net23147) );
  AOI22_X1 U38 ( .A1(rf_dout2_e[22]), .A2(n7), .B1(imm_e[22]), .B2(net40517), 
        .ZN(n255) );
  AOI22_X1 U39 ( .A1(n7), .A2(rf_dout2_e[5]), .B1(net34728), .B2(imm_e[5]), 
        .ZN(n242) );
  AOI22_X1 U40 ( .A1(rf_dout2_e[16]), .A2(net33900), .B1(n9), .B2(imm_e[16]), 
        .ZN(n262) );
  INV_X1 U41 ( .A(\CTRL_WORD[IMM_SEL] ), .ZN(n17) );
  OAI21_X1 U42 ( .B1(n50), .B2(n113), .A(n271), .ZN(alu_a_e[8]) );
  BUF_X1 U43 ( .A(n35), .Z(n31) );
  BUF_X1 U44 ( .A(net25878), .Z(net34727) );
  BUF_X2 U45 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n29) );
  CLKBUF_X1 U46 ( .A(n10), .Z(net40517) );
  BUF_X1 U47 ( .A(n10), .Z(net25872) );
  CLKBUF_X1 U48 ( .A(n49), .Z(n19) );
  BUF_X1 U49 ( .A(net25878), .Z(net34378) );
  CLKBUF_X3 U50 ( .A(n35), .Z(n36) );
  OAI21_X1 U51 ( .B1(n23), .B2(n114), .A(n272), .ZN(alu_a_e[7]) );
  BUF_X2 U52 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n35) );
  OAI21_X1 U53 ( .B1(n24), .B2(n97), .A(n285), .ZN(alu_a_e[24]) );
  OAI21_X1 U54 ( .B1(n34), .B2(n101), .A(n289), .ZN(alu_a_e[20]) );
  OAI21_X2 U55 ( .B1(n50), .B2(n116), .A(n274), .ZN(alu_a_e[5]) );
  NAND2_X1 U56 ( .A1(n25), .A2(n283), .ZN(alu_a_e[26]) );
  INV_X1 U57 ( .A(net34429), .ZN(net34744) );
  BUF_X1 U58 ( .A(net34429), .Z(net34734) );
  BUF_X1 U59 ( .A(net25878), .Z(net34728) );
  BUF_X1 U60 ( .A(n15), .Z(net34379) );
  INV_X1 U61 ( .A(n240), .ZN(n142) );
  BUF_X1 U62 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net25878) );
  NAND2_X1 U63 ( .A1(n26), .A2(n27), .ZN(n22) );
  BUF_X1 U64 ( .A(n35), .Z(n23) );
  BUF_X1 U65 ( .A(n35), .Z(n24) );
  OR2_X1 U66 ( .A1(n28), .A2(n95), .ZN(n25) );
  OAI21_X1 U67 ( .B1(n24), .B2(n100), .A(n288), .ZN(alu_a_e[21]) );
  OAI21_X1 U68 ( .B1(n28), .B2(n105), .A(n294), .ZN(alu_a_e[16]) );
  INV_X1 U69 ( .A(n259), .ZN(n131) );
  INV_X1 U70 ( .A(n265), .ZN(n136) );
  NAND2_X1 U71 ( .A1(rf_dout2_e[25]), .A2(net34744), .ZN(n26) );
  NAND2_X1 U72 ( .A1(imm_e[25]), .A2(n12), .ZN(n27) );
  INV_X1 U73 ( .A(n239), .ZN(n141) );
  OAI21_X1 U74 ( .B1(n24), .B2(n94), .A(n282), .ZN(alu_a_e[27]) );
  BUF_X1 U75 ( .A(n35), .Z(n28) );
  OAI21_X1 U76 ( .B1(n23), .B2(n112), .A(n270), .ZN(alu_a_e[9]) );
  OAI21_X1 U77 ( .B1(n28), .B2(n92), .A(n280), .ZN(alu_a_e[29]) );
  INV_X1 U78 ( .A(n244), .ZN(n185) );
  BUF_X2 U79 ( .A(alu_a_e[12]), .Z(n30) );
  OAI21_X1 U80 ( .B1(n28), .B2(n109), .A(n298), .ZN(alu_a_e[12]) );
  INV_X1 U81 ( .A(n11), .ZN(net33900) );
  INV_X1 U82 ( .A(n258), .ZN(n187) );
  INV_X1 U83 ( .A(n241), .ZN(n143) );
  INV_X1 U84 ( .A(n242), .ZN(net23121) );
  BUF_X1 U85 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n50) );
  OAI21_X1 U86 ( .B1(n29), .B2(n104), .A(n293), .ZN(alu_a_e[17]) );
  OAI21_X1 U87 ( .B1(n29), .B2(n99), .A(n287), .ZN(alu_a_e[22]) );
  OAI21_X1 U88 ( .B1(n24), .B2(n103), .A(n292), .ZN(alu_a_e[18]) );
  OAI21_X1 U89 ( .B1(n49), .B2(n108), .A(n297), .ZN(alu_a_e[13]) );
  OAI21_X1 U90 ( .B1(n50), .B2(n107), .A(n296), .ZN(alu_a_e[14]) );
  OAI21_X2 U91 ( .B1(n29), .B2(n93), .A(n281), .ZN(alu_a_e[28]) );
  OAI21_X1 U92 ( .B1(n29), .B2(n96), .A(n284), .ZN(alu_a_e[25]) );
  OAI21_X1 U93 ( .B1(n19), .B2(n90), .A(n277), .ZN(alu_a_e[31]) );
  NAND2_X1 U94 ( .A1(n32), .A2(n275), .ZN(alu_a_e[4]) );
  OAI21_X1 U95 ( .B1(n50), .B2(n111), .A(n300), .ZN(alu_a_e[10]) );
  OAI21_X1 U96 ( .B1(n28), .B2(n115), .A(n273), .ZN(alu_a_e[6]) );
  OR2_X1 U97 ( .A1(n29), .A2(n117), .ZN(n32) );
  INV_X1 U98 ( .A(n269), .ZN(n188) );
  BUF_X1 U99 ( .A(n54), .Z(n37) );
  BUF_X1 U100 ( .A(n54), .Z(n38) );
  BUF_X1 U101 ( .A(n54), .Z(n39) );
  BUF_X1 U102 ( .A(n150), .Z(n43) );
  BUF_X1 U103 ( .A(n150), .Z(n44) );
  BUF_X1 U104 ( .A(n151), .Z(n40) );
  BUF_X1 U105 ( .A(n151), .Z(n41) );
  BUF_X1 U106 ( .A(n150), .Z(n45) );
  BUF_X1 U107 ( .A(n151), .Z(n42) );
  INV_X1 U108 ( .A(rf_dout1_e[31]), .ZN(n90) );
  INV_X1 U109 ( .A(rf_dout1_e[30]), .ZN(n91) );
  INV_X1 U110 ( .A(rf_dout1_e[7]), .ZN(n114) );
  INV_X1 U111 ( .A(rf_dout1_e[16]), .ZN(n105) );
  INV_X1 U112 ( .A(rf_dout1_e[18]), .ZN(n103) );
  INV_X1 U113 ( .A(rf_dout1_e[20]), .ZN(n101) );
  INV_X1 U114 ( .A(rf_dout1_e[17]), .ZN(n104) );
  INV_X1 U115 ( .A(rf_dout1_e[19]), .ZN(n102) );
  INV_X1 U116 ( .A(rf_dout1_e[22]), .ZN(n99) );
  INV_X1 U117 ( .A(rf_dout1_e[21]), .ZN(n100) );
  INV_X1 U118 ( .A(rf_dout1_e[23]), .ZN(n98) );
  INV_X1 U119 ( .A(rf_dout1_e[8]), .ZN(n113) );
  INV_X1 U120 ( .A(rf_dout1_e[6]), .ZN(n115) );
  INV_X1 U121 ( .A(rf_dout1_e[29]), .ZN(n92) );
  INV_X1 U122 ( .A(rf_dout1_e[24]), .ZN(n97) );
  INV_X1 U123 ( .A(rf_dout1_e[26]), .ZN(n95) );
  INV_X1 U124 ( .A(rf_dout1_e[27]), .ZN(n94) );
  INV_X1 U125 ( .A(rf_dout1_e[9]), .ZN(n112) );
  INV_X1 U126 ( .A(rf_dout1_e[12]), .ZN(n109) );
  INV_X1 U127 ( .A(rf_dout1_e[10]), .ZN(n111) );
  INV_X1 U128 ( .A(rf_dout1_e[14]), .ZN(n107) );
  INV_X1 U129 ( .A(rf_dout1_e[11]), .ZN(n110) );
  INV_X1 U130 ( .A(rf_dout1_e[13]), .ZN(n108) );
  INV_X1 U131 ( .A(rf_dout1_e[15]), .ZN(n106) );
  INV_X1 U132 ( .A(rf_dout1_e[28]), .ZN(n93) );
  INV_X1 U133 ( .A(n182), .ZN(n306) );
  AOI222_X1 U134 ( .A1(dmem_dout_wb[0]), .A2(n46), .B1(alu_out_wb[0]), .B2(n43), .C1(pc_pls_4_wb[0]), .C2(n40), .ZN(n182) );
  INV_X1 U135 ( .A(n171), .ZN(n305) );
  AOI222_X1 U136 ( .A1(dmem_dout_wb[1]), .A2(n47), .B1(alu_out_wb[1]), .B2(n43), .C1(pc_pls_4_wb[1]), .C2(n40), .ZN(n171) );
  INV_X1 U137 ( .A(n160), .ZN(n304) );
  AOI222_X1 U138 ( .A1(dmem_dout_wb[2]), .A2(n48), .B1(alu_out_wb[2]), .B2(n44), .C1(pc_pls_4_wb[2]), .C2(n41), .ZN(n160) );
  INV_X1 U139 ( .A(n157), .ZN(n303) );
  AOI222_X1 U140 ( .A1(dmem_dout_wb[3]), .A2(n48), .B1(alu_out_wb[3]), .B2(n45), .C1(pc_pls_4_wb[3]), .C2(n42), .ZN(n157) );
  INV_X1 U141 ( .A(n156), .ZN(n252) );
  AOI222_X1 U142 ( .A1(dmem_dout_wb[4]), .A2(n48), .B1(alu_out_wb[4]), .B2(n45), .C1(pc_pls_4_wb[4]), .C2(n42), .ZN(n156) );
  INV_X1 U143 ( .A(n155), .ZN(n216) );
  AOI222_X1 U144 ( .A1(dmem_dout_wb[5]), .A2(n48), .B1(alu_out_wb[5]), .B2(n45), .C1(pc_pls_4_wb[5]), .C2(n42), .ZN(n155) );
  INV_X1 U145 ( .A(n154), .ZN(n215) );
  AOI222_X1 U146 ( .A1(dmem_dout_wb[6]), .A2(n48), .B1(alu_out_wb[6]), .B2(n45), .C1(pc_pls_4_wb[6]), .C2(n42), .ZN(n154) );
  INV_X1 U147 ( .A(n153), .ZN(n214) );
  AOI222_X1 U148 ( .A1(dmem_dout_wb[7]), .A2(n48), .B1(alu_out_wb[7]), .B2(n45), .C1(pc_pls_4_wb[7]), .C2(n42), .ZN(n153) );
  INV_X1 U149 ( .A(n152), .ZN(n213) );
  AOI222_X1 U150 ( .A1(dmem_dout_wb[8]), .A2(n48), .B1(alu_out_wb[8]), .B2(n45), .C1(pc_pls_4_wb[8]), .C2(n42), .ZN(n152) );
  INV_X1 U151 ( .A(n149), .ZN(n212) );
  AOI222_X1 U152 ( .A1(dmem_dout_wb[9]), .A2(n48), .B1(alu_out_wb[9]), .B2(n45), .C1(pc_pls_4_wb[9]), .C2(n42), .ZN(n149) );
  INV_X1 U153 ( .A(n181), .ZN(n211) );
  AOI222_X1 U154 ( .A1(dmem_dout_wb[10]), .A2(n46), .B1(alu_out_wb[10]), .B2(
        n43), .C1(pc_pls_4_wb[10]), .C2(n40), .ZN(n181) );
  INV_X1 U155 ( .A(n180), .ZN(n210) );
  AOI222_X1 U156 ( .A1(dmem_dout_wb[11]), .A2(n46), .B1(alu_out_wb[11]), .B2(
        n43), .C1(pc_pls_4_wb[11]), .C2(n40), .ZN(n180) );
  INV_X1 U157 ( .A(n179), .ZN(n209) );
  AOI222_X1 U158 ( .A1(dmem_dout_wb[12]), .A2(n46), .B1(alu_out_wb[12]), .B2(
        n43), .C1(pc_pls_4_wb[12]), .C2(n40), .ZN(n179) );
  INV_X1 U159 ( .A(n178), .ZN(n208) );
  AOI222_X1 U160 ( .A1(dmem_dout_wb[13]), .A2(n46), .B1(alu_out_wb[13]), .B2(
        n43), .C1(pc_pls_4_wb[13]), .C2(n40), .ZN(n178) );
  INV_X1 U161 ( .A(n177), .ZN(n207) );
  AOI222_X1 U162 ( .A1(dmem_dout_wb[14]), .A2(n46), .B1(alu_out_wb[14]), .B2(
        n43), .C1(pc_pls_4_wb[14]), .C2(n40), .ZN(n177) );
  INV_X1 U163 ( .A(n176), .ZN(n206) );
  AOI222_X1 U164 ( .A1(dmem_dout_wb[15]), .A2(n46), .B1(alu_out_wb[15]), .B2(
        n43), .C1(pc_pls_4_wb[15]), .C2(n40), .ZN(n176) );
  INV_X1 U165 ( .A(n175), .ZN(n205) );
  AOI222_X1 U166 ( .A1(dmem_dout_wb[16]), .A2(n46), .B1(alu_out_wb[16]), .B2(
        n43), .C1(pc_pls_4_wb[16]), .C2(n40), .ZN(n175) );
  INV_X1 U167 ( .A(n174), .ZN(n204) );
  AOI222_X1 U168 ( .A1(dmem_dout_wb[17]), .A2(n46), .B1(alu_out_wb[17]), .B2(
        n43), .C1(pc_pls_4_wb[17]), .C2(n40), .ZN(n174) );
  INV_X1 U169 ( .A(n173), .ZN(n203) );
  AOI222_X1 U170 ( .A1(dmem_dout_wb[18]), .A2(n46), .B1(alu_out_wb[18]), .B2(
        n43), .C1(pc_pls_4_wb[18]), .C2(n40), .ZN(n173) );
  INV_X1 U171 ( .A(n172), .ZN(n202) );
  AOI222_X1 U172 ( .A1(dmem_dout_wb[19]), .A2(n47), .B1(alu_out_wb[19]), .B2(
        n43), .C1(pc_pls_4_wb[19]), .C2(n40), .ZN(n172) );
  INV_X1 U173 ( .A(n170), .ZN(n201) );
  AOI222_X1 U174 ( .A1(dmem_dout_wb[20]), .A2(n47), .B1(alu_out_wb[20]), .B2(
        n44), .C1(pc_pls_4_wb[20]), .C2(n41), .ZN(n170) );
  INV_X1 U175 ( .A(n169), .ZN(n200) );
  AOI222_X1 U176 ( .A1(dmem_dout_wb[21]), .A2(n47), .B1(alu_out_wb[21]), .B2(
        n44), .C1(pc_pls_4_wb[21]), .C2(n41), .ZN(n169) );
  INV_X1 U177 ( .A(n168), .ZN(n199) );
  AOI222_X1 U178 ( .A1(dmem_dout_wb[22]), .A2(n47), .B1(alu_out_wb[22]), .B2(
        n44), .C1(pc_pls_4_wb[22]), .C2(n41), .ZN(n168) );
  INV_X1 U179 ( .A(n167), .ZN(n198) );
  AOI222_X1 U180 ( .A1(dmem_dout_wb[23]), .A2(n47), .B1(alu_out_wb[23]), .B2(
        n44), .C1(pc_pls_4_wb[23]), .C2(n41), .ZN(n167) );
  INV_X1 U181 ( .A(n166), .ZN(n197) );
  AOI222_X1 U182 ( .A1(dmem_dout_wb[24]), .A2(n47), .B1(alu_out_wb[24]), .B2(
        n44), .C1(pc_pls_4_wb[24]), .C2(n41), .ZN(n166) );
  INV_X1 U183 ( .A(n165), .ZN(n196) );
  AOI222_X1 U184 ( .A1(dmem_dout_wb[25]), .A2(n47), .B1(alu_out_wb[25]), .B2(
        n44), .C1(pc_pls_4_wb[25]), .C2(n41), .ZN(n165) );
  INV_X1 U185 ( .A(n164), .ZN(n195) );
  AOI222_X1 U186 ( .A1(dmem_dout_wb[26]), .A2(n47), .B1(alu_out_wb[26]), .B2(
        n44), .C1(pc_pls_4_wb[26]), .C2(n41), .ZN(n164) );
  INV_X1 U187 ( .A(n163), .ZN(n194) );
  AOI222_X1 U188 ( .A1(dmem_dout_wb[27]), .A2(n47), .B1(alu_out_wb[27]), .B2(
        n44), .C1(pc_pls_4_wb[27]), .C2(n41), .ZN(n163) );
  INV_X1 U189 ( .A(n162), .ZN(n193) );
  AOI222_X1 U190 ( .A1(dmem_dout_wb[28]), .A2(n47), .B1(alu_out_wb[28]), .B2(
        n44), .C1(pc_pls_4_wb[28]), .C2(n41), .ZN(n162) );
  INV_X1 U191 ( .A(n161), .ZN(n192) );
  AOI222_X1 U193 ( .A1(dmem_dout_wb[29]), .A2(n47), .B1(alu_out_wb[29]), .B2(
        n44), .C1(pc_pls_4_wb[29]), .C2(n41), .ZN(n161) );
  INV_X1 U194 ( .A(n159), .ZN(n191) );
  AOI222_X1 U195 ( .A1(dmem_dout_wb[30]), .A2(n48), .B1(alu_out_wb[30]), .B2(
        n44), .C1(pc_pls_4_wb[30]), .C2(n41), .ZN(n159) );
  INV_X1 U196 ( .A(n158), .ZN(n190) );
  AOI222_X1 U197 ( .A1(dmem_dout_wb[31]), .A2(n48), .B1(alu_out_wb[31]), .B2(
        n45), .C1(pc_pls_4_wb[31]), .C2(n42), .ZN(n158) );
  INV_X1 U198 ( .A(rf_dout1_e[5]), .ZN(n116) );
  INV_X1 U199 ( .A(rf_dout1_e[4]), .ZN(n117) );
  NAND2_X1 U201 ( .A1(instr_d[15]), .A2(n307), .ZN(n227) );
  INV_X1 U202 ( .A(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n307) );
  NOR4_X1 U203 ( .A1(rf_dout1_e[23]), .A2(rf_dout1_e[22]), .A3(rf_dout1_e[21]), 
        .A4(rf_dout1_e[20]), .ZN(n222) );
  NOR4_X1 U204 ( .A1(rf_dout1_e[9]), .A2(rf_dout1_e[8]), .A3(rf_dout1_e[7]), 
        .A4(rf_dout1_e[6]), .ZN(n226) );
  INV_X1 U205 ( .A(rf_dout1_e[3]), .ZN(n118) );
  NAND2_X1 U206 ( .A1(n227), .A2(n228), .ZN(imm_d[31]) );
  NAND2_X1 U207 ( .A1(instr_d[25]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n228) );
  INV_X1 U208 ( .A(rf_dout1_e[0]), .ZN(n121) );
  INV_X1 U209 ( .A(n255), .ZN(net23138) );
  INV_X1 U210 ( .A(n262), .ZN(net23132) );
  INV_X1 U211 ( .A(n256), .ZN(n129) );
  INV_X1 U212 ( .A(n251), .ZN(n126) );
  INV_X1 U213 ( .A(n260), .ZN(n132) );
  INV_X1 U214 ( .A(n261), .ZN(n133) );
  INV_X1 U215 ( .A(n238), .ZN(n140) );
  BUF_X1 U216 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n48) );
  INV_X1 U217 ( .A(n267), .ZN(n138) );
  BUF_X1 U218 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n46) );
  BUF_X1 U219 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n47) );
  INV_X1 U220 ( .A(n263), .ZN(n134) );
  INV_X1 U221 ( .A(n254), .ZN(n128) );
  INV_X1 U222 ( .A(n266), .ZN(n137) );
  INV_X1 U223 ( .A(n264), .ZN(n135) );
  INV_X1 U224 ( .A(n253), .ZN(n127) );
  INV_X1 U225 ( .A(n248), .ZN(n123) );
  INV_X1 U226 ( .A(n268), .ZN(n139) );
  INV_X1 U227 ( .A(n249), .ZN(n124) );
  INV_X1 U228 ( .A(n246), .ZN(n122) );
  INV_X1 U229 ( .A(\CTRL_WORD[R_TYPE_SEL] ), .ZN(n308) );
  NAND2_X1 U230 ( .A1(n227), .A2(n237), .ZN(imm_d[16]) );
  NAND2_X1 U231 ( .A1(instr_d[16]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n237) );
  NAND2_X1 U232 ( .A1(n227), .A2(n236), .ZN(imm_d[17]) );
  NAND2_X1 U233 ( .A1(instr_d[17]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n236) );
  NAND2_X1 U234 ( .A1(n227), .A2(n235), .ZN(imm_d[18]) );
  NAND2_X1 U235 ( .A1(instr_d[18]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n235) );
  NAND2_X1 U236 ( .A1(n227), .A2(n234), .ZN(imm_d[19]) );
  NAND2_X1 U237 ( .A1(instr_d[19]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n234) );
  NAND2_X1 U238 ( .A1(n227), .A2(n233), .ZN(imm_d[20]) );
  NAND2_X1 U239 ( .A1(instr_d[20]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n233) );
  NAND2_X1 U240 ( .A1(n227), .A2(n232), .ZN(imm_d[21]) );
  NAND2_X1 U241 ( .A1(instr_d[21]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n232) );
  INV_X1 U242 ( .A(rf_dout1_e[2]), .ZN(n119) );
  OR2_X1 U243 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[2]), .ZN(
        rf_waddr_d[2]) );
  OR2_X1 U244 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[0]), .ZN(
        rf_waddr_d[0]) );
  OR2_X1 U245 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[1]), .ZN(
        rf_waddr_d[1]) );
  INV_X1 U246 ( .A(n243), .ZN(n183) );
  NAND2_X1 U247 ( .A1(n227), .A2(n231), .ZN(imm_d[22]) );
  NAND2_X1 U248 ( .A1(instr_d[22]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n231) );
  NAND2_X1 U249 ( .A1(n227), .A2(n230), .ZN(imm_d[23]) );
  NAND2_X1 U250 ( .A1(instr_d[23]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n230) );
  NAND2_X1 U251 ( .A1(n227), .A2(n229), .ZN(imm_d[24]) );
  NAND2_X1 U252 ( .A1(instr_d[24]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n229) );
  NOR2_X1 U253 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(n46), .ZN(n150) );
  NAND4_X1 U254 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(n218) );
  NOR4_X1 U255 ( .A1(rf_dout1_e[12]), .A2(rf_dout1_e[11]), .A3(rf_dout1_e[10]), 
        .A4(rf_dout1_e[0]), .ZN(n219) );
  NOR4_X1 U256 ( .A1(rf_dout1_e[16]), .A2(rf_dout1_e[15]), .A3(rf_dout1_e[14]), 
        .A4(rf_dout1_e[13]), .ZN(n220) );
  NOR4_X1 U257 ( .A1(rf_dout1_e[1]), .A2(rf_dout1_e[19]), .A3(rf_dout1_e[18]), 
        .A4(rf_dout1_e[17]), .ZN(n221) );
  NAND4_X1 U258 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(n217) );
  NOR4_X1 U259 ( .A1(rf_dout1_e[27]), .A2(rf_dout1_e[26]), .A3(rf_dout1_e[25]), 
        .A4(rf_dout1_e[24]), .ZN(n223) );
  NOR4_X1 U260 ( .A1(rf_dout1_e[30]), .A2(rf_dout1_e[2]), .A3(rf_dout1_e[29]), 
        .A4(rf_dout1_e[28]), .ZN(n224) );
  NOR4_X1 U261 ( .A1(rf_dout1_e[5]), .A2(rf_dout1_e[4]), .A3(rf_dout1_e[3]), 
        .A4(rf_dout1_e[31]), .ZN(n225) );
  NOR2_X1 U262 ( .A1(n309), .A2(n46), .ZN(n151) );
  INV_X1 U263 ( .A(\CTRL_WORD[JAL_EN] ), .ZN(n309) );
  INV_X1 U264 ( .A(rf_dout1_e[25]), .ZN(n96) );
  INV_X1 U265 ( .A(rf_dout1_e[1]), .ZN(n120) );
  OR2_X1 U266 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[4]), .ZN(
        rf_waddr_d[4]) );
  OR2_X1 U267 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[3]), .ZN(
        rf_waddr_d[3]) );
  NOR2_X1 U268 ( .A1(n217), .A2(n218), .ZN(n302) );
  AND2_X1 U269 ( .A1(DMEM_RWADDR[31]), .A2(n184), .ZN(\npc_f[31] ) );
  INV_X1 U270 ( .A(n148), .ZN(n89) );
  AOI22_X1 U271 ( .A1(rs2_e[0]), .A2(n308), .B1(rs3_e[0]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n148) );
  INV_X1 U272 ( .A(n147), .ZN(n88) );
  AOI22_X1 U273 ( .A1(rs2_e[1]), .A2(n308), .B1(rs3_e[1]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n147) );
  INV_X1 U274 ( .A(n146), .ZN(n87) );
  AOI22_X1 U275 ( .A1(rs2_e[2]), .A2(n308), .B1(rs3_e[2]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n146) );
  INV_X1 U276 ( .A(n145), .ZN(n86) );
  AOI22_X1 U277 ( .A1(rs2_e[3]), .A2(n308), .B1(rs3_e[3]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n145) );
  INV_X1 U278 ( .A(n144), .ZN(n85) );
  AOI22_X1 U279 ( .A1(rs2_e[4]), .A2(n308), .B1(rs3_e[4]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n144) );
  BUF_X2 U280 ( .A(RST_AN), .Z(n51) );
  BUF_X2 U281 ( .A(RST_AN), .Z(n52) );
  BUF_X2 U282 ( .A(n35), .Z(n34) );
  NAND2_X1 U283 ( .A1(pc_pls_4_e[26]), .A2(n34), .ZN(n283) );
  NAND2_X1 U284 ( .A1(n36), .A2(pc_pls_4_e[23]), .ZN(n286) );
  NAND2_X1 U285 ( .A1(pc_pls_4_e[21]), .A2(n34), .ZN(n288) );
  NAND2_X1 U286 ( .A1(pc_pls_4_e[22]), .A2(n36), .ZN(n287) );
  NAND2_X1 U287 ( .A1(pc_pls_4_e[19]), .A2(n24), .ZN(n291) );
  NAND2_X1 U288 ( .A1(pc_pls_4_e[20]), .A2(n29), .ZN(n289) );
  NAND2_X1 U289 ( .A1(pc_pls_4_e[17]), .A2(n33), .ZN(n293) );
  NAND2_X1 U290 ( .A1(pc_pls_4_e[18]), .A2(n36), .ZN(n292) );
  NAND2_X1 U291 ( .A1(pc_pls_4_e[3]), .A2(n29), .ZN(n276) );
  NAND2_X1 U292 ( .A1(pc_pls_4_e[5]), .A2(n49), .ZN(n274) );
  INV_X1 U293 ( .A(net25874), .ZN(net25862) );
  NAND2_X1 U294 ( .A1(pc_pls_4_e[1]), .A2(n29), .ZN(n290) );
  OAI21_X1 U295 ( .B1(n23), .B2(n118), .A(n276), .ZN(alu_a_e[3]) );
  NAND2_X1 U296 ( .A1(pc_pls_4_e[4]), .A2(n19), .ZN(n275) );
  OAI21_X1 U297 ( .B1(n50), .B2(n121), .A(n301), .ZN(alu_a_e[0]) );
  NAND2_X1 U298 ( .A1(pc_pls_4_e[30]), .A2(n23), .ZN(n278) );
  NAND2_X1 U299 ( .A1(pc_pls_4_e[28]), .A2(n31), .ZN(n281) );
  NAND2_X1 U300 ( .A1(pc_pls_4_e[29]), .A2(n50), .ZN(n280) );
  NAND2_X1 U301 ( .A1(pc_pls_4_e[25]), .A2(n19), .ZN(n284) );
  NAND2_X1 U302 ( .A1(pc_pls_4_e[27]), .A2(n33), .ZN(n282) );
  NAND2_X1 U303 ( .A1(pc_pls_4_e[24]), .A2(n29), .ZN(n285) );
  NAND2_X1 U304 ( .A1(pc_pls_4_e[31]), .A2(n36), .ZN(n277) );
  NAND2_X1 U305 ( .A1(n49), .A2(pc_pls_4_e[2]), .ZN(n279) );
  NAND2_X1 U306 ( .A1(pc_pls_4_e[15]), .A2(n34), .ZN(n295) );
  NAND2_X1 U307 ( .A1(pc_pls_4_e[16]), .A2(n31), .ZN(n294) );
  NAND2_X1 U308 ( .A1(pc_pls_4_e[13]), .A2(n36), .ZN(n297) );
  NAND2_X1 U309 ( .A1(pc_pls_4_e[14]), .A2(n31), .ZN(n296) );
  NAND2_X1 U310 ( .A1(pc_pls_4_e[11]), .A2(n31), .ZN(n299) );
  NAND2_X1 U311 ( .A1(pc_pls_4_e[9]), .A2(n24), .ZN(n270) );
  NAND2_X1 U312 ( .A1(pc_pls_4_e[10]), .A2(n28), .ZN(n300) );
  NAND2_X1 U313 ( .A1(pc_pls_4_e[12]), .A2(n29), .ZN(n298) );
  NAND2_X1 U314 ( .A1(pc_pls_4_e[7]), .A2(n34), .ZN(n272) );
  NAND2_X1 U315 ( .A1(pc_pls_4_e[8]), .A2(n49), .ZN(n271) );
  NAND2_X1 U316 ( .A1(pc_pls_4_e[6]), .A2(n36), .ZN(n273) );
  INV_X1 U317 ( .A(net25888), .ZN(net25860) );
  INV_X1 U318 ( .A(n247), .ZN(n186) );
  OAI21_X1 U319 ( .B1(n29), .B2(n119), .A(n279), .ZN(alu_a_e[2]) );
  AOI22_X1 U320 ( .A1(rf_dout2_e[9]), .A2(n7), .B1(imm_e[9]), .B2(n12), .ZN(
        n238) );
  AOI22_X1 U321 ( .A1(rf_dout2_e[7]), .A2(n16), .B1(net34728), .B2(imm_e[7]), 
        .ZN(n240) );
  AOI22_X1 U322 ( .A1(rf_dout2_e[8]), .A2(net25862), .B1(n9), .B2(imm_e[8]), 
        .ZN(n239) );
  AOI22_X1 U323 ( .A1(net25860), .A2(rf_dout2_e[6]), .B1(net25872), .B2(
        imm_e[6]), .ZN(n241) );
  AOI22_X1 U324 ( .A1(rf_dout2_e[3]), .A2(n13), .B1(n9), .B2(imm_e[3]), .ZN(
        n244) );
  AOI22_X1 U325 ( .A1(net34744), .A2(rf_dout2_e[4]), .B1(net25868), .B2(
        imm_e[4]), .ZN(n243) );
  NAND2_X1 U326 ( .A1(n49), .A2(pc_pls_4_e[0]), .ZN(n301) );
  AOI22_X1 U327 ( .A1(rf_dout2_e[26]), .A2(n16), .B1(net34734), .B2(imm_e[26]), 
        .ZN(n251) );
  AOI22_X1 U328 ( .A1(rf_dout2_e[21]), .A2(net25862), .B1(net34727), .B2(
        imm_e[21]), .ZN(n256) );
  AOI22_X1 U329 ( .A1(rf_dout2_e[28]), .A2(n16), .B1(net34378), .B2(imm_e[28]), 
        .ZN(n249) );
  AOI22_X1 U330 ( .A1(rf_dout2_e[20]), .A2(n14), .B1(imm_e[20]), .B2(net40517), 
        .ZN(n257) );
  AOI22_X1 U331 ( .A1(rf_dout2_e[27]), .A2(net25860), .B1(imm_e[27]), .B2(n12), 
        .ZN(n250) );
  AOI22_X1 U332 ( .A1(rf_dout2_e[30]), .A2(net40540), .B1(net34734), .B2(
        imm_e[30]), .ZN(n246) );
  AOI22_X1 U333 ( .A1(rf_dout2_e[23]), .A2(net25860), .B1(imm_e[23]), .B2(
        net25872), .ZN(n254) );
  AOI22_X1 U334 ( .A1(net25860), .A2(rf_dout2_e[29]), .B1(imm_e[29]), .B2(
        net34379), .ZN(n248) );
  AOI22_X1 U335 ( .A1(n16), .A2(rf_dout2_e[24]), .B1(n9), .B2(imm_e[24]), .ZN(
        n253) );
  AOI22_X1 U336 ( .A1(net27502), .A2(rf_dout2_e[2]), .B1(net25888), .B2(
        imm_e[2]), .ZN(n247) );
  AOI22_X1 U337 ( .A1(rf_dout2_e[19]), .A2(net34744), .B1(imm_e[19]), .B2(n15), 
        .ZN(n259) );
  AOI22_X1 U338 ( .A1(net33900), .A2(rf_dout2_e[15]), .B1(imm_e[15]), .B2(
        net34727), .ZN(n263) );
  AOI22_X1 U339 ( .A1(rf_dout2_e[13]), .A2(net33900), .B1(n1), .B2(imm_e[13]), 
        .ZN(n265) );
  AOI22_X1 U340 ( .A1(rf_dout2_e[18]), .A2(n14), .B1(imm_e[18]), .B2(net34379), 
        .ZN(n260) );
  AOI22_X1 U341 ( .A1(net25862), .A2(rf_dout2_e[17]), .B1(imm_e[17]), .B2(n15), 
        .ZN(n261) );
  AOI22_X1 U342 ( .A1(rf_dout2_e[14]), .A2(net34744), .B1(net25868), .B2(
        imm_e[14]), .ZN(n264) );
  AOI22_X1 U343 ( .A1(n14), .A2(rf_dout2_e[11]), .B1(net25872), .B2(imm_e[11]), 
        .ZN(n267) );
  AOI22_X1 U344 ( .A1(n14), .A2(rf_dout2_e[12]), .B1(n1), .B2(imm_e[12]), .ZN(
        n266) );
  AOI22_X1 U345 ( .A1(rf_dout2_e[10]), .A2(n7), .B1(imm_e[10]), .B2(net34728), 
        .ZN(n268) );
  AOI22_X1 U346 ( .A1(net40540), .A2(rf_dout2_e[0]), .B1(n11), .B2(imm_e[0]), 
        .ZN(n269) );
  AOI22_X1 U347 ( .A1(n13), .A2(rf_dout2_e[1]), .B1(net34378), .B2(imm_e[1]), 
        .ZN(n258) );
  XOR2_X1 U348 ( .A(\DP_SIG[CMPR_0_IS_0_M] ), .B(\CTRL_WORD[COMP_0_INVERT] ), 
        .Z(n53) );
  MUX2_X1 U349 ( .A(\CTRL_WORD[JUMP_EN] ), .B(n53), .S(\CTRL_WORD[BRANCH_EN] ), 
        .Z(n184) );
  INV_X1 U350 ( .A(n184), .ZN(n54) );
  MUX2_X1 U351 ( .A(DMEM_RWADDR[0]), .B(pc_pls_4_f[0]), .S(n37), .Z(n189) );
  MUX2_X1 U352 ( .A(DMEM_RWADDR[1]), .B(pc_pls_4_f[1]), .S(n37), .Z(n84) );
  MUX2_X1 U353 ( .A(DMEM_RWADDR[2]), .B(pc_pls_4_f[2]), .S(n37), .Z(n83) );
  MUX2_X1 U354 ( .A(DMEM_RWADDR[3]), .B(pc_pls_4_f[3]), .S(n37), .Z(n82) );
  MUX2_X1 U355 ( .A(DMEM_RWADDR[4]), .B(pc_pls_4_f[4]), .S(n37), .Z(n81) );
  MUX2_X1 U356 ( .A(DMEM_RWADDR[5]), .B(pc_pls_4_f[5]), .S(n37), .Z(n80) );
  MUX2_X1 U357 ( .A(DMEM_RWADDR[6]), .B(pc_pls_4_f[6]), .S(n37), .Z(n79) );
  MUX2_X1 U358 ( .A(DMEM_RWADDR[7]), .B(pc_pls_4_f[7]), .S(n37), .Z(n78) );
  MUX2_X1 U359 ( .A(DMEM_RWADDR[8]), .B(pc_pls_4_f[8]), .S(n37), .Z(n77) );
  MUX2_X1 U360 ( .A(DMEM_RWADDR[9]), .B(pc_pls_4_f[9]), .S(n37), .Z(n76) );
  MUX2_X1 U361 ( .A(DMEM_RWADDR[10]), .B(pc_pls_4_f[10]), .S(n37), .Z(n75) );
  MUX2_X1 U362 ( .A(DMEM_RWADDR[11]), .B(pc_pls_4_f[11]), .S(n38), .Z(n74) );
  MUX2_X1 U363 ( .A(DMEM_RWADDR[12]), .B(pc_pls_4_f[12]), .S(n38), .Z(n73) );
  MUX2_X1 U364 ( .A(DMEM_RWADDR[13]), .B(pc_pls_4_f[13]), .S(n38), .Z(n72) );
  MUX2_X1 U365 ( .A(DMEM_RWADDR[14]), .B(pc_pls_4_f[14]), .S(n38), .Z(n71) );
  MUX2_X1 U366 ( .A(DMEM_RWADDR[15]), .B(pc_pls_4_f[15]), .S(n38), .Z(n70) );
  MUX2_X1 U367 ( .A(DMEM_RWADDR[16]), .B(pc_pls_4_f[16]), .S(n38), .Z(n69) );
  MUX2_X1 U368 ( .A(DMEM_RWADDR[17]), .B(pc_pls_4_f[17]), .S(n38), .Z(n68) );
  MUX2_X1 U369 ( .A(DMEM_RWADDR[18]), .B(pc_pls_4_f[18]), .S(n38), .Z(n67) );
  MUX2_X1 U370 ( .A(DMEM_RWADDR[19]), .B(pc_pls_4_f[19]), .S(n38), .Z(n66) );
  MUX2_X1 U371 ( .A(DMEM_RWADDR[20]), .B(pc_pls_4_f[20]), .S(n38), .Z(n65) );
  MUX2_X1 U372 ( .A(DMEM_RWADDR[21]), .B(pc_pls_4_f[21]), .S(n38), .Z(n64) );
  MUX2_X1 U373 ( .A(DMEM_RWADDR[22]), .B(pc_pls_4_f[22]), .S(n39), .Z(n63) );
  MUX2_X1 U374 ( .A(DMEM_RWADDR[23]), .B(pc_pls_4_f[23]), .S(n39), .Z(n62) );
  MUX2_X1 U375 ( .A(DMEM_RWADDR[24]), .B(pc_pls_4_f[24]), .S(n39), .Z(n61) );
  MUX2_X1 U376 ( .A(DMEM_RWADDR[25]), .B(pc_pls_4_f[25]), .S(n39), .Z(n60) );
  MUX2_X1 U377 ( .A(DMEM_RWADDR[26]), .B(pc_pls_4_f[26]), .S(n39), .Z(n59) );
  MUX2_X1 U378 ( .A(DMEM_RWADDR[27]), .B(pc_pls_4_f[27]), .S(n39), .Z(n58) );
  MUX2_X1 U379 ( .A(DMEM_RWADDR[28]), .B(pc_pls_4_f[28]), .S(n39), .Z(n57) );
  MUX2_X1 U380 ( .A(DMEM_RWADDR[29]), .B(pc_pls_4_f[29]), .S(n39), .Z(n56) );
  MUX2_X1 U381 ( .A(DMEM_RWADDR[30]), .B(pc_pls_4_f[30]), .S(n39), .Z(n55) );
endmodule


module HU ( CLK, RST_AN, .DP_SIG({\DP_SIG[CMPR_0_IS_0_M] , 
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }), 
    .HZRD_SIG({\HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , 
        \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , 
        \HZRD_SIG[FLUSH_MWB] }) );
  input CLK, RST_AN, \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  output \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] ,
         \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] ;
  wire   n2, n3, n4, n7, \HZRD_SIG[FLUSH_DE] , n9;
  assign \HZRD_SIG[FLUSH_MWB]  = 1'b0;
  assign \HZRD_SIG[STALL_DE]  = 1'b0;
  assign \HZRD_SIG[STALL_FD]  = 1'b0;
  assign \HZRD_SIG[FLUSH_FD]  = \HZRD_SIG[FLUSH_DE] ;
  assign \HZRD_SIG[FLUSH_EM]  = \HZRD_SIG[FLUSH_DE] ;

  INV_X1 U3 ( .A(n7), .ZN(\HZRD_SIG[FLUSH_DE] ) );
  OR4_X1 U4 ( .A1(\DP_SIG[INSTR_OPCODE_M][5] ), .A2(
        \DP_SIG[INSTR_OPCODE_M][4] ), .A3(\DP_SIG[INSTR_OPCODE_M][3] ), .A4(n2), .ZN(n7) );
  AOI22_X1 U5 ( .A1(n3), .A2(\DP_SIG[INSTR_OPCODE_M][2] ), .B1(
        \DP_SIG[INSTR_OPCODE_M][1] ), .B2(n9), .ZN(n2) );
  INV_X1 U6 ( .A(\DP_SIG[INSTR_OPCODE_M][2] ), .ZN(n9) );
  NOR2_X1 U7 ( .A1(\DP_SIG[INSTR_OPCODE_M][1] ), .A2(n4), .ZN(n3) );
  XNOR2_X1 U8 ( .A(\DP_SIG[INSTR_OPCODE_M][0] ), .B(\DP_SIG[CMPR_0_IS_0_M] ), 
        .ZN(n4) );
endmodule


module CPU_1 ( CLK, RST_AN, IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, DMEM_WEN, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN;
  output DMEM_WEN;
  wire   \hzrd_sig[FLUSH_FD] , \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] ,
         \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] ,
         \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] ,
         \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] ,
         \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] ,
         \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] ,
         \ctrl_word[COMP_0_INVERT] , \ctrl_word[RF_WB_DMEM_DOUT_SEL] ,
         \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] , \dp_sig[CMPR_0_IS_0_M] ,
         \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] ,
         \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] ,
         \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] ;
  wire   [31:0] instr_cu;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  CU U_CU ( .CLK(CLK), .RST_AN(RST_AN), .INSTR(instr_cu), .HZRD_SIG({1'b0, 
        \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        1'b0}), .CTRL_WORD({\ctrl_word[J_TYPE_IMM_SEL] , 
        \ctrl_word[R_TYPE_SEL] , \ctrl_word[IMM_SEL] , 
        \ctrl_word[PC_PLS_4_SEL] , \ctrl_word[ALU_FUNC][3] , 
        \ctrl_word[ALU_FUNC][2] , \ctrl_word[ALU_FUNC][1] , 
        \ctrl_word[ALU_FUNC][0] , \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }) );
  DATAPATH_1 U_DATAPATH ( .CLK(CLK), .RST_AN(RST_AN), .CTRL_WORD({
        \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] , 
        \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] , 
        \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] , 
        \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] , 
        \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }), .INSTR_CU(instr_cu), 
        .HZRD_SIG({1'b0, \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , 
        \hzrd_sig[FLUSH_EM] , 1'b0}), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), 
        .IMEM_ADDR(IMEM_ADDR), .IMEM_DOUT(IMEM_DOUT), .DMEM_RWADDR(DMEM_RWADDR), .DMEM_DIN(DMEM_DIN), .DMEM_DOUT(DMEM_DOUT) );
  HU U_HU ( .CLK(CLK), .RST_AN(RST_AN), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), .HZRD_SIG(
        {SYNOPSYS_UNCONNECTED__0, \hzrd_sig[FLUSH_FD] , 
        SYNOPSYS_UNCONNECTED__1, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        SYNOPSYS_UNCONNECTED__2}) );
endmodule

