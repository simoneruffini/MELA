
module CU ( CLK, RST_AN, INSTR, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .CTRL_WORD({
        \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] , 
        \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] , 
        \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] , 
        \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] , 
        \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }) );
  input [31:0] INSTR;
  input CLK, RST_AN, \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] ;
  wire   INSTR_31, INSTR_30, INSTR_29, INSTR_28, INSTR_27, INSTR_26,
         \execute_sig_d1[R_TYPE_SEL] , \execute_sig_d1[IMM_SEL] ,
         \execute_sig_d1[PC_PLS_4_SEL] , \execute_sig_d1[ALU_FUNC][3] ,
         \execute_sig_d1[ALU_FUNC][2] , \execute_sig_d1[ALU_FUNC][1] ,
         \execute_sig_d1[ALU_FUNC][0] , \memory_sig_d1[DMEM_WEN] ,
         \memory_sig_d1[BRANCH_EN] , \memory_sig_d1[JUMP_EN] ,
         \memory_sig_d1[COMP_0_INVERT] ,
         \writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d1[JAL_EN] ,
         \writeback_sig_d1[RF_WEN] , \memory_sig_d2[DMEM_WEN] ,
         \memory_sig_d2[BRANCH_EN] , \memory_sig_d2[JUMP_EN] ,
         \memory_sig_d2[COMP_0_INVERT] ,
         \writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d2[JAL_EN] ,
         \writeback_sig_d2[RF_WEN] , \writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ,
         \writeback_sig_d3[JAL_EN] , \writeback_sig_d3[RF_WEN] , N213, N214,
         N215, N216, N217, N218, N224, N228, N229, N231, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n117, n118, n119, n120, n121, n122
;
  assign INSTR_31 = INSTR[31];
  assign INSTR_30 = INSTR[30];
  assign INSTR_29 = INSTR[29];
  assign INSTR_28 = INSTR[28];
  assign INSTR_27 = INSTR[27];
  assign INSTR_26 = INSTR[26];

  DFFR_X1 \decode_sig_d1_reg[J_TYPE_IMM_SEL]  ( .D(n36), .CK(CLK), .RN(n28), 
        .Q(\CTRL_WORD[J_TYPE_IMM_SEL] ) );
  SDFFR_X1 \execute_sig_d1_reg[R_TYPE_SEL]  ( .D(1'b0), .SI(n39), .SE(n42), 
        .CK(CLK), .RN(n29), .Q(\execute_sig_d1[R_TYPE_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[IMM_SEL]  ( .D(N218), .CK(CLK), .RN(n28), .Q(
        \execute_sig_d1[IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[PC_PLS_4_SEL]  ( .D(N217), .CK(CLK), .RN(n28), 
        .Q(\execute_sig_d1[PC_PLS_4_SEL] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][3]  ( .D(N216), .CK(CLK), .SN(n31), 
        .Q(\execute_sig_d1[ALU_FUNC][3] ) );
  DFFR_X1 \execute_sig_d1_reg[ALU_FUNC][2]  ( .D(N215), .CK(CLK), .RN(n28), 
        .Q(\execute_sig_d1[ALU_FUNC][2] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][1]  ( .D(N214), .CK(CLK), .SN(n31), 
        .Q(\execute_sig_d1[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][0]  ( .D(N213), .CK(CLK), .SN(n31), 
        .Q(\execute_sig_d1[ALU_FUNC][0] ) );
  SDFFR_X1 \memory_sig_d1_reg[DMEM_WEN]  ( .D(1'b0), .SI(n34), .SE(INSTR_29), 
        .CK(CLK), .RN(n29), .Q(\memory_sig_d1[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d1_reg[BRANCH_EN]  ( .D(n37), .CK(CLK), .RN(n28), .Q(
        \memory_sig_d1[BRANCH_EN] ) );
  DFFR_X1 \memory_sig_d1_reg[JUMP_EN]  ( .D(n36), .CK(CLK), .RN(n28), .Q(
        \memory_sig_d1[JUMP_EN] ) );
  SDFFR_X1 \memory_sig_d1_reg[COMP_0_INVERT]  ( .D(1'b0), .SI(n37), .SE(
        INSTR_26), .CK(CLK), .RN(n28), .Q(\memory_sig_d1[COMP_0_INVERT] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n34), .CK(CLK), 
        .RN(n28), .Q(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ) );
  SDFFR_X1 \writeback_sig_d1_reg[JAL_EN]  ( .D(1'b0), .SI(n36), .SE(INSTR_26), 
        .CK(CLK), .RN(n28), .Q(\writeback_sig_d1[JAL_EN] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WEN]  ( .D(N224), .CK(CLK), .RN(n28), .Q(
        \writeback_sig_d1[RF_WEN] ) );
  SDFFR_X1 \execute_sig_d2_reg[R_TYPE_SEL]  ( .D(1'b0), .SI(n33), .SE(
        \execute_sig_d1[R_TYPE_SEL] ), .CK(CLK), .RN(n29), .Q(
        \CTRL_WORD[R_TYPE_SEL] ) );
  SDFFR_X1 \execute_sig_d2_reg[IMM_SEL]  ( .D(1'b0), .SI(n33), .SE(
        \execute_sig_d1[IMM_SEL] ), .CK(CLK), .RN(n29), .Q(
        \CTRL_WORD[IMM_SEL] ) );
  SDFFR_X1 \execute_sig_d2_reg[PC_PLS_4_SEL]  ( .D(1'b0), .SI(n33), .SE(
        \execute_sig_d1[PC_PLS_4_SEL] ), .CK(CLK), .RN(n29), .Q(
        \CTRL_WORD[PC_PLS_4_SEL] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][3]  ( .D(N231), .CK(CLK), .SN(n30), 
        .Q(\CTRL_WORD[ALU_FUNC][3] ) );
  SDFFR_X1 \execute_sig_d2_reg[ALU_FUNC][2]  ( .D(1'b0), .SI(n33), .SE(
        \execute_sig_d1[ALU_FUNC][2] ), .CK(CLK), .RN(n29), .Q(
        \CTRL_WORD[ALU_FUNC][2] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][1]  ( .D(N229), .CK(CLK), .SN(n31), 
        .Q(\CTRL_WORD[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][0]  ( .D(N228), .CK(CLK), .SN(n30), 
        .Q(\CTRL_WORD[ALU_FUNC][0] ) );
  SDFFR_X1 \memory_sig_d2_reg[DMEM_WEN]  ( .D(1'b0), .SI(n33), .SE(
        \memory_sig_d1[DMEM_WEN] ), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d2[DMEM_WEN] ) );
  SDFFR_X1 \memory_sig_d2_reg[BRANCH_EN]  ( .D(1'b0), .SI(n33), .SE(
        \memory_sig_d1[BRANCH_EN] ), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d2[BRANCH_EN] ) );
  SDFFR_X1 \memory_sig_d2_reg[JUMP_EN]  ( .D(1'b0), .SI(n33), .SE(
        \memory_sig_d1[JUMP_EN] ), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d2[JUMP_EN] ) );
  SDFFR_X1 \memory_sig_d2_reg[COMP_0_INVERT]  ( .D(1'b0), .SI(n33), .SE(
        \memory_sig_d1[COMP_0_INVERT] ), .CK(CLK), .RN(n29), .Q(
        \memory_sig_d2[COMP_0_INVERT] ) );
  SDFFR_X1 \writeback_sig_d2_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(1'b0), .SI(n33), 
        .SE(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ), .CK(CLK), .RN(n29), .Q(
        \writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ) );
  SDFFR_X1 \writeback_sig_d2_reg[JAL_EN]  ( .D(1'b0), .SI(n33), .SE(
        \writeback_sig_d1[JAL_EN] ), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d2[JAL_EN] ) );
  SDFFR_X1 \writeback_sig_d2_reg[RF_WEN]  ( .D(1'b0), .SI(n33), .SE(
        \writeback_sig_d1[RF_WEN] ), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d2[RF_WEN] ) );
  SDFFR_X1 \memory_sig_d3_reg[DMEM_WEN]  ( .D(1'b0), .SI(n32), .SE(
        \memory_sig_d2[DMEM_WEN] ), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[DMEM_WEN] ) );
  SDFFR_X1 \memory_sig_d3_reg[BRANCH_EN]  ( .D(1'b0), .SI(n32), .SE(
        \memory_sig_d2[BRANCH_EN] ), .CK(CLK), .RN(n29), .Q(
        \CTRL_WORD[BRANCH_EN] ) );
  SDFFR_X1 \memory_sig_d3_reg[JUMP_EN]  ( .D(1'b0), .SI(n32), .SE(
        \memory_sig_d2[JUMP_EN] ), .CK(CLK), .RN(n30), .Q(\CTRL_WORD[JUMP_EN] ) );
  SDFFR_X1 \memory_sig_d3_reg[COMP_0_INVERT]  ( .D(1'b0), .SI(n32), .SE(
        \memory_sig_d2[COMP_0_INVERT] ), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[COMP_0_INVERT] ) );
  SDFFR_X1 \writeback_sig_d3_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(1'b0), .SI(n32), 
        .SE(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ) );
  SDFFR_X1 \writeback_sig_d4_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(1'b0), .SI(n40), 
        .SE(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ) );
  SDFFR_X1 \writeback_sig_d3_reg[JAL_EN]  ( .D(1'b0), .SI(n32), .SE(
        \writeback_sig_d2[JAL_EN] ), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d3[JAL_EN] ) );
  SDFFR_X1 \writeback_sig_d4_reg[JAL_EN]  ( .D(1'b0), .SI(n40), .SE(
        \writeback_sig_d3[JAL_EN] ), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[JAL_EN] ) );
  SDFFR_X1 \writeback_sig_d3_reg[RF_WEN]  ( .D(1'b0), .SI(n32), .SE(
        \writeback_sig_d2[RF_WEN] ), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d3[RF_WEN] ) );
  SDFFR_X1 \writeback_sig_d4_reg[RF_WEN]  ( .D(1'b0), .SI(n40), .SE(
        \writeback_sig_d3[RF_WEN] ), .CK(CLK), .RN(n28), .Q(
        \CTRL_WORD[RF_WEN] ) );
  OR2_X2 U28 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][3] ), 
        .ZN(N231) );
  OR2_X2 U29 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][1] ), 
        .ZN(N229) );
  OR2_X2 U30 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][0] ), 
        .ZN(N228) );
  AOI21_X2 U31 ( .B1(n56), .B2(n57), .A(\HZRD_SIG[FLUSH_FD] ), .ZN(N224) );
  OAI211_X2 U32 ( .C1(n58), .C2(n59), .A(n50), .B(n44), .ZN(n57) );
  NOR3_X2 U33 ( .A1(INSTR_26), .A2(INSTR_31), .A3(INSTR_27), .ZN(n59) );
  AOI211_X2 U34 ( .C1(INSTR_29), .C2(n41), .A(n52), .B(n53), .ZN(n58) );
  OAI21_X2 U35 ( .B1(n60), .B2(n61), .A(n41), .ZN(n56) );
  OAI22_X2 U36 ( .A1(n50), .A2(n47), .B1(n49), .B2(n62), .ZN(n61) );
  OAI211_X2 U37 ( .C1(n66), .C2(n67), .A(n55), .B(n54), .ZN(N218) );
  AOI21_X2 U38 ( .B1(n51), .B2(n69), .A(n60), .ZN(n66) );
  OAI211_X2 U39 ( .C1(n44), .C2(n70), .A(n71), .B(n72), .ZN(n60) );
  NAND2_X2 U40 ( .A1(n64), .A2(n55), .ZN(N217) );
  NAND4_X2 U41 ( .A1(n48), .A2(n38), .A3(n52), .A4(n44), .ZN(n64) );
  OAI221_X2 U42 ( .B1(n73), .B2(n74), .C1(n42), .C2(n75), .A(n39), .ZN(N216)
         );
  AOI221_X2 U43 ( .B1(n76), .B2(n49), .C1(INSTR_31), .C2(n77), .A(n78), .ZN(
        n75) );
  OAI221_X2 U44 ( .B1(INSTR_27), .B2(n69), .C1(n48), .C2(n44), .A(n79), .ZN(
        n78) );
  OAI22_X2 U45 ( .A1(INSTR_31), .A2(INSTR_28), .B1(n52), .B2(n50), .ZN(n80) );
  AOI21_X2 U46 ( .B1(INSTR[0]), .B2(n117), .A(n81), .ZN(n73) );
  OAI21_X2 U47 ( .B1(n82), .B2(n65), .A(n83), .ZN(N215) );
  OAI211_X2 U48 ( .C1(n84), .C2(n63), .A(n38), .B(INSTR_28), .ZN(n83) );
  NOR2_X2 U49 ( .A1(n85), .A2(INSTR_26), .ZN(n63) );
  AOI21_X2 U50 ( .B1(n72), .B2(n85), .A(n52), .ZN(n84) );
  NAND2_X2 U51 ( .A1(n86), .A2(n53), .ZN(n72) );
  NAND2_X2 U52 ( .A1(n42), .A2(n39), .ZN(n65) );
  AOI211_X2 U53 ( .C1(INSTR[1]), .C2(n87), .A(n88), .B(n89), .ZN(n82) );
  OAI211_X2 U54 ( .C1(n90), .C2(n74), .A(n91), .B(n35), .ZN(N214) );
  OAI211_X2 U55 ( .C1(n92), .C2(n46), .A(n74), .B(n41), .ZN(n91) );
  AOI22_X2 U56 ( .A1(n86), .A2(n51), .B1(n62), .B2(INSTR_30), .ZN(n93) );
  NAND2_X2 U57 ( .A1(INSTR_28), .A2(n52), .ZN(n62) );
  OAI211_X2 U58 ( .C1(INSTR_29), .C2(n94), .A(n70), .B(n95), .ZN(n92) );
  NAND2_X2 U59 ( .A1(n48), .A2(INSTR_27), .ZN(n70) );
  AOI21_X2 U60 ( .B1(n52), .B2(n50), .A(n45), .ZN(n94) );
  AOI21_X2 U61 ( .B1(n87), .B2(n119), .A(n97), .ZN(n90) );
  OAI211_X2 U62 ( .C1(n99), .C2(n74), .A(n100), .B(n35), .ZN(N213) );
  OAI221_X2 U63 ( .B1(n68), .B2(n41), .C1(n102), .C2(n74), .A(n39), .ZN(n101)
         );
  NOR2_X2 U64 ( .A1(n103), .A2(n89), .ZN(n102) );
  NOR4_X2 U65 ( .A1(n121), .A2(n104), .A3(n122), .A4(INSTR[5]), .ZN(n89) );
  NOR3_X2 U66 ( .A1(n104), .A2(n105), .A3(n122), .ZN(n103) );
  NOR2_X2 U67 ( .A1(n77), .A2(INSTR_30), .ZN(n68) );
  OAI211_X2 U68 ( .C1(n106), .C2(n107), .A(n74), .B(n41), .ZN(n100) );
  OAI22_X2 U69 ( .A1(INSTR_29), .A2(n43), .B1(INSTR_27), .B2(n85), .ZN(n107)
         );
  NAND2_X2 U70 ( .A1(INSTR_30), .A2(n49), .ZN(n85) );
  OAI21_X2 U71 ( .B1(INSTR_28), .B2(INSTR_27), .A(n108), .ZN(n76) );
  OAI211_X2 U72 ( .C1(n109), .C2(n52), .A(n110), .B(n95), .ZN(n106) );
  NAND2_X2 U73 ( .A1(n86), .A2(INSTR_26), .ZN(n95) );
  NOR2_X2 U74 ( .A1(n49), .A2(INSTR_30), .ZN(n86) );
  NAND2_X2 U75 ( .A1(INSTR_28), .A2(n49), .ZN(n96) );
  AOI21_X2 U76 ( .B1(INSTR_29), .B2(n50), .A(n45), .ZN(n109) );
  NAND2_X2 U77 ( .A1(INSTR_30), .A2(INSTR_26), .ZN(n69) );
  NAND4_X2 U78 ( .A1(n52), .A2(n50), .A3(n53), .A4(n111), .ZN(n74) );
  NOR3_X2 U79 ( .A1(INSTR_29), .A2(INSTR_31), .A3(INSTR_30), .ZN(n111) );
  NOR3_X2 U80 ( .A1(n112), .A2(n81), .A3(n88), .ZN(n99) );
  NOR3_X2 U81 ( .A1(INSTR[1]), .A2(INSTR[5]), .A3(n118), .ZN(n88) );
  NOR2_X2 U82 ( .A1(n104), .A2(INSTR[0]), .ZN(n87) );
  AND3_X2 U83 ( .A1(n117), .A2(n122), .A3(INSTR[2]), .ZN(n81) );
  NAND2_X2 U84 ( .A1(INSTR[5]), .A2(n121), .ZN(n105) );
  NOR4_X2 U85 ( .A1(n114), .A2(INSTR[0]), .A3(INSTR[3]), .A4(INSTR[2]), .ZN(
        n112) );
  NOR4_X2 U86 ( .A1(INSTR[6]), .A2(INSTR[4]), .A3(INSTR[10]), .A4(n115), .ZN(
        n113) );
  OR3_X4 U87 ( .A1(INSTR[9]), .A2(INSTR[8]), .A3(INSTR[7]), .ZN(n115) );
  NOR3_X2 U88 ( .A1(INSTR_28), .A2(INSTR_30), .A3(INSTR_29), .ZN(n116) );
  NAND2_X2 U89 ( .A1(n39), .A2(n41), .ZN(n67) );
  NAND3_X1 U118 ( .A1(n68), .A2(n39), .A3(INSTR_31), .ZN(n54) );
  NAND3_X1 U119 ( .A1(INSTR_29), .A2(n52), .A3(n45), .ZN(n71) );
  NAND3_X1 U120 ( .A1(INSTR_26), .A2(n80), .A3(INSTR_29), .ZN(n79) );
  OAI33_X1 U121 ( .A1(n121), .A2(INSTR[5]), .A3(n118), .B1(n122), .B2(INSTR[2]), .B3(n98), .ZN(n97) );
  NAND3_X1 U122 ( .A1(INSTR_26), .A2(n50), .A3(INSTR_27), .ZN(n77) );
  NAND3_X1 U123 ( .A1(INSTR_27), .A2(n44), .A3(INSTR_28), .ZN(n108) );
  NAND3_X1 U124 ( .A1(n96), .A2(n53), .A3(INSTR_30), .ZN(n110) );
  NAND3_X1 U125 ( .A1(n113), .A2(n120), .A3(INSTR[2]), .ZN(n104) );
  NAND3_X1 U126 ( .A1(n113), .A2(n119), .A3(INSTR[3]), .ZN(n98) );
  NAND3_X1 U127 ( .A1(n113), .A2(INSTR[5]), .A3(INSTR[1]), .ZN(n114) );
  NAND3_X1 U128 ( .A1(n38), .A2(INSTR_27), .A3(n116), .ZN(n55) );
  CLKBUF_X2 U90 ( .A(RST_AN), .Z(n26) );
  CLKBUF_X2 U91 ( .A(RST_AN), .Z(n27) );
  CLKBUF_X3 U92 ( .A(n26), .Z(n28) );
  CLKBUF_X3 U93 ( .A(n26), .Z(n29) );
  CLKBUF_X3 U94 ( .A(n27), .Z(n30) );
  CLKBUF_X3 U95 ( .A(n27), .Z(n31) );
  INV_X2 U96 ( .A(\HZRD_SIG[FLUSH_EM] ), .ZN(n32) );
  INV_X2 U97 ( .A(\HZRD_SIG[FLUSH_DE] ), .ZN(n33) );
  INV_X2 U98 ( .A(n54), .ZN(n34) );
  INV_X2 U99 ( .A(n101), .ZN(n35) );
  INV_X2 U100 ( .A(n55), .ZN(n36) );
  INV_X2 U101 ( .A(n64), .ZN(n37) );
  INV_X2 U102 ( .A(n67), .ZN(n38) );
  INV_X2 U103 ( .A(\HZRD_SIG[FLUSH_FD] ), .ZN(n39) );
  INV_X2 U104 ( .A(\HZRD_SIG[FLUSH_MWB] ), .ZN(n40) );
  INV_X2 U105 ( .A(INSTR_31), .ZN(n41) );
  INV_X2 U106 ( .A(n74), .ZN(n42) );
  INV_X2 U107 ( .A(n76), .ZN(n43) );
  INV_X2 U108 ( .A(INSTR_30), .ZN(n44) );
  INV_X2 U109 ( .A(n69), .ZN(n45) );
  INV_X2 U110 ( .A(n93), .ZN(n46) );
  INV_X2 U111 ( .A(n63), .ZN(n47) );
  INV_X2 U112 ( .A(n96), .ZN(n48) );
  INV_X2 U113 ( .A(INSTR_29), .ZN(n49) );
  INV_X2 U114 ( .A(INSTR_28), .ZN(n50) );
  INV_X2 U115 ( .A(n62), .ZN(n51) );
  INV_X2 U116 ( .A(INSTR_27), .ZN(n52) );
  INV_X2 U117 ( .A(INSTR_26), .ZN(n53) );
  INV_X2 U129 ( .A(n98), .ZN(n117) );
  INV_X2 U130 ( .A(n87), .ZN(n118) );
  INV_X2 U131 ( .A(n105), .ZN(n119) );
  INV_X2 U132 ( .A(INSTR[3]), .ZN(n120) );
  INV_X2 U133 ( .A(INSTR[1]), .ZN(n121) );
  INV_X2 U134 ( .A(INSTR[0]), .ZN(n122) );
endmodule


module REG_PIPO_32_fffffffc_fffffffc ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n97, n98, n99;

  DFFS_X1 \reg_mem_reg[31]  ( .D(n96), .CK(CLK), .SN(n21), .Q(DOUT[31]), .QN(
        n64) );
  DFFS_X1 \reg_mem_reg[30]  ( .D(n95), .CK(CLK), .SN(n21), .Q(DOUT[30]), .QN(
        n63) );
  DFFS_X1 \reg_mem_reg[29]  ( .D(n94), .CK(CLK), .SN(n21), .Q(DOUT[29]), .QN(
        n62) );
  DFFS_X1 \reg_mem_reg[28]  ( .D(n93), .CK(CLK), .SN(n21), .Q(DOUT[28]), .QN(
        n61) );
  DFFS_X1 \reg_mem_reg[27]  ( .D(n92), .CK(CLK), .SN(n21), .Q(DOUT[27]), .QN(
        n60) );
  DFFS_X1 \reg_mem_reg[26]  ( .D(n91), .CK(CLK), .SN(n21), .Q(DOUT[26]), .QN(
        n59) );
  DFFS_X1 \reg_mem_reg[25]  ( .D(n90), .CK(CLK), .SN(n20), .Q(DOUT[25]), .QN(
        n58) );
  DFFS_X1 \reg_mem_reg[24]  ( .D(n89), .CK(CLK), .SN(n20), .Q(DOUT[24]), .QN(
        n57) );
  DFFS_X1 \reg_mem_reg[23]  ( .D(n88), .CK(CLK), .SN(n20), .Q(DOUT[23]), .QN(
        n56) );
  DFFS_X1 \reg_mem_reg[22]  ( .D(n87), .CK(CLK), .SN(n20), .Q(DOUT[22]), .QN(
        n55) );
  DFFS_X1 \reg_mem_reg[21]  ( .D(n86), .CK(CLK), .SN(n20), .Q(DOUT[21]), .QN(
        n54) );
  DFFS_X1 \reg_mem_reg[20]  ( .D(n85), .CK(CLK), .SN(n20), .Q(DOUT[20]), .QN(
        n53) );
  DFFS_X1 \reg_mem_reg[19]  ( .D(n84), .CK(CLK), .SN(n20), .Q(DOUT[19]), .QN(
        n52) );
  DFFS_X1 \reg_mem_reg[18]  ( .D(n83), .CK(CLK), .SN(n20), .Q(DOUT[18]), .QN(
        n51) );
  DFFS_X1 \reg_mem_reg[17]  ( .D(n82), .CK(CLK), .SN(n20), .Q(DOUT[17]), .QN(
        n50) );
  DFFS_X1 \reg_mem_reg[16]  ( .D(n81), .CK(CLK), .SN(n20), .Q(DOUT[16]), .QN(
        n49) );
  DFFS_X1 \reg_mem_reg[15]  ( .D(n80), .CK(CLK), .SN(n20), .Q(DOUT[15]), .QN(
        n48) );
  DFFS_X1 \reg_mem_reg[14]  ( .D(n79), .CK(CLK), .SN(n20), .Q(DOUT[14]), .QN(
        n47) );
  DFFS_X1 \reg_mem_reg[13]  ( .D(n78), .CK(CLK), .SN(n20), .Q(DOUT[13]), .QN(
        n46) );
  DFFS_X1 \reg_mem_reg[12]  ( .D(n77), .CK(CLK), .SN(n19), .Q(DOUT[12]), .QN(
        n45) );
  DFFS_X1 \reg_mem_reg[11]  ( .D(n76), .CK(CLK), .SN(n19), .Q(DOUT[11]), .QN(
        n44) );
  DFFS_X1 \reg_mem_reg[10]  ( .D(n75), .CK(CLK), .SN(n19), .Q(DOUT[10]), .QN(
        n43) );
  DFFS_X1 \reg_mem_reg[9]  ( .D(n74), .CK(CLK), .SN(n19), .Q(DOUT[9]), .QN(n42) );
  DFFS_X1 \reg_mem_reg[8]  ( .D(n73), .CK(CLK), .SN(n19), .Q(DOUT[8]), .QN(n41) );
  DFFS_X1 \reg_mem_reg[7]  ( .D(n72), .CK(CLK), .SN(n19), .Q(DOUT[7]), .QN(n40) );
  DFFS_X1 \reg_mem_reg[6]  ( .D(n71), .CK(CLK), .SN(n19), .Q(DOUT[6]), .QN(n39) );
  DFFS_X1 \reg_mem_reg[5]  ( .D(n70), .CK(CLK), .SN(n19), .Q(DOUT[5]), .QN(n38) );
  DFFS_X1 \reg_mem_reg[4]  ( .D(n69), .CK(CLK), .SN(n19), .Q(DOUT[4]), .QN(n37) );
  DFFS_X1 \reg_mem_reg[3]  ( .D(n68), .CK(CLK), .SN(n19), .Q(DOUT[3]), .QN(n36) );
  DFFS_X1 \reg_mem_reg[2]  ( .D(n67), .CK(CLK), .SN(n19), .Q(DOUT[2]), .QN(n35) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n66), .CK(CLK), .RN(n19), .Q(DOUT[1]), .QN(n34) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n65), .CK(CLK), .RN(n19), .Q(DOUT[0]), .QN(n33) );
  OAI21_X2 U2 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X2 U3 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X2 U4 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X2 U5 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X2 U6 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X2 U7 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X2 U8 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X2 U9 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  OAI21_X2 U10 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  NAND2_X2 U11 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X2 U12 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  NAND2_X2 U13 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X2 U14 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X2 U15 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  OAI21_X2 U16 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  NAND2_X2 U17 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  OAI21_X2 U18 ( .B1(n41), .B2(EN), .A(n9), .ZN(n73) );
  NAND2_X2 U19 ( .A1(DIN[8]), .A2(EN), .ZN(n9) );
  OAI21_X2 U20 ( .B1(n42), .B2(EN), .A(n10), .ZN(n74) );
  NAND2_X2 U21 ( .A1(DIN[9]), .A2(EN), .ZN(n10) );
  OAI21_X2 U22 ( .B1(n43), .B2(EN), .A(n11), .ZN(n75) );
  NAND2_X2 U23 ( .A1(DIN[10]), .A2(EN), .ZN(n11) );
  OAI21_X2 U24 ( .B1(n44), .B2(EN), .A(n12), .ZN(n76) );
  NAND2_X2 U25 ( .A1(DIN[11]), .A2(EN), .ZN(n12) );
  OAI21_X2 U26 ( .B1(n45), .B2(EN), .A(n13), .ZN(n77) );
  NAND2_X2 U27 ( .A1(DIN[12]), .A2(EN), .ZN(n13) );
  OAI21_X2 U28 ( .B1(n46), .B2(EN), .A(n14), .ZN(n78) );
  NAND2_X2 U29 ( .A1(DIN[13]), .A2(EN), .ZN(n14) );
  OAI21_X2 U30 ( .B1(n47), .B2(EN), .A(n15), .ZN(n79) );
  NAND2_X2 U31 ( .A1(DIN[14]), .A2(EN), .ZN(n15) );
  OAI21_X2 U32 ( .B1(n48), .B2(EN), .A(n16), .ZN(n80) );
  NAND2_X2 U33 ( .A1(DIN[15]), .A2(EN), .ZN(n16) );
  OAI21_X2 U34 ( .B1(n49), .B2(EN), .A(n17), .ZN(n81) );
  NAND2_X2 U35 ( .A1(DIN[16]), .A2(EN), .ZN(n17) );
  OAI21_X2 U36 ( .B1(n50), .B2(EN), .A(n18), .ZN(n82) );
  NAND2_X2 U37 ( .A1(DIN[17]), .A2(EN), .ZN(n18) );
  OAI21_X2 U64 ( .B1(n64), .B2(EN), .A(n32), .ZN(n96) );
  NAND2_X2 U65 ( .A1(DIN[31]), .A2(EN), .ZN(n32) );
  CLKBUF_X3 U38 ( .A(RST_AN), .Z(n19) );
  CLKBUF_X3 U39 ( .A(RST_AN), .Z(n20) );
  CLKBUF_X3 U40 ( .A(RST_AN), .Z(n21) );
  INV_X1 U41 ( .A(n51), .ZN(n22) );
  MUX2_X1 U42 ( .A(n22), .B(DIN[18]), .S(EN), .Z(n83) );
  INV_X1 U43 ( .A(n52), .ZN(n23) );
  MUX2_X1 U44 ( .A(n23), .B(DIN[19]), .S(EN), .Z(n84) );
  INV_X1 U45 ( .A(n53), .ZN(n24) );
  MUX2_X1 U46 ( .A(n24), .B(DIN[20]), .S(EN), .Z(n85) );
  INV_X1 U47 ( .A(n54), .ZN(n25) );
  MUX2_X1 U48 ( .A(n25), .B(DIN[21]), .S(EN), .Z(n86) );
  INV_X1 U49 ( .A(n55), .ZN(n26) );
  MUX2_X1 U50 ( .A(n26), .B(DIN[22]), .S(EN), .Z(n87) );
  INV_X1 U51 ( .A(n56), .ZN(n27) );
  MUX2_X1 U52 ( .A(n27), .B(DIN[23]), .S(EN), .Z(n88) );
  INV_X1 U53 ( .A(n57), .ZN(n28) );
  MUX2_X1 U54 ( .A(n28), .B(DIN[24]), .S(EN), .Z(n89) );
  INV_X1 U55 ( .A(n58), .ZN(n29) );
  MUX2_X1 U56 ( .A(n29), .B(DIN[25]), .S(EN), .Z(n90) );
  INV_X1 U57 ( .A(n59), .ZN(n30) );
  MUX2_X1 U58 ( .A(n30), .B(DIN[26]), .S(EN), .Z(n91) );
  INV_X1 U59 ( .A(n60), .ZN(n31) );
  MUX2_X1 U60 ( .A(n31), .B(DIN[27]), .S(EN), .Z(n92) );
  INV_X1 U61 ( .A(n61), .ZN(n97) );
  MUX2_X1 U62 ( .A(n97), .B(DIN[28]), .S(EN), .Z(n93) );
  INV_X1 U63 ( .A(n62), .ZN(n98) );
  MUX2_X1 U66 ( .A(n98), .B(DIN[29]), .S(EN), .Z(n94) );
  INV_X1 U67 ( .A(n63), .ZN(n99) );
  MUX2_X1 U68 ( .A(n99), .B(DIN[30]), .S(EN), .Z(n95) );
endmodule


module REG_PIPO_32_00000000_00000000_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n99,
         n100, n101, n102;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n98), .CK(CLK), .RN(n4), .Q(DOUT[31]), .QN(
        n66) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n97), .CK(CLK), .RN(n4), .Q(DOUT[30]), .QN(
        n65) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n96), .CK(CLK), .RN(n4), .Q(DOUT[29]), .QN(
        n64) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n95), .CK(CLK), .RN(n4), .Q(DOUT[28]), .QN(
        n63) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n94), .CK(CLK), .RN(n4), .Q(DOUT[27]), .QN(
        n62) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n93), .CK(CLK), .RN(n4), .Q(DOUT[26]), .QN(
        n61) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n92), .CK(CLK), .RN(n4), .Q(DOUT[25]), .QN(
        n60) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n91), .CK(CLK), .RN(n4), .Q(DOUT[24]), .QN(
        n59) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n90), .CK(CLK), .RN(n4), .Q(DOUT[23]), .QN(
        n58) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n89), .CK(CLK), .RN(n4), .Q(DOUT[22]), .QN(
        n57) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n88), .CK(CLK), .RN(n3), .Q(DOUT[21]), .QN(
        n56) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n87), .CK(CLK), .RN(n3), .Q(DOUT[20]), .QN(
        n55) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n86), .CK(CLK), .RN(n3), .Q(DOUT[19]), .QN(
        n54) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n85), .CK(CLK), .RN(n3), .Q(DOUT[18]), .QN(
        n53) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n84), .CK(CLK), .RN(n3), .Q(DOUT[17]), .QN(
        n52) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n83), .CK(CLK), .RN(n3), .Q(DOUT[16]), .QN(
        n51) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n82), .CK(CLK), .RN(n3), .Q(DOUT[15]), .QN(
        n50) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n81), .CK(CLK), .RN(n3), .Q(DOUT[14]), .QN(
        n49) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n80), .CK(CLK), .RN(n3), .Q(DOUT[13]), .QN(
        n48) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n79), .CK(CLK), .RN(n3), .Q(DOUT[12]), .QN(
        n47) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n78), .CK(CLK), .RN(n3), .Q(DOUT[11]), .QN(
        n46) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n77), .CK(CLK), .RN(n2), .Q(DOUT[10]), .QN(
        n45) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n76), .CK(CLK), .RN(n2), .Q(DOUT[9]), .QN(n44)
         );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n75), .CK(CLK), .RN(n2), .Q(DOUT[8]), .QN(n43)
         );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n74), .CK(CLK), .RN(n2), .Q(DOUT[7]), .QN(n42)
         );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n73), .CK(CLK), .RN(n2), .Q(DOUT[6]), .QN(n41)
         );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n72), .CK(CLK), .RN(n2), .Q(DOUT[5]), .QN(n40)
         );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n71), .CK(CLK), .RN(n2), .Q(DOUT[4]), .QN(n39)
         );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n70), .CK(CLK), .RN(n2), .Q(DOUT[3]), .QN(n38)
         );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n69), .CK(CLK), .RN(n2), .Q(DOUT[2]), .QN(n37)
         );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n68), .CK(CLK), .RN(n2), .Q(DOUT[1]), .QN(n36)
         );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n67), .CK(CLK), .RN(n2), .Q(DOUT[0]), .QN(n35)
         );
  OAI22_X2 U2 ( .A1(n35), .A2(EN), .B1(n1), .B2(n101), .ZN(n67) );
  OAI22_X2 U4 ( .A1(n36), .A2(EN), .B1(n1), .B2(n100), .ZN(n68) );
  OAI22_X2 U6 ( .A1(n37), .A2(EN), .B1(n1), .B2(n99), .ZN(n69) );
  OAI22_X2 U8 ( .A1(n38), .A2(EN), .B1(n1), .B2(n34), .ZN(n70) );
  OAI22_X2 U10 ( .A1(n39), .A2(EN), .B1(n1), .B2(n33), .ZN(n71) );
  OAI22_X2 U12 ( .A1(n40), .A2(EN), .B1(n1), .B2(n32), .ZN(n72) );
  OAI22_X2 U14 ( .A1(n41), .A2(EN), .B1(n1), .B2(n31), .ZN(n73) );
  OAI22_X2 U16 ( .A1(n42), .A2(EN), .B1(n1), .B2(n30), .ZN(n74) );
  OAI22_X2 U18 ( .A1(n43), .A2(EN), .B1(n1), .B2(n29), .ZN(n75) );
  OAI22_X2 U20 ( .A1(n44), .A2(EN), .B1(n1), .B2(n28), .ZN(n76) );
  OAI22_X2 U22 ( .A1(n45), .A2(EN), .B1(n1), .B2(n27), .ZN(n77) );
  OAI22_X2 U24 ( .A1(n46), .A2(EN), .B1(n1), .B2(n26), .ZN(n78) );
  OAI22_X2 U26 ( .A1(n47), .A2(EN), .B1(n1), .B2(n25), .ZN(n79) );
  OAI22_X2 U28 ( .A1(n48), .A2(EN), .B1(n1), .B2(n24), .ZN(n80) );
  OAI22_X2 U30 ( .A1(n49), .A2(EN), .B1(n1), .B2(n23), .ZN(n81) );
  OAI22_X2 U32 ( .A1(n50), .A2(EN), .B1(n1), .B2(n22), .ZN(n82) );
  OAI22_X2 U34 ( .A1(n51), .A2(EN), .B1(n1), .B2(n21), .ZN(n83) );
  OAI22_X2 U36 ( .A1(n52), .A2(EN), .B1(n1), .B2(n20), .ZN(n84) );
  OAI22_X2 U64 ( .A1(n66), .A2(EN), .B1(n1), .B2(n102), .ZN(n98) );
  CLKBUF_X3 U3 ( .A(RST_AN), .Z(n2) );
  CLKBUF_X3 U5 ( .A(RST_AN), .Z(n3) );
  CLKBUF_X3 U7 ( .A(RST_AN), .Z(n4) );
  INV_X1 U9 ( .A(EN), .ZN(n5) );
  OR2_X1 U11 ( .A1(INIT), .A2(n5), .ZN(n1) );
  INV_X1 U13 ( .A(n1), .ZN(n18) );
  NAND2_X1 U15 ( .A1(DIN[18]), .A2(n18), .ZN(n6) );
  OAI21_X1 U17 ( .B1(n53), .B2(EN), .A(n6), .ZN(n85) );
  NAND2_X1 U19 ( .A1(DIN[19]), .A2(n18), .ZN(n7) );
  OAI21_X1 U21 ( .B1(n54), .B2(EN), .A(n7), .ZN(n86) );
  NAND2_X1 U23 ( .A1(DIN[20]), .A2(n18), .ZN(n8) );
  OAI21_X1 U25 ( .B1(n55), .B2(EN), .A(n8), .ZN(n87) );
  NAND2_X1 U27 ( .A1(DIN[21]), .A2(n18), .ZN(n9) );
  OAI21_X1 U29 ( .B1(n56), .B2(EN), .A(n9), .ZN(n88) );
  NAND2_X1 U31 ( .A1(DIN[22]), .A2(n18), .ZN(n10) );
  OAI21_X1 U33 ( .B1(n57), .B2(EN), .A(n10), .ZN(n89) );
  NAND2_X1 U35 ( .A1(DIN[23]), .A2(n18), .ZN(n11) );
  OAI21_X1 U37 ( .B1(n58), .B2(EN), .A(n11), .ZN(n90) );
  NAND2_X1 U38 ( .A1(DIN[24]), .A2(n18), .ZN(n12) );
  OAI21_X1 U39 ( .B1(n59), .B2(EN), .A(n12), .ZN(n91) );
  NAND2_X1 U40 ( .A1(DIN[25]), .A2(n18), .ZN(n13) );
  OAI21_X1 U41 ( .B1(n60), .B2(EN), .A(n13), .ZN(n92) );
  NAND2_X1 U42 ( .A1(DIN[26]), .A2(n18), .ZN(n14) );
  OAI21_X1 U43 ( .B1(n61), .B2(EN), .A(n14), .ZN(n93) );
  NAND2_X1 U44 ( .A1(DIN[27]), .A2(n18), .ZN(n15) );
  OAI21_X1 U45 ( .B1(n62), .B2(EN), .A(n15), .ZN(n94) );
  NAND2_X1 U46 ( .A1(DIN[28]), .A2(n18), .ZN(n16) );
  OAI21_X1 U47 ( .B1(n63), .B2(EN), .A(n16), .ZN(n95) );
  NAND2_X1 U48 ( .A1(DIN[29]), .A2(n18), .ZN(n17) );
  OAI21_X1 U49 ( .B1(n64), .B2(EN), .A(n17), .ZN(n96) );
  NAND2_X1 U50 ( .A1(DIN[30]), .A2(n18), .ZN(n19) );
  OAI21_X1 U51 ( .B1(n65), .B2(EN), .A(n19), .ZN(n97) );
  INV_X2 U52 ( .A(DIN[17]), .ZN(n20) );
  INV_X2 U53 ( .A(DIN[16]), .ZN(n21) );
  INV_X2 U54 ( .A(DIN[15]), .ZN(n22) );
  INV_X2 U55 ( .A(DIN[14]), .ZN(n23) );
  INV_X2 U56 ( .A(DIN[13]), .ZN(n24) );
  INV_X2 U57 ( .A(DIN[12]), .ZN(n25) );
  INV_X2 U58 ( .A(DIN[11]), .ZN(n26) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n27) );
  INV_X2 U60 ( .A(DIN[9]), .ZN(n28) );
  INV_X2 U61 ( .A(DIN[8]), .ZN(n29) );
  INV_X2 U62 ( .A(DIN[7]), .ZN(n30) );
  INV_X2 U63 ( .A(DIN[6]), .ZN(n31) );
  INV_X2 U65 ( .A(DIN[5]), .ZN(n32) );
  INV_X2 U66 ( .A(DIN[4]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[3]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[2]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[1]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[0]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[31]), .ZN(n102) );
endmodule


module REG_PIPO_32_00000000_00000000_11 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module RF_ADDR_W5_DATA_W32 ( CLK, RST_AN, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST_AN, ENABLE, RD1, RD2, WR;
  wire   \registers[1][31] , \registers[1][30] , \registers[1][29] ,
         \registers[1][28] , \registers[1][27] , \registers[1][26] ,
         \registers[1][25] , \registers[1][24] , \registers[1][23] ,
         \registers[1][22] , \registers[1][21] , \registers[1][20] ,
         \registers[1][19] , \registers[1][18] , \registers[1][17] ,
         \registers[1][16] , \registers[1][15] , \registers[1][14] ,
         \registers[1][13] , \registers[1][12] , \registers[1][11] ,
         \registers[1][10] , \registers[1][9] , \registers[1][8] ,
         \registers[1][7] , \registers[1][6] , \registers[1][5] ,
         \registers[1][4] , \registers[1][3] , \registers[1][2] ,
         \registers[1][1] , \registers[1][0] , \registers[6][31] ,
         \registers[6][30] , \registers[6][29] , \registers[6][28] ,
         \registers[6][27] , \registers[6][26] , \registers[6][25] ,
         \registers[6][24] , \registers[6][23] , \registers[6][22] ,
         \registers[6][21] , \registers[6][20] , \registers[6][19] ,
         \registers[6][18] , \registers[6][17] , \registers[6][16] ,
         \registers[6][15] , \registers[6][14] , \registers[6][13] ,
         \registers[6][12] , \registers[6][11] , \registers[6][10] ,
         \registers[6][9] , \registers[6][8] , \registers[6][7] ,
         \registers[6][6] , \registers[6][5] , \registers[6][4] ,
         \registers[6][3] , \registers[6][2] , \registers[6][1] ,
         \registers[6][0] , \registers[7][31] , \registers[7][30] ,
         \registers[7][29] , \registers[7][28] , \registers[7][27] ,
         \registers[7][26] , \registers[7][25] , \registers[7][24] ,
         \registers[7][23] , \registers[7][22] , \registers[7][21] ,
         \registers[7][20] , \registers[7][19] , \registers[7][18] ,
         \registers[7][17] , \registers[7][16] , \registers[7][15] ,
         \registers[7][14] , \registers[7][13] , \registers[7][12] ,
         \registers[7][11] , \registers[7][10] , \registers[7][9] ,
         \registers[7][8] , \registers[7][7] , \registers[7][6] ,
         \registers[7][5] , \registers[7][4] , \registers[7][3] ,
         \registers[7][2] , \registers[7][1] , \registers[7][0] ,
         \registers[8][31] , \registers[8][30] , \registers[8][29] ,
         \registers[8][28] , \registers[8][27] , \registers[8][26] ,
         \registers[8][25] , \registers[8][24] , \registers[8][23] ,
         \registers[8][22] , \registers[8][21] , \registers[8][20] ,
         \registers[8][19] , \registers[8][18] , \registers[8][17] ,
         \registers[8][16] , \registers[8][15] , \registers[8][14] ,
         \registers[8][13] , \registers[8][12] , \registers[8][11] ,
         \registers[8][10] , \registers[8][9] , \registers[8][8] ,
         \registers[8][7] , \registers[8][6] , \registers[8][5] ,
         \registers[8][4] , \registers[8][3] , \registers[8][2] ,
         \registers[8][1] , \registers[8][0] , \registers[9][31] ,
         \registers[9][30] , \registers[9][29] , \registers[9][28] ,
         \registers[9][27] , \registers[9][26] , \registers[9][25] ,
         \registers[9][24] , \registers[9][23] , \registers[9][22] ,
         \registers[9][21] , \registers[9][20] , \registers[9][19] ,
         \registers[9][18] , \registers[9][17] , \registers[9][16] ,
         \registers[9][15] , \registers[9][14] , \registers[9][13] ,
         \registers[9][12] , \registers[9][11] , \registers[9][10] ,
         \registers[9][9] , \registers[9][8] , \registers[9][7] ,
         \registers[9][6] , \registers[9][5] , \registers[9][4] ,
         \registers[9][3] , \registers[9][2] , \registers[9][1] ,
         \registers[9][0] , \registers[12][31] , \registers[12][30] ,
         \registers[12][29] , \registers[12][28] , \registers[12][27] ,
         \registers[12][26] , \registers[12][25] , \registers[12][24] ,
         \registers[12][23] , \registers[12][22] , \registers[12][21] ,
         \registers[12][20] , \registers[12][19] , \registers[12][18] ,
         \registers[12][17] , \registers[12][16] , \registers[12][15] ,
         \registers[12][14] , \registers[12][13] , \registers[12][12] ,
         \registers[12][11] , \registers[12][10] , \registers[12][9] ,
         \registers[12][8] , \registers[12][7] , \registers[12][6] ,
         \registers[12][5] , \registers[12][4] , \registers[12][3] ,
         \registers[12][2] , \registers[12][1] , \registers[12][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[18][31] ,
         \registers[18][30] , \registers[18][29] , \registers[18][28] ,
         \registers[18][27] , \registers[18][26] , \registers[18][25] ,
         \registers[18][24] , \registers[18][23] , \registers[18][22] ,
         \registers[18][21] , \registers[18][20] , \registers[18][19] ,
         \registers[18][18] , \registers[18][17] , \registers[18][16] ,
         \registers[18][15] , \registers[18][14] , \registers[18][13] ,
         \registers[18][12] , \registers[18][11] , \registers[18][10] ,
         \registers[18][9] , \registers[18][8] , \registers[18][7] ,
         \registers[18][6] , \registers[18][5] , \registers[18][4] ,
         \registers[18][3] , \registers[18][2] , \registers[18][1] ,
         \registers[18][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[22][31] , \registers[22][30] , \registers[22][29] ,
         \registers[22][28] , \registers[22][27] , \registers[22][26] ,
         \registers[22][25] , \registers[22][24] , \registers[22][23] ,
         \registers[22][22] , \registers[22][21] , \registers[22][20] ,
         \registers[22][19] , \registers[22][18] , \registers[22][17] ,
         \registers[22][16] , \registers[22][15] , \registers[22][14] ,
         \registers[22][13] , \registers[22][12] , \registers[22][11] ,
         \registers[22][10] , \registers[22][9] , \registers[22][8] ,
         \registers[22][7] , \registers[22][6] , \registers[22][5] ,
         \registers[22][4] , \registers[22][3] , \registers[22][2] ,
         \registers[22][1] , \registers[22][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[24][31] , \registers[24][30] ,
         \registers[24][29] , \registers[24][28] , \registers[24][27] ,
         \registers[24][26] , \registers[24][25] , \registers[24][24] ,
         \registers[24][23] , \registers[24][22] , \registers[24][21] ,
         \registers[24][20] , \registers[24][19] , \registers[24][18] ,
         \registers[24][17] , \registers[24][16] , \registers[24][15] ,
         \registers[24][14] , \registers[24][13] , \registers[24][12] ,
         \registers[24][11] , \registers[24][10] , \registers[24][9] ,
         \registers[24][8] , \registers[24][7] , \registers[24][6] ,
         \registers[24][5] , \registers[24][4] , \registers[24][3] ,
         \registers[24][2] , \registers[24][1] , \registers[24][0] ,
         \registers[25][31] , \registers[25][30] , \registers[25][29] ,
         \registers[25][28] , \registers[25][27] , \registers[25][26] ,
         \registers[25][25] , \registers[25][24] , \registers[25][23] ,
         \registers[25][22] , \registers[25][21] , \registers[25][20] ,
         \registers[25][19] , \registers[25][18] , \registers[25][17] ,
         \registers[25][16] , \registers[25][15] , \registers[25][14] ,
         \registers[25][13] , \registers[25][12] , \registers[25][11] ,
         \registers[25][10] , \registers[25][9] , \registers[25][8] ,
         \registers[25][7] , \registers[25][6] , \registers[25][5] ,
         \registers[25][4] , \registers[25][3] , \registers[25][2] ,
         \registers[25][1] , \registers[25][0] , \registers[28][31] ,
         \registers[28][30] , \registers[28][29] , \registers[28][28] ,
         \registers[28][27] , \registers[28][26] , \registers[28][25] ,
         \registers[28][24] , \registers[28][23] , \registers[28][22] ,
         \registers[28][21] , \registers[28][20] , \registers[28][19] ,
         \registers[28][18] , \registers[28][17] , \registers[28][16] ,
         \registers[28][15] , \registers[28][14] , \registers[28][13] ,
         \registers[28][12] , \registers[28][11] , \registers[28][10] ,
         \registers[28][9] , \registers[28][8] , \registers[28][7] ,
         \registers[28][6] , \registers[28][5] , \registers[28][4] ,
         \registers[28][3] , \registers[28][2] , \registers[28][1] ,
         \registers[28][0] , \registers[29][31] , \registers[29][30] ,
         \registers[29][29] , \registers[29][28] , \registers[29][27] ,
         \registers[29][26] , \registers[29][25] , \registers[29][24] ,
         \registers[29][23] , \registers[29][22] , \registers[29][21] ,
         \registers[29][20] , \registers[29][19] , \registers[29][18] ,
         \registers[29][17] , \registers[29][16] , \registers[29][15] ,
         \registers[29][14] , \registers[29][13] , \registers[29][12] ,
         \registers[29][11] , \registers[29][10] , \registers[29][9] ,
         \registers[29][8] , \registers[29][7] , \registers[29][6] ,
         \registers[29][5] , \registers[29][4] , \registers[29][3] ,
         \registers[29][2] , \registers[29][1] , \registers[29][0] , N83, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891;

  DFFR_X1 \registers_reg[1][31]  ( .D(n3527), .CK(n3891), .RN(n3351), .Q(
        \registers[1][31] ) );
  DFFR_X1 \registers_reg[1][30]  ( .D(n3526), .CK(n3891), .RN(n3351), .Q(
        \registers[1][30] ) );
  DFFR_X1 \registers_reg[1][29]  ( .D(n3525), .CK(n3891), .RN(n3350), .Q(
        \registers[1][29] ) );
  DFFR_X1 \registers_reg[1][28]  ( .D(n3524), .CK(n3891), .RN(n3350), .Q(
        \registers[1][28] ) );
  DFFR_X1 \registers_reg[1][27]  ( .D(n3523), .CK(n3891), .RN(n3350), .Q(
        \registers[1][27] ) );
  DFFR_X1 \registers_reg[1][26]  ( .D(n3522), .CK(n3891), .RN(n3350), .Q(
        \registers[1][26] ) );
  DFFR_X1 \registers_reg[1][25]  ( .D(n3521), .CK(n3891), .RN(n3350), .Q(
        \registers[1][25] ) );
  DFFR_X1 \registers_reg[1][24]  ( .D(n3520), .CK(n3891), .RN(n3350), .Q(
        \registers[1][24] ) );
  DFFR_X1 \registers_reg[1][23]  ( .D(n3519), .CK(n3891), .RN(n3350), .Q(
        \registers[1][23] ) );
  DFFR_X1 \registers_reg[1][22]  ( .D(n3518), .CK(n3891), .RN(n3350), .Q(
        \registers[1][22] ) );
  DFFR_X1 \registers_reg[1][21]  ( .D(n3517), .CK(n3891), .RN(n3350), .Q(
        \registers[1][21] ) );
  DFFR_X1 \registers_reg[1][20]  ( .D(n3516), .CK(n3891), .RN(n3350), .Q(
        \registers[1][20] ) );
  DFFR_X1 \registers_reg[1][19]  ( .D(n3515), .CK(n3891), .RN(n3350), .Q(
        \registers[1][19] ) );
  DFFR_X1 \registers_reg[1][18]  ( .D(n3514), .CK(n3891), .RN(n3349), .Q(
        \registers[1][18] ) );
  DFFR_X1 \registers_reg[1][17]  ( .D(n3513), .CK(n3891), .RN(n3349), .Q(
        \registers[1][17] ) );
  DFFR_X1 \registers_reg[1][16]  ( .D(n3512), .CK(n3891), .RN(n3349), .Q(
        \registers[1][16] ) );
  DFFR_X1 \registers_reg[1][15]  ( .D(n3511), .CK(n3891), .RN(n3349), .Q(
        \registers[1][15] ) );
  DFFR_X1 \registers_reg[1][14]  ( .D(n3510), .CK(n3891), .RN(n3349), .Q(
        \registers[1][14] ) );
  DFFR_X1 \registers_reg[1][13]  ( .D(n3509), .CK(n3891), .RN(n3349), .Q(
        \registers[1][13] ) );
  DFFR_X1 \registers_reg[1][12]  ( .D(n3508), .CK(n3891), .RN(n3349), .Q(
        \registers[1][12] ) );
  DFFR_X1 \registers_reg[1][11]  ( .D(n3507), .CK(n3891), .RN(n3349), .Q(
        \registers[1][11] ) );
  DFFR_X1 \registers_reg[1][10]  ( .D(n3506), .CK(n3891), .RN(n3349), .Q(
        \registers[1][10] ) );
  DFFR_X1 \registers_reg[1][9]  ( .D(n3505), .CK(n3891), .RN(n3349), .Q(
        \registers[1][9] ) );
  DFFR_X1 \registers_reg[1][8]  ( .D(n3504), .CK(n3891), .RN(n3349), .Q(
        \registers[1][8] ) );
  DFFR_X1 \registers_reg[1][7]  ( .D(n3503), .CK(n3891), .RN(n3348), .Q(
        \registers[1][7] ) );
  DFFR_X1 \registers_reg[1][6]  ( .D(n3502), .CK(n3891), .RN(n3348), .Q(
        \registers[1][6] ) );
  DFFR_X1 \registers_reg[1][5]  ( .D(n3501), .CK(n3891), .RN(n3348), .Q(
        \registers[1][5] ) );
  DFFR_X1 \registers_reg[1][4]  ( .D(n3500), .CK(n3891), .RN(n3348), .Q(
        \registers[1][4] ) );
  DFFR_X1 \registers_reg[1][3]  ( .D(n3499), .CK(n3891), .RN(n3348), .Q(
        \registers[1][3] ) );
  DFFR_X1 \registers_reg[1][2]  ( .D(n3498), .CK(n3891), .RN(n3348), .Q(
        \registers[1][2] ) );
  DFFR_X1 \registers_reg[1][1]  ( .D(n3497), .CK(n3891), .RN(n3348), .Q(
        \registers[1][1] ) );
  DFFR_X1 \registers_reg[1][0]  ( .D(n3496), .CK(n3891), .RN(n3348), .Q(
        \registers[1][0] ) );
  DFFR_X1 \registers_reg[2][31]  ( .D(n3285), .CK(n3891), .RN(n3348), .QN(n33)
         );
  DFFR_X1 \registers_reg[2][30]  ( .D(n3284), .CK(n3891), .RN(n3348), .QN(n34)
         );
  DFFR_X1 \registers_reg[2][29]  ( .D(n3283), .CK(n3891), .RN(n3348), .QN(n35)
         );
  DFFR_X1 \registers_reg[2][28]  ( .D(n3282), .CK(n3891), .RN(n3347), .QN(n36)
         );
  DFFR_X1 \registers_reg[2][27]  ( .D(n3281), .CK(n3891), .RN(n3347), .QN(n37)
         );
  DFFR_X1 \registers_reg[2][26]  ( .D(n3280), .CK(n3891), .RN(n3347), .QN(n38)
         );
  DFFR_X1 \registers_reg[2][25]  ( .D(n3279), .CK(n3891), .RN(n3347), .QN(n39)
         );
  DFFR_X1 \registers_reg[2][24]  ( .D(n3278), .CK(n3891), .RN(n3347), .QN(n40)
         );
  DFFR_X1 \registers_reg[2][23]  ( .D(n3277), .CK(n3891), .RN(n3347), .QN(n41)
         );
  DFFR_X1 \registers_reg[2][22]  ( .D(n3276), .CK(n3891), .RN(n3347), .QN(n42)
         );
  DFFR_X1 \registers_reg[2][21]  ( .D(n3275), .CK(n3891), .RN(n3347), .QN(n43)
         );
  DFFR_X1 \registers_reg[2][20]  ( .D(n3274), .CK(n3891), .RN(n3347), .QN(n44)
         );
  DFFR_X1 \registers_reg[2][19]  ( .D(n3273), .CK(n3891), .RN(n3347), .QN(n45)
         );
  DFFR_X1 \registers_reg[2][18]  ( .D(n3272), .CK(n3891), .RN(n3347), .QN(n46)
         );
  DFFR_X1 \registers_reg[2][17]  ( .D(n3271), .CK(n3891), .RN(n3346), .QN(n47)
         );
  DFFR_X1 \registers_reg[2][16]  ( .D(n3270), .CK(n3891), .RN(n3346), .QN(n48)
         );
  DFFR_X1 \registers_reg[2][15]  ( .D(n3269), .CK(n3891), .RN(n3346), .QN(n49)
         );
  DFFR_X1 \registers_reg[2][14]  ( .D(n3268), .CK(n3891), .RN(n3346), .QN(n50)
         );
  DFFR_X1 \registers_reg[2][13]  ( .D(n3267), .CK(n3891), .RN(n3346), .QN(n51)
         );
  DFFR_X1 \registers_reg[2][12]  ( .D(n3266), .CK(n3891), .RN(n3346), .QN(n52)
         );
  DFFR_X1 \registers_reg[2][11]  ( .D(n3265), .CK(n3891), .RN(n3346), .QN(n53)
         );
  DFFR_X1 \registers_reg[2][10]  ( .D(n3264), .CK(n3891), .RN(n3346), .QN(n54)
         );
  DFFR_X1 \registers_reg[2][9]  ( .D(n3263), .CK(n3891), .RN(n3346), .QN(n55)
         );
  DFFR_X1 \registers_reg[2][8]  ( .D(n3262), .CK(n3891), .RN(n3346), .QN(n56)
         );
  DFFR_X1 \registers_reg[2][7]  ( .D(n3261), .CK(n3891), .RN(n3346), .QN(n57)
         );
  DFFR_X1 \registers_reg[2][6]  ( .D(n3260), .CK(n3891), .RN(n3345), .QN(n58)
         );
  DFFR_X1 \registers_reg[2][5]  ( .D(n3259), .CK(n3891), .RN(n3345), .QN(n59)
         );
  DFFR_X1 \registers_reg[2][4]  ( .D(n3258), .CK(n3891), .RN(n3345), .QN(n60)
         );
  DFFR_X1 \registers_reg[2][3]  ( .D(n3257), .CK(n3891), .RN(n3345), .QN(n61)
         );
  DFFR_X1 \registers_reg[2][2]  ( .D(n3256), .CK(n3891), .RN(n3345), .QN(n62)
         );
  DFFR_X1 \registers_reg[2][1]  ( .D(n3255), .CK(n3891), .RN(n3345), .QN(n63)
         );
  DFFR_X1 \registers_reg[2][0]  ( .D(n3254), .CK(n3891), .RN(n3345), .QN(n64)
         );
  DFFR_X1 \registers_reg[3][31]  ( .D(n3253), .CK(n3891), .RN(n3345), .QN(n65)
         );
  DFFR_X1 \registers_reg[3][30]  ( .D(n3252), .CK(n3891), .RN(n3345), .QN(n66)
         );
  DFFR_X1 \registers_reg[3][29]  ( .D(n3251), .CK(n3891), .RN(n3345), .QN(n67)
         );
  DFFR_X1 \registers_reg[3][28]  ( .D(n3250), .CK(n3891), .RN(n3345), .QN(n68)
         );
  DFFR_X1 \registers_reg[3][27]  ( .D(n3249), .CK(n3891), .RN(n3344), .QN(n69)
         );
  DFFR_X1 \registers_reg[3][26]  ( .D(n3248), .CK(n3891), .RN(n3344), .QN(n70)
         );
  DFFR_X1 \registers_reg[3][25]  ( .D(n3247), .CK(n3891), .RN(n3344), .QN(n71)
         );
  DFFR_X1 \registers_reg[3][24]  ( .D(n3246), .CK(n3891), .RN(n3344), .QN(n72)
         );
  DFFR_X1 \registers_reg[3][23]  ( .D(n3245), .CK(n3891), .RN(n3344), .QN(n73)
         );
  DFFR_X1 \registers_reg[3][22]  ( .D(n3244), .CK(n3891), .RN(n3344), .QN(n74)
         );
  DFFR_X1 \registers_reg[3][21]  ( .D(n3243), .CK(n3891), .RN(n3344), .QN(n75)
         );
  DFFR_X1 \registers_reg[3][20]  ( .D(n3242), .CK(n3891), .RN(n3344), .QN(n76)
         );
  DFFR_X1 \registers_reg[3][19]  ( .D(n3241), .CK(n3891), .RN(n3344), .QN(n77)
         );
  DFFR_X1 \registers_reg[3][18]  ( .D(n3240), .CK(n3891), .RN(n3344), .QN(n78)
         );
  DFFR_X1 \registers_reg[3][17]  ( .D(n3239), .CK(n3891), .RN(n3344), .QN(n79)
         );
  DFFR_X1 \registers_reg[3][16]  ( .D(n3238), .CK(n3891), .RN(n3343), .QN(n80)
         );
  DFFR_X1 \registers_reg[3][15]  ( .D(n3237), .CK(n3891), .RN(n3343), .QN(n81)
         );
  DFFR_X1 \registers_reg[3][14]  ( .D(n3236), .CK(n3891), .RN(n3343), .QN(n82)
         );
  DFFR_X1 \registers_reg[3][13]  ( .D(n3235), .CK(n3891), .RN(n3343), .QN(n83)
         );
  DFFR_X1 \registers_reg[3][12]  ( .D(n3234), .CK(n3891), .RN(n3343), .QN(n84)
         );
  DFFR_X1 \registers_reg[3][11]  ( .D(n3233), .CK(n3891), .RN(n3343), .QN(n85)
         );
  DFFR_X1 \registers_reg[3][10]  ( .D(n3232), .CK(n3891), .RN(n3343), .QN(n86)
         );
  DFFR_X1 \registers_reg[3][9]  ( .D(n3231), .CK(n3891), .RN(n3343), .QN(n87)
         );
  DFFR_X1 \registers_reg[3][8]  ( .D(n3230), .CK(n3891), .RN(n3343), .QN(n88)
         );
  DFFR_X1 \registers_reg[3][7]  ( .D(n3229), .CK(n3891), .RN(n3343), .QN(n89)
         );
  DFFR_X1 \registers_reg[3][6]  ( .D(n3228), .CK(n3891), .RN(n3343), .QN(n90)
         );
  DFFR_X1 \registers_reg[3][5]  ( .D(n3227), .CK(n3891), .RN(n3342), .QN(n91)
         );
  DFFR_X1 \registers_reg[3][4]  ( .D(n3226), .CK(n3891), .RN(n3342), .QN(n92)
         );
  DFFR_X1 \registers_reg[3][3]  ( .D(n3225), .CK(n3891), .RN(n3342), .QN(n93)
         );
  DFFR_X1 \registers_reg[3][2]  ( .D(n3224), .CK(n3891), .RN(n3342), .QN(n94)
         );
  DFFR_X1 \registers_reg[3][1]  ( .D(n3223), .CK(n3891), .RN(n3342), .QN(n95)
         );
  DFFR_X1 \registers_reg[3][0]  ( .D(n3222), .CK(n3891), .RN(n3342), .QN(n96)
         );
  DFFR_X1 \registers_reg[4][31]  ( .D(n3221), .CK(n3891), .RN(n3342), .QN(n97)
         );
  DFFR_X1 \registers_reg[4][30]  ( .D(n3220), .CK(n3891), .RN(n3342), .QN(n98)
         );
  DFFR_X1 \registers_reg[4][29]  ( .D(n3219), .CK(n3891), .RN(n3342), .QN(n99)
         );
  DFFR_X1 \registers_reg[4][28]  ( .D(n3218), .CK(n3891), .RN(n3342), .QN(n100) );
  DFFR_X1 \registers_reg[4][27]  ( .D(n3217), .CK(n3891), .RN(n3342), .QN(n101) );
  DFFR_X1 \registers_reg[4][26]  ( .D(n3216), .CK(n3891), .RN(n3341), .QN(n102) );
  DFFR_X1 \registers_reg[4][25]  ( .D(n3215), .CK(n3891), .RN(n3341), .QN(n103) );
  DFFR_X1 \registers_reg[4][24]  ( .D(n3214), .CK(n3891), .RN(n3341), .QN(n104) );
  DFFR_X1 \registers_reg[4][23]  ( .D(n3213), .CK(n3891), .RN(n3341), .QN(n105) );
  DFFR_X1 \registers_reg[4][22]  ( .D(n3212), .CK(n3891), .RN(n3341), .QN(n106) );
  DFFR_X1 \registers_reg[4][21]  ( .D(n3211), .CK(n3891), .RN(n3341), .QN(n107) );
  DFFR_X1 \registers_reg[4][20]  ( .D(n3210), .CK(n3891), .RN(n3341), .QN(n108) );
  DFFR_X1 \registers_reg[4][19]  ( .D(n3209), .CK(n3891), .RN(n3341), .QN(n109) );
  DFFR_X1 \registers_reg[4][18]  ( .D(n3208), .CK(n3891), .RN(n3341), .QN(n110) );
  DFFR_X1 \registers_reg[4][17]  ( .D(n3207), .CK(n3891), .RN(n3341), .QN(n111) );
  DFFR_X1 \registers_reg[4][16]  ( .D(n3206), .CK(n3891), .RN(n3341), .QN(n112) );
  DFFR_X1 \registers_reg[4][15]  ( .D(n3205), .CK(n3891), .RN(n3340), .QN(n113) );
  DFFR_X1 \registers_reg[4][14]  ( .D(n3204), .CK(n3891), .RN(n3340), .QN(n114) );
  DFFR_X1 \registers_reg[4][13]  ( .D(n3203), .CK(n3891), .RN(n3340), .QN(n115) );
  DFFR_X1 \registers_reg[4][12]  ( .D(n3202), .CK(n3891), .RN(n3340), .QN(n116) );
  DFFR_X1 \registers_reg[4][11]  ( .D(n3201), .CK(n3891), .RN(n3340), .QN(n117) );
  DFFR_X1 \registers_reg[4][10]  ( .D(n3200), .CK(n3891), .RN(n3340), .QN(n118) );
  DFFR_X1 \registers_reg[4][9]  ( .D(n3199), .CK(n3891), .RN(n3340), .QN(n119)
         );
  DFFR_X1 \registers_reg[4][8]  ( .D(n3198), .CK(n3891), .RN(n3340), .QN(n120)
         );
  DFFR_X1 \registers_reg[4][7]  ( .D(n3197), .CK(n3891), .RN(n3340), .QN(n121)
         );
  DFFR_X1 \registers_reg[4][6]  ( .D(n3196), .CK(n3891), .RN(n3340), .QN(n122)
         );
  DFFR_X1 \registers_reg[4][5]  ( .D(n3195), .CK(n3891), .RN(n3340), .QN(n123)
         );
  DFFR_X1 \registers_reg[4][4]  ( .D(n3194), .CK(n3891), .RN(n3339), .QN(n124)
         );
  DFFR_X1 \registers_reg[4][3]  ( .D(n3193), .CK(n3891), .RN(n3339), .QN(n125)
         );
  DFFR_X1 \registers_reg[4][2]  ( .D(n3192), .CK(n3891), .RN(n3339), .QN(n126)
         );
  DFFR_X1 \registers_reg[4][1]  ( .D(n3191), .CK(n3891), .RN(n3339), .QN(n127)
         );
  DFFR_X1 \registers_reg[4][0]  ( .D(n3190), .CK(n3891), .RN(n3339), .QN(n128)
         );
  DFFR_X1 \registers_reg[5][31]  ( .D(n3189), .CK(n3891), .RN(n3339), .QN(n129) );
  DFFR_X1 \registers_reg[5][30]  ( .D(n3188), .CK(n3891), .RN(n3339), .QN(n130) );
  DFFR_X1 \registers_reg[5][29]  ( .D(n3187), .CK(n3891), .RN(n3339), .QN(n131) );
  DFFR_X1 \registers_reg[5][28]  ( .D(n3186), .CK(n3891), .RN(n3339), .QN(n132) );
  DFFR_X1 \registers_reg[5][27]  ( .D(n3185), .CK(n3891), .RN(n3339), .QN(n133) );
  DFFR_X1 \registers_reg[5][26]  ( .D(n3184), .CK(n3891), .RN(n3339), .QN(n134) );
  DFFR_X1 \registers_reg[5][25]  ( .D(n3183), .CK(n3891), .RN(n3338), .QN(n135) );
  DFFR_X1 \registers_reg[5][24]  ( .D(n3182), .CK(n3891), .RN(n3338), .QN(n136) );
  DFFR_X1 \registers_reg[5][23]  ( .D(n3181), .CK(n3891), .RN(n3338), .QN(n137) );
  DFFR_X1 \registers_reg[5][22]  ( .D(n3180), .CK(n3891), .RN(n3338), .QN(n138) );
  DFFR_X1 \registers_reg[5][21]  ( .D(n3179), .CK(n3891), .RN(n3338), .QN(n139) );
  DFFR_X1 \registers_reg[5][20]  ( .D(n3178), .CK(n3891), .RN(n3338), .QN(n140) );
  DFFR_X1 \registers_reg[5][19]  ( .D(n3177), .CK(n3891), .RN(n3338), .QN(n141) );
  DFFR_X1 \registers_reg[5][18]  ( .D(n3176), .CK(n3891), .RN(n3338), .QN(n142) );
  DFFR_X1 \registers_reg[5][17]  ( .D(n3175), .CK(n3891), .RN(n3338), .QN(n143) );
  DFFR_X1 \registers_reg[5][16]  ( .D(n3174), .CK(n3891), .RN(n3338), .QN(n144) );
  DFFR_X1 \registers_reg[5][15]  ( .D(n3173), .CK(n3891), .RN(n3338), .QN(n145) );
  DFFR_X1 \registers_reg[5][14]  ( .D(n3172), .CK(n3891), .RN(n3337), .QN(n146) );
  DFFR_X1 \registers_reg[5][13]  ( .D(n3171), .CK(n3891), .RN(n3337), .QN(n147) );
  DFFR_X1 \registers_reg[5][12]  ( .D(n3170), .CK(n3891), .RN(n3337), .QN(n148) );
  DFFR_X1 \registers_reg[5][11]  ( .D(n3169), .CK(n3891), .RN(n3337), .QN(n149) );
  DFFR_X1 \registers_reg[5][10]  ( .D(n3168), .CK(n3891), .RN(n3337), .QN(n150) );
  DFFR_X1 \registers_reg[5][9]  ( .D(n3167), .CK(n3891), .RN(n3337), .QN(n151)
         );
  DFFR_X1 \registers_reg[5][8]  ( .D(n3166), .CK(n3891), .RN(n3337), .QN(n152)
         );
  DFFR_X1 \registers_reg[5][7]  ( .D(n3165), .CK(n3891), .RN(n3337), .QN(n153)
         );
  DFFR_X1 \registers_reg[5][6]  ( .D(n3164), .CK(n3891), .RN(n3337), .QN(n154)
         );
  DFFR_X1 \registers_reg[5][5]  ( .D(n3163), .CK(n3891), .RN(n3337), .QN(n155)
         );
  DFFR_X1 \registers_reg[5][4]  ( .D(n3162), .CK(n3891), .RN(n3337), .QN(n156)
         );
  DFFR_X1 \registers_reg[5][3]  ( .D(n3161), .CK(n3891), .RN(n3336), .QN(n157)
         );
  DFFR_X1 \registers_reg[5][2]  ( .D(n3160), .CK(n3891), .RN(n3336), .QN(n158)
         );
  DFFR_X1 \registers_reg[5][1]  ( .D(n3159), .CK(n3891), .RN(n3336), .QN(n159)
         );
  DFFR_X1 \registers_reg[5][0]  ( .D(n3158), .CK(n3891), .RN(n3336), .QN(n160)
         );
  DFFR_X1 \registers_reg[6][31]  ( .D(n3559), .CK(n3891), .RN(n3336), .Q(
        \registers[6][31] ) );
  DFFR_X1 \registers_reg[6][30]  ( .D(n3558), .CK(n3891), .RN(n3336), .Q(
        \registers[6][30] ) );
  DFFR_X1 \registers_reg[6][29]  ( .D(n3557), .CK(n3891), .RN(n3336), .Q(
        \registers[6][29] ) );
  DFFR_X1 \registers_reg[6][28]  ( .D(n3556), .CK(n3891), .RN(n3336), .Q(
        \registers[6][28] ) );
  DFFR_X1 \registers_reg[6][27]  ( .D(n3555), .CK(n3891), .RN(n3336), .Q(
        \registers[6][27] ) );
  DFFR_X1 \registers_reg[6][26]  ( .D(n3554), .CK(n3891), .RN(n3336), .Q(
        \registers[6][26] ) );
  DFFR_X1 \registers_reg[6][25]  ( .D(n3553), .CK(n3891), .RN(n3336), .Q(
        \registers[6][25] ) );
  DFFR_X1 \registers_reg[6][24]  ( .D(n3552), .CK(n3891), .RN(n3335), .Q(
        \registers[6][24] ) );
  DFFR_X1 \registers_reg[6][23]  ( .D(n3551), .CK(n3891), .RN(n3335), .Q(
        \registers[6][23] ) );
  DFFR_X1 \registers_reg[6][22]  ( .D(n3550), .CK(n3891), .RN(n3335), .Q(
        \registers[6][22] ) );
  DFFR_X1 \registers_reg[6][21]  ( .D(n3549), .CK(n3891), .RN(n3335), .Q(
        \registers[6][21] ) );
  DFFR_X1 \registers_reg[6][20]  ( .D(n3548), .CK(n3891), .RN(n3335), .Q(
        \registers[6][20] ) );
  DFFR_X1 \registers_reg[6][19]  ( .D(n3547), .CK(n3891), .RN(n3335), .Q(
        \registers[6][19] ) );
  DFFR_X1 \registers_reg[6][18]  ( .D(n3546), .CK(n3891), .RN(n3335), .Q(
        \registers[6][18] ) );
  DFFR_X1 \registers_reg[6][17]  ( .D(n3545), .CK(n3891), .RN(n3335), .Q(
        \registers[6][17] ) );
  DFFR_X1 \registers_reg[6][16]  ( .D(n3544), .CK(n3891), .RN(n3335), .Q(
        \registers[6][16] ) );
  DFFR_X1 \registers_reg[6][15]  ( .D(n3543), .CK(n3891), .RN(n3335), .Q(
        \registers[6][15] ) );
  DFFR_X1 \registers_reg[6][14]  ( .D(n3542), .CK(n3891), .RN(n3335), .Q(
        \registers[6][14] ) );
  DFFR_X1 \registers_reg[6][13]  ( .D(n3541), .CK(n3891), .RN(n3334), .Q(
        \registers[6][13] ) );
  DFFR_X1 \registers_reg[6][12]  ( .D(n3540), .CK(n3891), .RN(n3334), .Q(
        \registers[6][12] ) );
  DFFR_X1 \registers_reg[6][11]  ( .D(n3539), .CK(n3891), .RN(n3334), .Q(
        \registers[6][11] ) );
  DFFR_X1 \registers_reg[6][10]  ( .D(n3538), .CK(n3891), .RN(n3334), .Q(
        \registers[6][10] ) );
  DFFR_X1 \registers_reg[6][9]  ( .D(n3537), .CK(n3891), .RN(n3334), .Q(
        \registers[6][9] ) );
  DFFR_X1 \registers_reg[6][8]  ( .D(n3536), .CK(n3891), .RN(n3334), .Q(
        \registers[6][8] ) );
  DFFR_X1 \registers_reg[6][7]  ( .D(n3535), .CK(n3891), .RN(n3334), .Q(
        \registers[6][7] ) );
  DFFR_X1 \registers_reg[6][6]  ( .D(n3534), .CK(n3891), .RN(n3334), .Q(
        \registers[6][6] ) );
  DFFR_X1 \registers_reg[6][5]  ( .D(n3533), .CK(n3891), .RN(n3334), .Q(
        \registers[6][5] ) );
  DFFR_X1 \registers_reg[6][4]  ( .D(n3532), .CK(n3891), .RN(n3334), .Q(
        \registers[6][4] ) );
  DFFR_X1 \registers_reg[6][3]  ( .D(n3531), .CK(n3891), .RN(n3334), .Q(
        \registers[6][3] ) );
  DFFR_X1 \registers_reg[6][2]  ( .D(n3530), .CK(n3891), .RN(n3333), .Q(
        \registers[6][2] ) );
  DFFR_X1 \registers_reg[6][1]  ( .D(n3529), .CK(n3891), .RN(n3333), .Q(
        \registers[6][1] ) );
  DFFR_X1 \registers_reg[6][0]  ( .D(n3528), .CK(n3891), .RN(n3333), .Q(
        \registers[6][0] ) );
  DFFR_X1 \registers_reg[7][31]  ( .D(n3591), .CK(n3891), .RN(n3333), .Q(
        \registers[7][31] ) );
  DFFR_X1 \registers_reg[7][30]  ( .D(n3590), .CK(n3891), .RN(n3333), .Q(
        \registers[7][30] ) );
  DFFR_X1 \registers_reg[7][29]  ( .D(n3589), .CK(n3891), .RN(n3333), .Q(
        \registers[7][29] ) );
  DFFR_X1 \registers_reg[7][28]  ( .D(n3588), .CK(n3891), .RN(n3333), .Q(
        \registers[7][28] ) );
  DFFR_X1 \registers_reg[7][27]  ( .D(n3587), .CK(n3891), .RN(n3333), .Q(
        \registers[7][27] ) );
  DFFR_X1 \registers_reg[7][26]  ( .D(n3586), .CK(n3891), .RN(n3333), .Q(
        \registers[7][26] ) );
  DFFR_X1 \registers_reg[7][25]  ( .D(n3585), .CK(n3891), .RN(n3333), .Q(
        \registers[7][25] ) );
  DFFR_X1 \registers_reg[7][24]  ( .D(n3584), .CK(n3891), .RN(n3333), .Q(
        \registers[7][24] ) );
  DFFR_X1 \registers_reg[7][23]  ( .D(n3583), .CK(n3891), .RN(n3332), .Q(
        \registers[7][23] ) );
  DFFR_X1 \registers_reg[7][22]  ( .D(n3582), .CK(n3891), .RN(n3332), .Q(
        \registers[7][22] ) );
  DFFR_X1 \registers_reg[7][21]  ( .D(n3581), .CK(n3891), .RN(n3332), .Q(
        \registers[7][21] ) );
  DFFR_X1 \registers_reg[7][20]  ( .D(n3580), .CK(n3891), .RN(n3332), .Q(
        \registers[7][20] ) );
  DFFR_X1 \registers_reg[7][19]  ( .D(n3579), .CK(n3891), .RN(n3332), .Q(
        \registers[7][19] ) );
  DFFR_X1 \registers_reg[7][18]  ( .D(n3578), .CK(n3891), .RN(n3332), .Q(
        \registers[7][18] ) );
  DFFR_X1 \registers_reg[7][17]  ( .D(n3577), .CK(n3891), .RN(n3332), .Q(
        \registers[7][17] ) );
  DFFR_X1 \registers_reg[7][16]  ( .D(n3576), .CK(n3891), .RN(n3332), .Q(
        \registers[7][16] ) );
  DFFR_X1 \registers_reg[7][15]  ( .D(n3575), .CK(n3891), .RN(n3332), .Q(
        \registers[7][15] ) );
  DFFR_X1 \registers_reg[7][14]  ( .D(n3574), .CK(n3891), .RN(n3332), .Q(
        \registers[7][14] ) );
  DFFR_X1 \registers_reg[7][13]  ( .D(n3573), .CK(n3891), .RN(n3332), .Q(
        \registers[7][13] ) );
  DFFR_X1 \registers_reg[7][12]  ( .D(n3572), .CK(n3891), .RN(n3331), .Q(
        \registers[7][12] ) );
  DFFR_X1 \registers_reg[7][11]  ( .D(n3571), .CK(n3891), .RN(n3331), .Q(
        \registers[7][11] ) );
  DFFR_X1 \registers_reg[7][10]  ( .D(n3570), .CK(n3891), .RN(n3331), .Q(
        \registers[7][10] ) );
  DFFR_X1 \registers_reg[7][9]  ( .D(n3569), .CK(n3891), .RN(n3331), .Q(
        \registers[7][9] ) );
  DFFR_X1 \registers_reg[7][8]  ( .D(n3568), .CK(n3891), .RN(n3331), .Q(
        \registers[7][8] ) );
  DFFR_X1 \registers_reg[7][7]  ( .D(n3567), .CK(n3891), .RN(n3331), .Q(
        \registers[7][7] ) );
  DFFR_X1 \registers_reg[7][6]  ( .D(n3566), .CK(n3891), .RN(n3331), .Q(
        \registers[7][6] ) );
  DFFR_X1 \registers_reg[7][5]  ( .D(n3565), .CK(n3891), .RN(n3331), .Q(
        \registers[7][5] ) );
  DFFR_X1 \registers_reg[7][4]  ( .D(n3564), .CK(n3891), .RN(n3331), .Q(
        \registers[7][4] ) );
  DFFR_X1 \registers_reg[7][3]  ( .D(n3563), .CK(n3891), .RN(n3331), .Q(
        \registers[7][3] ) );
  DFFR_X1 \registers_reg[7][2]  ( .D(n3562), .CK(n3891), .RN(n3331), .Q(
        \registers[7][2] ) );
  DFFR_X1 \registers_reg[7][1]  ( .D(n3561), .CK(n3891), .RN(n3330), .Q(
        \registers[7][1] ) );
  DFFR_X1 \registers_reg[7][0]  ( .D(n3560), .CK(n3891), .RN(n3330), .Q(
        \registers[7][0] ) );
  DFFR_X1 \registers_reg[8][31]  ( .D(n3399), .CK(n3891), .RN(n3330), .Q(
        \registers[8][31] ) );
  DFFR_X1 \registers_reg[8][30]  ( .D(n3398), .CK(n3891), .RN(n3330), .Q(
        \registers[8][30] ) );
  DFFR_X1 \registers_reg[8][29]  ( .D(n3397), .CK(n3891), .RN(n3330), .Q(
        \registers[8][29] ) );
  DFFR_X1 \registers_reg[8][28]  ( .D(n3396), .CK(n3891), .RN(n3330), .Q(
        \registers[8][28] ) );
  DFFR_X1 \registers_reg[8][27]  ( .D(n3395), .CK(n3891), .RN(n3330), .Q(
        \registers[8][27] ) );
  DFFR_X1 \registers_reg[8][26]  ( .D(n3394), .CK(n3891), .RN(n3330), .Q(
        \registers[8][26] ) );
  DFFR_X1 \registers_reg[8][25]  ( .D(n3393), .CK(n3891), .RN(n3330), .Q(
        \registers[8][25] ) );
  DFFR_X1 \registers_reg[8][24]  ( .D(n3392), .CK(n3891), .RN(n3330), .Q(
        \registers[8][24] ) );
  DFFR_X1 \registers_reg[8][23]  ( .D(n3391), .CK(n3891), .RN(n3330), .Q(
        \registers[8][23] ) );
  DFFR_X1 \registers_reg[8][22]  ( .D(n3390), .CK(n3891), .RN(n3329), .Q(
        \registers[8][22] ) );
  DFFR_X1 \registers_reg[8][21]  ( .D(n3389), .CK(n3891), .RN(n3329), .Q(
        \registers[8][21] ) );
  DFFR_X1 \registers_reg[8][20]  ( .D(n3388), .CK(n3891), .RN(n3329), .Q(
        \registers[8][20] ) );
  DFFR_X1 \registers_reg[8][19]  ( .D(n3387), .CK(n3891), .RN(n3329), .Q(
        \registers[8][19] ) );
  DFFR_X1 \registers_reg[8][18]  ( .D(n3386), .CK(n3891), .RN(n3329), .Q(
        \registers[8][18] ) );
  DFFR_X1 \registers_reg[8][17]  ( .D(n3385), .CK(n3891), .RN(n3329), .Q(
        \registers[8][17] ) );
  DFFR_X1 \registers_reg[8][16]  ( .D(n3384), .CK(n3891), .RN(n3329), .Q(
        \registers[8][16] ) );
  DFFR_X1 \registers_reg[8][15]  ( .D(n3383), .CK(n3891), .RN(n3329), .Q(
        \registers[8][15] ) );
  DFFR_X1 \registers_reg[8][14]  ( .D(n3382), .CK(n3891), .RN(n3329), .Q(
        \registers[8][14] ) );
  DFFR_X1 \registers_reg[8][13]  ( .D(n3381), .CK(n3891), .RN(n3329), .Q(
        \registers[8][13] ) );
  DFFR_X1 \registers_reg[8][12]  ( .D(n3380), .CK(n3891), .RN(n3329), .Q(
        \registers[8][12] ) );
  DFFR_X1 \registers_reg[8][11]  ( .D(n3379), .CK(n3891), .RN(n3328), .Q(
        \registers[8][11] ) );
  DFFR_X1 \registers_reg[8][10]  ( .D(n3378), .CK(n3891), .RN(n3328), .Q(
        \registers[8][10] ) );
  DFFR_X1 \registers_reg[8][9]  ( .D(n3377), .CK(n3891), .RN(n3328), .Q(
        \registers[8][9] ) );
  DFFR_X1 \registers_reg[8][8]  ( .D(n3376), .CK(n3891), .RN(n3328), .Q(
        \registers[8][8] ) );
  DFFR_X1 \registers_reg[8][7]  ( .D(n3375), .CK(n3891), .RN(n3328), .Q(
        \registers[8][7] ) );
  DFFR_X1 \registers_reg[8][6]  ( .D(n3374), .CK(n3891), .RN(n3328), .Q(
        \registers[8][6] ) );
  DFFR_X1 \registers_reg[8][5]  ( .D(n3373), .CK(n3891), .RN(n3328), .Q(
        \registers[8][5] ) );
  DFFR_X1 \registers_reg[8][4]  ( .D(n3372), .CK(n3891), .RN(n3328), .Q(
        \registers[8][4] ) );
  DFFR_X1 \registers_reg[8][3]  ( .D(n3371), .CK(n3891), .RN(n3328), .Q(
        \registers[8][3] ) );
  DFFR_X1 \registers_reg[8][2]  ( .D(n3370), .CK(n3891), .RN(n3328), .Q(
        \registers[8][2] ) );
  DFFR_X1 \registers_reg[8][1]  ( .D(n3369), .CK(n3891), .RN(n3328), .Q(
        \registers[8][1] ) );
  DFFR_X1 \registers_reg[8][0]  ( .D(n3368), .CK(n3891), .RN(n3327), .Q(
        \registers[8][0] ) );
  DFFR_X1 \registers_reg[9][31]  ( .D(n3431), .CK(n3891), .RN(n3327), .Q(
        \registers[9][31] ) );
  DFFR_X1 \registers_reg[9][30]  ( .D(n3430), .CK(n3891), .RN(n3327), .Q(
        \registers[9][30] ) );
  DFFR_X1 \registers_reg[9][29]  ( .D(n3429), .CK(n3891), .RN(n3327), .Q(
        \registers[9][29] ) );
  DFFR_X1 \registers_reg[9][28]  ( .D(n3428), .CK(n3891), .RN(n3327), .Q(
        \registers[9][28] ) );
  DFFR_X1 \registers_reg[9][27]  ( .D(n3427), .CK(n3891), .RN(n3327), .Q(
        \registers[9][27] ) );
  DFFR_X1 \registers_reg[9][26]  ( .D(n3426), .CK(n3891), .RN(n3327), .Q(
        \registers[9][26] ) );
  DFFR_X1 \registers_reg[9][25]  ( .D(n3425), .CK(n3891), .RN(n3327), .Q(
        \registers[9][25] ) );
  DFFR_X1 \registers_reg[9][24]  ( .D(n3424), .CK(n3891), .RN(n3327), .Q(
        \registers[9][24] ) );
  DFFR_X1 \registers_reg[9][23]  ( .D(n3423), .CK(n3891), .RN(n3327), .Q(
        \registers[9][23] ) );
  DFFR_X1 \registers_reg[9][22]  ( .D(n3422), .CK(n3891), .RN(n3327), .Q(
        \registers[9][22] ) );
  DFFR_X1 \registers_reg[9][21]  ( .D(n3421), .CK(n3891), .RN(n3326), .Q(
        \registers[9][21] ) );
  DFFR_X1 \registers_reg[9][20]  ( .D(n3420), .CK(n3891), .RN(n3326), .Q(
        \registers[9][20] ) );
  DFFR_X1 \registers_reg[9][19]  ( .D(n3419), .CK(n3891), .RN(n3326), .Q(
        \registers[9][19] ) );
  DFFR_X1 \registers_reg[9][18]  ( .D(n3418), .CK(n3891), .RN(n3326), .Q(
        \registers[9][18] ) );
  DFFR_X1 \registers_reg[9][17]  ( .D(n3417), .CK(n3891), .RN(n3326), .Q(
        \registers[9][17] ) );
  DFFR_X1 \registers_reg[9][16]  ( .D(n3416), .CK(n3891), .RN(n3326), .Q(
        \registers[9][16] ) );
  DFFR_X1 \registers_reg[9][15]  ( .D(n3415), .CK(n3891), .RN(n3326), .Q(
        \registers[9][15] ) );
  DFFR_X1 \registers_reg[9][14]  ( .D(n3414), .CK(n3891), .RN(n3326), .Q(
        \registers[9][14] ) );
  DFFR_X1 \registers_reg[9][13]  ( .D(n3413), .CK(n3891), .RN(n3326), .Q(
        \registers[9][13] ) );
  DFFR_X1 \registers_reg[9][12]  ( .D(n3412), .CK(n3891), .RN(n3326), .Q(
        \registers[9][12] ) );
  DFFR_X1 \registers_reg[9][11]  ( .D(n3411), .CK(n3891), .RN(n3326), .Q(
        \registers[9][11] ) );
  DFFR_X1 \registers_reg[9][10]  ( .D(n3410), .CK(n3891), .RN(n3325), .Q(
        \registers[9][10] ) );
  DFFR_X1 \registers_reg[9][9]  ( .D(n3409), .CK(n3891), .RN(n3325), .Q(
        \registers[9][9] ) );
  DFFR_X1 \registers_reg[9][8]  ( .D(n3408), .CK(n3891), .RN(n3325), .Q(
        \registers[9][8] ) );
  DFFR_X1 \registers_reg[9][7]  ( .D(n3407), .CK(n3891), .RN(n3325), .Q(
        \registers[9][7] ) );
  DFFR_X1 \registers_reg[9][6]  ( .D(n3406), .CK(n3891), .RN(n3325), .Q(
        \registers[9][6] ) );
  DFFR_X1 \registers_reg[9][5]  ( .D(n3405), .CK(n3891), .RN(n3325), .Q(
        \registers[9][5] ) );
  DFFR_X1 \registers_reg[9][4]  ( .D(n3404), .CK(n3891), .RN(n3325), .Q(
        \registers[9][4] ) );
  DFFR_X1 \registers_reg[9][3]  ( .D(n3403), .CK(n3891), .RN(n3325), .Q(
        \registers[9][3] ) );
  DFFR_X1 \registers_reg[9][2]  ( .D(n3402), .CK(n3891), .RN(n3325), .Q(
        \registers[9][2] ) );
  DFFR_X1 \registers_reg[9][1]  ( .D(n3401), .CK(n3891), .RN(n3325), .Q(
        \registers[9][1] ) );
  DFFR_X1 \registers_reg[9][0]  ( .D(n3400), .CK(n3891), .RN(n3325), .Q(
        \registers[9][0] ) );
  DFFR_X1 \registers_reg[10][31]  ( .D(n3157), .CK(n3891), .RN(n3324), .QN(
        n289) );
  DFFR_X1 \registers_reg[10][30]  ( .D(n3156), .CK(n3891), .RN(n3324), .QN(
        n290) );
  DFFR_X1 \registers_reg[10][29]  ( .D(n3155), .CK(n3891), .RN(n3324), .QN(
        n291) );
  DFFR_X1 \registers_reg[10][28]  ( .D(n3154), .CK(n3891), .RN(n3324), .QN(
        n292) );
  DFFR_X1 \registers_reg[10][27]  ( .D(n3153), .CK(n3891), .RN(n3324), .QN(
        n293) );
  DFFR_X1 \registers_reg[10][26]  ( .D(n3152), .CK(n3891), .RN(n3324), .QN(
        n294) );
  DFFR_X1 \registers_reg[10][25]  ( .D(n3151), .CK(n3891), .RN(n3324), .QN(
        n295) );
  DFFR_X1 \registers_reg[10][24]  ( .D(n3150), .CK(n3891), .RN(n3324), .QN(
        n296) );
  DFFR_X1 \registers_reg[10][23]  ( .D(n3149), .CK(n3891), .RN(n3324), .QN(
        n297) );
  DFFR_X1 \registers_reg[10][22]  ( .D(n3148), .CK(n3891), .RN(n3324), .QN(
        n298) );
  DFFR_X1 \registers_reg[10][21]  ( .D(n3147), .CK(n3891), .RN(n3324), .QN(
        n299) );
  DFFR_X1 \registers_reg[10][20]  ( .D(n3146), .CK(n3891), .RN(n3323), .QN(
        n300) );
  DFFR_X1 \registers_reg[10][19]  ( .D(n3145), .CK(n3891), .RN(n3323), .QN(
        n301) );
  DFFR_X1 \registers_reg[10][18]  ( .D(n3144), .CK(n3891), .RN(n3323), .QN(
        n302) );
  DFFR_X1 \registers_reg[10][17]  ( .D(n3143), .CK(n3891), .RN(n3323), .QN(
        n303) );
  DFFR_X1 \registers_reg[10][16]  ( .D(n3142), .CK(n3891), .RN(n3323), .QN(
        n304) );
  DFFR_X1 \registers_reg[10][15]  ( .D(n3141), .CK(n3891), .RN(n3323), .QN(
        n305) );
  DFFR_X1 \registers_reg[10][14]  ( .D(n3140), .CK(n3891), .RN(n3323), .QN(
        n306) );
  DFFR_X1 \registers_reg[10][13]  ( .D(n3139), .CK(n3891), .RN(n3323), .QN(
        n307) );
  DFFR_X1 \registers_reg[10][12]  ( .D(n3138), .CK(n3891), .RN(n3323), .QN(
        n308) );
  DFFR_X1 \registers_reg[10][11]  ( .D(n3137), .CK(n3891), .RN(n3323), .QN(
        n309) );
  DFFR_X1 \registers_reg[10][10]  ( .D(n3136), .CK(n3891), .RN(n3323), .QN(
        n310) );
  DFFR_X1 \registers_reg[10][9]  ( .D(n3135), .CK(n3891), .RN(n3322), .QN(n311) );
  DFFR_X1 \registers_reg[10][8]  ( .D(n3134), .CK(n3891), .RN(n3322), .QN(n312) );
  DFFR_X1 \registers_reg[10][7]  ( .D(n3133), .CK(n3891), .RN(n3322), .QN(n313) );
  DFFR_X1 \registers_reg[10][6]  ( .D(n3132), .CK(n3891), .RN(n3322), .QN(n314) );
  DFFR_X1 \registers_reg[10][5]  ( .D(n3131), .CK(n3891), .RN(n3322), .QN(n315) );
  DFFR_X1 \registers_reg[10][4]  ( .D(n3130), .CK(n3891), .RN(n3322), .QN(n316) );
  DFFR_X1 \registers_reg[10][3]  ( .D(n3129), .CK(n3891), .RN(n3322), .QN(n317) );
  DFFR_X1 \registers_reg[10][2]  ( .D(n3128), .CK(n3891), .RN(n3322), .QN(n318) );
  DFFR_X1 \registers_reg[10][1]  ( .D(n3127), .CK(n3891), .RN(n3322), .QN(n319) );
  DFFR_X1 \registers_reg[10][0]  ( .D(n3126), .CK(n3891), .RN(n3322), .QN(n320) );
  DFFR_X1 \registers_reg[11][31]  ( .D(n3125), .CK(n3891), .RN(n3322), .QN(
        n321) );
  DFFR_X1 \registers_reg[11][30]  ( .D(n3124), .CK(n3891), .RN(n3321), .QN(
        n322) );
  DFFR_X1 \registers_reg[11][29]  ( .D(n3123), .CK(n3891), .RN(n3321), .QN(
        n323) );
  DFFR_X1 \registers_reg[11][28]  ( .D(n3122), .CK(n3891), .RN(n3321), .QN(
        n324) );
  DFFR_X1 \registers_reg[11][27]  ( .D(n3121), .CK(n3891), .RN(n3321), .QN(
        n325) );
  DFFR_X1 \registers_reg[11][26]  ( .D(n3120), .CK(n3891), .RN(n3321), .QN(
        n326) );
  DFFR_X1 \registers_reg[11][25]  ( .D(n3119), .CK(n3891), .RN(n3321), .QN(
        n327) );
  DFFR_X1 \registers_reg[11][24]  ( .D(n3118), .CK(n3891), .RN(n3321), .QN(
        n328) );
  DFFR_X1 \registers_reg[11][23]  ( .D(n3117), .CK(n3891), .RN(n3321), .QN(
        n329) );
  DFFR_X1 \registers_reg[11][22]  ( .D(n3116), .CK(n3891), .RN(n3321), .QN(
        n330) );
  DFFR_X1 \registers_reg[11][21]  ( .D(n3115), .CK(n3891), .RN(n3321), .QN(
        n331) );
  DFFR_X1 \registers_reg[11][20]  ( .D(n3114), .CK(n3891), .RN(n3321), .QN(
        n332) );
  DFFR_X1 \registers_reg[11][19]  ( .D(n3113), .CK(n3891), .RN(n3320), .QN(
        n333) );
  DFFR_X1 \registers_reg[11][18]  ( .D(n3112), .CK(n3891), .RN(n3320), .QN(
        n334) );
  DFFR_X1 \registers_reg[11][17]  ( .D(n3111), .CK(n3891), .RN(n3320), .QN(
        n335) );
  DFFR_X1 \registers_reg[11][16]  ( .D(n3110), .CK(n3891), .RN(n3320), .QN(
        n336) );
  DFFR_X1 \registers_reg[11][15]  ( .D(n3109), .CK(n3891), .RN(n3320), .QN(
        n337) );
  DFFR_X1 \registers_reg[11][14]  ( .D(n3108), .CK(n3891), .RN(n3320), .QN(
        n338) );
  DFFR_X1 \registers_reg[11][13]  ( .D(n3107), .CK(n3891), .RN(n3320), .QN(
        n339) );
  DFFR_X1 \registers_reg[11][12]  ( .D(n3106), .CK(n3891), .RN(n3320), .QN(
        n340) );
  DFFR_X1 \registers_reg[11][11]  ( .D(n3105), .CK(n3891), .RN(n3320), .QN(
        n341) );
  DFFR_X1 \registers_reg[11][10]  ( .D(n3104), .CK(n3891), .RN(n3320), .QN(
        n342) );
  DFFR_X1 \registers_reg[11][9]  ( .D(n3103), .CK(n3891), .RN(n3320), .QN(n343) );
  DFFR_X1 \registers_reg[11][8]  ( .D(n3102), .CK(n3891), .RN(n3319), .QN(n344) );
  DFFR_X1 \registers_reg[11][7]  ( .D(n3101), .CK(n3891), .RN(n3319), .QN(n345) );
  DFFR_X1 \registers_reg[11][6]  ( .D(n3100), .CK(n3891), .RN(n3319), .QN(n346) );
  DFFR_X1 \registers_reg[11][5]  ( .D(n3099), .CK(n3891), .RN(n3319), .QN(n347) );
  DFFR_X1 \registers_reg[11][4]  ( .D(n3098), .CK(n3891), .RN(n3319), .QN(n348) );
  DFFR_X1 \registers_reg[11][3]  ( .D(n3097), .CK(n3891), .RN(n3319), .QN(n349) );
  DFFR_X1 \registers_reg[11][2]  ( .D(n3096), .CK(n3891), .RN(n3319), .QN(n350) );
  DFFR_X1 \registers_reg[11][1]  ( .D(n3095), .CK(n3891), .RN(n3319), .QN(n351) );
  DFFR_X1 \registers_reg[11][0]  ( .D(n3094), .CK(n3891), .RN(n3319), .QN(n352) );
  DFFR_X1 \registers_reg[12][31]  ( .D(n3463), .CK(n3891), .RN(n3319), .Q(
        \registers[12][31] ) );
  DFFR_X1 \registers_reg[12][30]  ( .D(n3462), .CK(n3891), .RN(n3319), .Q(
        \registers[12][30] ) );
  DFFR_X1 \registers_reg[12][29]  ( .D(n3461), .CK(n3891), .RN(n3318), .Q(
        \registers[12][29] ) );
  DFFR_X1 \registers_reg[12][28]  ( .D(n3460), .CK(n3891), .RN(n3318), .Q(
        \registers[12][28] ) );
  DFFR_X1 \registers_reg[12][27]  ( .D(n3459), .CK(n3891), .RN(n3318), .Q(
        \registers[12][27] ) );
  DFFR_X1 \registers_reg[12][26]  ( .D(n3458), .CK(n3891), .RN(n3318), .Q(
        \registers[12][26] ) );
  DFFR_X1 \registers_reg[12][25]  ( .D(n3457), .CK(n3891), .RN(n3318), .Q(
        \registers[12][25] ) );
  DFFR_X1 \registers_reg[12][24]  ( .D(n3456), .CK(n3891), .RN(n3318), .Q(
        \registers[12][24] ) );
  DFFR_X1 \registers_reg[12][23]  ( .D(n3455), .CK(n3891), .RN(n3318), .Q(
        \registers[12][23] ) );
  DFFR_X1 \registers_reg[12][22]  ( .D(n3454), .CK(n3891), .RN(n3318), .Q(
        \registers[12][22] ) );
  DFFR_X1 \registers_reg[12][21]  ( .D(n3453), .CK(n3891), .RN(n3318), .Q(
        \registers[12][21] ) );
  DFFR_X1 \registers_reg[12][20]  ( .D(n3452), .CK(n3891), .RN(n3318), .Q(
        \registers[12][20] ) );
  DFFR_X1 \registers_reg[12][19]  ( .D(n3451), .CK(n3891), .RN(n3318), .Q(
        \registers[12][19] ) );
  DFFR_X1 \registers_reg[12][18]  ( .D(n3450), .CK(n3891), .RN(n3317), .Q(
        \registers[12][18] ) );
  DFFR_X1 \registers_reg[12][17]  ( .D(n3449), .CK(n3891), .RN(n3317), .Q(
        \registers[12][17] ) );
  DFFR_X1 \registers_reg[12][16]  ( .D(n3448), .CK(n3891), .RN(n3317), .Q(
        \registers[12][16] ) );
  DFFR_X1 \registers_reg[12][15]  ( .D(n3447), .CK(n3891), .RN(n3317), .Q(
        \registers[12][15] ) );
  DFFR_X1 \registers_reg[12][14]  ( .D(n3446), .CK(n3891), .RN(n3317), .Q(
        \registers[12][14] ) );
  DFFR_X1 \registers_reg[12][13]  ( .D(n3445), .CK(n3891), .RN(n3317), .Q(
        \registers[12][13] ) );
  DFFR_X1 \registers_reg[12][12]  ( .D(n3444), .CK(n3891), .RN(n3317), .Q(
        \registers[12][12] ) );
  DFFR_X1 \registers_reg[12][11]  ( .D(n3443), .CK(n3891), .RN(n3317), .Q(
        \registers[12][11] ) );
  DFFR_X1 \registers_reg[12][10]  ( .D(n3442), .CK(n3891), .RN(n3317), .Q(
        \registers[12][10] ) );
  DFFR_X1 \registers_reg[12][9]  ( .D(n3441), .CK(n3891), .RN(n3317), .Q(
        \registers[12][9] ) );
  DFFR_X1 \registers_reg[12][8]  ( .D(n3440), .CK(n3891), .RN(n3317), .Q(
        \registers[12][8] ) );
  DFFR_X1 \registers_reg[12][7]  ( .D(n3439), .CK(n3891), .RN(n3316), .Q(
        \registers[12][7] ) );
  DFFR_X1 \registers_reg[12][6]  ( .D(n3438), .CK(n3891), .RN(n3316), .Q(
        \registers[12][6] ) );
  DFFR_X1 \registers_reg[12][5]  ( .D(n3437), .CK(n3891), .RN(n3316), .Q(
        \registers[12][5] ) );
  DFFR_X1 \registers_reg[12][4]  ( .D(n3436), .CK(n3891), .RN(n3316), .Q(
        \registers[12][4] ) );
  DFFR_X1 \registers_reg[12][3]  ( .D(n3435), .CK(n3891), .RN(n3316), .Q(
        \registers[12][3] ) );
  DFFR_X1 \registers_reg[12][2]  ( .D(n3434), .CK(n3891), .RN(n3316), .Q(
        \registers[12][2] ) );
  DFFR_X1 \registers_reg[12][1]  ( .D(n3433), .CK(n3891), .RN(n3316), .Q(
        \registers[12][1] ) );
  DFFR_X1 \registers_reg[12][0]  ( .D(n3432), .CK(n3891), .RN(n3316), .Q(
        \registers[12][0] ) );
  DFFR_X1 \registers_reg[13][31]  ( .D(n3495), .CK(n3891), .RN(n3316), .Q(
        \registers[13][31] ) );
  DFFR_X1 \registers_reg[13][30]  ( .D(n3494), .CK(n3891), .RN(n3316), .Q(
        \registers[13][30] ) );
  DFFR_X1 \registers_reg[13][29]  ( .D(n3493), .CK(n3891), .RN(n3316), .Q(
        \registers[13][29] ) );
  DFFR_X1 \registers_reg[13][28]  ( .D(n3492), .CK(n3891), .RN(n3315), .Q(
        \registers[13][28] ) );
  DFFR_X1 \registers_reg[13][27]  ( .D(n3491), .CK(n3891), .RN(n3315), .Q(
        \registers[13][27] ) );
  DFFR_X1 \registers_reg[13][26]  ( .D(n3490), .CK(n3891), .RN(n3315), .Q(
        \registers[13][26] ) );
  DFFR_X1 \registers_reg[13][25]  ( .D(n3489), .CK(n3891), .RN(n3315), .Q(
        \registers[13][25] ) );
  DFFR_X1 \registers_reg[13][24]  ( .D(n3488), .CK(n3891), .RN(n3315), .Q(
        \registers[13][24] ) );
  DFFR_X1 \registers_reg[13][23]  ( .D(n3487), .CK(n3891), .RN(n3315), .Q(
        \registers[13][23] ) );
  DFFR_X1 \registers_reg[13][22]  ( .D(n3486), .CK(n3891), .RN(n3315), .Q(
        \registers[13][22] ) );
  DFFR_X1 \registers_reg[13][21]  ( .D(n3485), .CK(n3891), .RN(n3315), .Q(
        \registers[13][21] ) );
  DFFR_X1 \registers_reg[13][20]  ( .D(n3484), .CK(n3891), .RN(n3315), .Q(
        \registers[13][20] ) );
  DFFR_X1 \registers_reg[13][19]  ( .D(n3483), .CK(n3891), .RN(n3315), .Q(
        \registers[13][19] ) );
  DFFR_X1 \registers_reg[13][18]  ( .D(n3482), .CK(n3891), .RN(n3315), .Q(
        \registers[13][18] ) );
  DFFR_X1 \registers_reg[13][17]  ( .D(n3481), .CK(n3891), .RN(n3314), .Q(
        \registers[13][17] ) );
  DFFR_X1 \registers_reg[13][16]  ( .D(n3480), .CK(n3891), .RN(n3314), .Q(
        \registers[13][16] ) );
  DFFR_X1 \registers_reg[13][15]  ( .D(n3479), .CK(n3891), .RN(n3314), .Q(
        \registers[13][15] ) );
  DFFR_X1 \registers_reg[13][14]  ( .D(n3478), .CK(n3891), .RN(n3314), .Q(
        \registers[13][14] ) );
  DFFR_X1 \registers_reg[13][13]  ( .D(n3477), .CK(n3891), .RN(n3314), .Q(
        \registers[13][13] ) );
  DFFR_X1 \registers_reg[13][12]  ( .D(n3476), .CK(n3891), .RN(n3314), .Q(
        \registers[13][12] ) );
  DFFR_X1 \registers_reg[13][11]  ( .D(n3475), .CK(n3891), .RN(n3314), .Q(
        \registers[13][11] ) );
  DFFR_X1 \registers_reg[13][10]  ( .D(n3474), .CK(n3891), .RN(n3314), .Q(
        \registers[13][10] ) );
  DFFR_X1 \registers_reg[13][9]  ( .D(n3473), .CK(n3891), .RN(n3314), .Q(
        \registers[13][9] ) );
  DFFR_X1 \registers_reg[13][8]  ( .D(n3472), .CK(n3891), .RN(n3314), .Q(
        \registers[13][8] ) );
  DFFR_X1 \registers_reg[13][7]  ( .D(n3471), .CK(n3891), .RN(n3314), .Q(
        \registers[13][7] ) );
  DFFR_X1 \registers_reg[13][6]  ( .D(n3470), .CK(n3891), .RN(n3313), .Q(
        \registers[13][6] ) );
  DFFR_X1 \registers_reg[13][5]  ( .D(n3469), .CK(n3891), .RN(n3313), .Q(
        \registers[13][5] ) );
  DFFR_X1 \registers_reg[13][4]  ( .D(n3468), .CK(n3891), .RN(n3313), .Q(
        \registers[13][4] ) );
  DFFR_X1 \registers_reg[13][3]  ( .D(n3467), .CK(n3891), .RN(n3313), .Q(
        \registers[13][3] ) );
  DFFR_X1 \registers_reg[13][2]  ( .D(n3466), .CK(n3891), .RN(n3313), .Q(
        \registers[13][2] ) );
  DFFR_X1 \registers_reg[13][1]  ( .D(n3465), .CK(n3891), .RN(n3313), .Q(
        \registers[13][1] ) );
  DFFR_X1 \registers_reg[13][0]  ( .D(n3464), .CK(n3891), .RN(n3313), .Q(
        \registers[13][0] ) );
  DFFR_X1 \registers_reg[14][31]  ( .D(n3093), .CK(n3891), .RN(n3313), .QN(
        n417) );
  DFFR_X1 \registers_reg[14][30]  ( .D(n3092), .CK(n3891), .RN(n3313), .QN(
        n418) );
  DFFR_X1 \registers_reg[14][29]  ( .D(n3091), .CK(n3891), .RN(n3313), .QN(
        n419) );
  DFFR_X1 \registers_reg[14][28]  ( .D(n3090), .CK(n3891), .RN(n3313), .QN(
        n420) );
  DFFR_X1 \registers_reg[14][27]  ( .D(n3089), .CK(n3891), .RN(n3312), .QN(
        n421) );
  DFFR_X1 \registers_reg[14][26]  ( .D(n3088), .CK(n3891), .RN(n3312), .QN(
        n422) );
  DFFR_X1 \registers_reg[14][25]  ( .D(n3087), .CK(n3891), .RN(n3312), .QN(
        n423) );
  DFFR_X1 \registers_reg[14][24]  ( .D(n3086), .CK(n3891), .RN(n3312), .QN(
        n424) );
  DFFR_X1 \registers_reg[14][23]  ( .D(n3085), .CK(n3891), .RN(n3312), .QN(
        n425) );
  DFFR_X1 \registers_reg[14][22]  ( .D(n3084), .CK(n3891), .RN(n3312), .QN(
        n426) );
  DFFR_X1 \registers_reg[14][21]  ( .D(n3083), .CK(n3891), .RN(n3312), .QN(
        n427) );
  DFFR_X1 \registers_reg[14][20]  ( .D(n3082), .CK(n3891), .RN(n3312), .QN(
        n428) );
  DFFR_X1 \registers_reg[14][19]  ( .D(n3081), .CK(n3891), .RN(n3312), .QN(
        n429) );
  DFFR_X1 \registers_reg[14][18]  ( .D(n3080), .CK(n3891), .RN(n3312), .QN(
        n430) );
  DFFR_X1 \registers_reg[14][17]  ( .D(n3079), .CK(n3891), .RN(n3312), .QN(
        n431) );
  DFFR_X1 \registers_reg[14][16]  ( .D(n3078), .CK(n3891), .RN(n3311), .QN(
        n432) );
  DFFR_X1 \registers_reg[14][15]  ( .D(n3077), .CK(n3891), .RN(n3311), .QN(
        n433) );
  DFFR_X1 \registers_reg[14][14]  ( .D(n3076), .CK(n3891), .RN(n3311), .QN(
        n434) );
  DFFR_X1 \registers_reg[14][13]  ( .D(n3075), .CK(n3891), .RN(n3311), .QN(
        n435) );
  DFFR_X1 \registers_reg[14][12]  ( .D(n3074), .CK(n3891), .RN(n3311), .QN(
        n436) );
  DFFR_X1 \registers_reg[14][11]  ( .D(n3073), .CK(n3891), .RN(n3311), .QN(
        n437) );
  DFFR_X1 \registers_reg[14][10]  ( .D(n3072), .CK(n3891), .RN(n3311), .QN(
        n438) );
  DFFR_X1 \registers_reg[14][9]  ( .D(n3071), .CK(n3891), .RN(n3311), .QN(n439) );
  DFFR_X1 \registers_reg[14][8]  ( .D(n3070), .CK(n3891), .RN(n3311), .QN(n440) );
  DFFR_X1 \registers_reg[14][7]  ( .D(n3069), .CK(n3891), .RN(n3311), .QN(n441) );
  DFFR_X1 \registers_reg[14][6]  ( .D(n3068), .CK(n3891), .RN(n3311), .QN(n442) );
  DFFR_X1 \registers_reg[14][5]  ( .D(n3067), .CK(n3891), .RN(n3310), .QN(n443) );
  DFFR_X1 \registers_reg[14][4]  ( .D(n3066), .CK(n3891), .RN(n3310), .QN(n444) );
  DFFR_X1 \registers_reg[14][3]  ( .D(n3065), .CK(n3891), .RN(n3310), .QN(n445) );
  DFFR_X1 \registers_reg[14][2]  ( .D(n3064), .CK(n3891), .RN(n3310), .QN(n446) );
  DFFR_X1 \registers_reg[14][1]  ( .D(n3063), .CK(n3891), .RN(n3310), .QN(n447) );
  DFFR_X1 \registers_reg[14][0]  ( .D(n3062), .CK(n3891), .RN(n3310), .QN(n448) );
  DFFR_X1 \registers_reg[15][31]  ( .D(n3061), .CK(n3891), .RN(n3310), .QN(
        n449) );
  DFFR_X1 \registers_reg[15][30]  ( .D(n3060), .CK(n3891), .RN(n3310), .QN(
        n450) );
  DFFR_X1 \registers_reg[15][29]  ( .D(n3059), .CK(n3891), .RN(n3310), .QN(
        n451) );
  DFFR_X1 \registers_reg[15][28]  ( .D(n3058), .CK(n3891), .RN(n3310), .QN(
        n452) );
  DFFR_X1 \registers_reg[15][27]  ( .D(n3057), .CK(n3891), .RN(n3310), .QN(
        n453) );
  DFFR_X1 \registers_reg[15][26]  ( .D(n3056), .CK(n3891), .RN(n3309), .QN(
        n454) );
  DFFR_X1 \registers_reg[15][25]  ( .D(n3055), .CK(n3891), .RN(n3309), .QN(
        n455) );
  DFFR_X1 \registers_reg[15][24]  ( .D(n3054), .CK(n3891), .RN(n3309), .QN(
        n456) );
  DFFR_X1 \registers_reg[15][23]  ( .D(n3053), .CK(n3891), .RN(n3309), .QN(
        n457) );
  DFFR_X1 \registers_reg[15][22]  ( .D(n3052), .CK(n3891), .RN(n3309), .QN(
        n458) );
  DFFR_X1 \registers_reg[15][21]  ( .D(n3051), .CK(n3891), .RN(n3309), .QN(
        n459) );
  DFFR_X1 \registers_reg[15][20]  ( .D(n3050), .CK(n3891), .RN(n3309), .QN(
        n460) );
  DFFR_X1 \registers_reg[15][19]  ( .D(n3049), .CK(n3891), .RN(n3309), .QN(
        n461) );
  DFFR_X1 \registers_reg[15][18]  ( .D(n3048), .CK(n3891), .RN(n3309), .QN(
        n462) );
  DFFR_X1 \registers_reg[15][17]  ( .D(n3047), .CK(n3891), .RN(n3309), .QN(
        n463) );
  DFFR_X1 \registers_reg[15][16]  ( .D(n3046), .CK(n3891), .RN(n3309), .QN(
        n464) );
  DFFR_X1 \registers_reg[15][15]  ( .D(n3045), .CK(n3891), .RN(n3308), .QN(
        n465) );
  DFFR_X1 \registers_reg[15][14]  ( .D(n3044), .CK(n3891), .RN(n3308), .QN(
        n466) );
  DFFR_X1 \registers_reg[15][13]  ( .D(n3043), .CK(n3891), .RN(n3308), .QN(
        n467) );
  DFFR_X1 \registers_reg[15][12]  ( .D(n3042), .CK(n3891), .RN(n3308), .QN(
        n468) );
  DFFR_X1 \registers_reg[15][11]  ( .D(n3041), .CK(n3891), .RN(n3308), .QN(
        n469) );
  DFFR_X1 \registers_reg[15][10]  ( .D(n3040), .CK(n3891), .RN(n3308), .QN(
        n470) );
  DFFR_X1 \registers_reg[15][9]  ( .D(n3039), .CK(n3891), .RN(n3308), .QN(n471) );
  DFFR_X1 \registers_reg[15][8]  ( .D(n3038), .CK(n3891), .RN(n3308), .QN(n472) );
  DFFR_X1 \registers_reg[15][7]  ( .D(n3037), .CK(n3891), .RN(n3308), .QN(n473) );
  DFFR_X1 \registers_reg[15][6]  ( .D(n3036), .CK(n3891), .RN(n3308), .QN(n474) );
  DFFR_X1 \registers_reg[15][5]  ( .D(n3035), .CK(n3891), .RN(n3308), .QN(n475) );
  DFFR_X1 \registers_reg[15][4]  ( .D(n3034), .CK(n3891), .RN(n3307), .QN(n476) );
  DFFR_X1 \registers_reg[15][3]  ( .D(n3033), .CK(n3891), .RN(n3307), .QN(n477) );
  DFFR_X1 \registers_reg[15][2]  ( .D(n3032), .CK(n3891), .RN(n3307), .QN(n478) );
  DFFR_X1 \registers_reg[15][1]  ( .D(n3031), .CK(n3891), .RN(n3307), .QN(n479) );
  DFFR_X1 \registers_reg[15][0]  ( .D(n3030), .CK(n3891), .RN(n3307), .QN(n480) );
  DFFR_X1 \registers_reg[16][31]  ( .D(n3029), .CK(n3891), .RN(n3307), .QN(
        n481) );
  DFFR_X1 \registers_reg[16][30]  ( .D(n3028), .CK(n3891), .RN(n3307), .QN(
        n482) );
  DFFR_X1 \registers_reg[16][29]  ( .D(n3027), .CK(n3891), .RN(n3307), .QN(
        n483) );
  DFFR_X1 \registers_reg[16][28]  ( .D(n3026), .CK(n3891), .RN(n3307), .QN(
        n484) );
  DFFR_X1 \registers_reg[16][27]  ( .D(n3025), .CK(n3891), .RN(n3307), .QN(
        n485) );
  DFFR_X1 \registers_reg[16][26]  ( .D(n3024), .CK(n3891), .RN(n3307), .QN(
        n486) );
  DFFR_X1 \registers_reg[16][25]  ( .D(n3023), .CK(n3891), .RN(n3306), .QN(
        n487) );
  DFFR_X1 \registers_reg[16][24]  ( .D(n3022), .CK(n3891), .RN(n3306), .QN(
        n488) );
  DFFR_X1 \registers_reg[16][23]  ( .D(n3021), .CK(n3891), .RN(n3306), .QN(
        n489) );
  DFFR_X1 \registers_reg[16][22]  ( .D(n3020), .CK(n3891), .RN(n3306), .QN(
        n490) );
  DFFR_X1 \registers_reg[16][21]  ( .D(n3019), .CK(n3891), .RN(n3306), .QN(
        n491) );
  DFFR_X1 \registers_reg[16][20]  ( .D(n3018), .CK(n3891), .RN(n3306), .QN(
        n492) );
  DFFR_X1 \registers_reg[16][19]  ( .D(n3017), .CK(n3891), .RN(n3306), .QN(
        n493) );
  DFFR_X1 \registers_reg[16][18]  ( .D(n3016), .CK(n3891), .RN(n3306), .QN(
        n494) );
  DFFR_X1 \registers_reg[16][17]  ( .D(n3015), .CK(n3891), .RN(n3306), .QN(
        n495) );
  DFFR_X1 \registers_reg[16][16]  ( .D(n3014), .CK(n3891), .RN(n3306), .QN(
        n496) );
  DFFR_X1 \registers_reg[16][15]  ( .D(n3013), .CK(n3891), .RN(n3306), .QN(
        n497) );
  DFFR_X1 \registers_reg[16][14]  ( .D(n3012), .CK(n3891), .RN(n3305), .QN(
        n498) );
  DFFR_X1 \registers_reg[16][13]  ( .D(n3011), .CK(n3891), .RN(n3305), .QN(
        n499) );
  DFFR_X1 \registers_reg[16][12]  ( .D(n3010), .CK(n3891), .RN(n3305), .QN(
        n500) );
  DFFR_X1 \registers_reg[16][11]  ( .D(n3009), .CK(n3891), .RN(n3305), .QN(
        n501) );
  DFFR_X1 \registers_reg[16][10]  ( .D(n3008), .CK(n3891), .RN(n3305), .QN(
        n502) );
  DFFR_X1 \registers_reg[16][9]  ( .D(n3007), .CK(n3891), .RN(n3305), .QN(n503) );
  DFFR_X1 \registers_reg[16][8]  ( .D(n3006), .CK(n3891), .RN(n3305), .QN(n504) );
  DFFR_X1 \registers_reg[16][7]  ( .D(n3005), .CK(n3891), .RN(n3305), .QN(n505) );
  DFFR_X1 \registers_reg[16][6]  ( .D(n3004), .CK(n3891), .RN(n3305), .QN(n506) );
  DFFR_X1 \registers_reg[16][5]  ( .D(n3003), .CK(n3891), .RN(n3305), .QN(n507) );
  DFFR_X1 \registers_reg[16][4]  ( .D(n3002), .CK(n3891), .RN(n3305), .QN(n508) );
  DFFR_X1 \registers_reg[16][3]  ( .D(n3001), .CK(n3891), .RN(n3304), .QN(n509) );
  DFFR_X1 \registers_reg[16][2]  ( .D(n3000), .CK(n3891), .RN(n3304), .QN(n510) );
  DFFR_X1 \registers_reg[16][1]  ( .D(n2999), .CK(n3891), .RN(n3304), .QN(n511) );
  DFFR_X1 \registers_reg[16][0]  ( .D(n2998), .CK(n3891), .RN(n3304), .QN(n512) );
  DFFR_X1 \registers_reg[17][31]  ( .D(n2997), .CK(n3891), .RN(n3304), .QN(
        n513) );
  DFFR_X1 \registers_reg[17][30]  ( .D(n2996), .CK(n3891), .RN(n3304), .QN(
        n514) );
  DFFR_X1 \registers_reg[17][29]  ( .D(n2995), .CK(n3891), .RN(n3304), .QN(
        n515) );
  DFFR_X1 \registers_reg[17][28]  ( .D(n2994), .CK(n3891), .RN(n3304), .QN(
        n516) );
  DFFR_X1 \registers_reg[17][27]  ( .D(n2993), .CK(n3891), .RN(n3304), .QN(
        n517) );
  DFFR_X1 \registers_reg[17][26]  ( .D(n2992), .CK(n3891), .RN(n3304), .QN(
        n518) );
  DFFR_X1 \registers_reg[17][25]  ( .D(n2991), .CK(n3891), .RN(n3304), .QN(
        n519) );
  DFFR_X1 \registers_reg[17][24]  ( .D(n2990), .CK(n3891), .RN(n3303), .QN(
        n520) );
  DFFR_X1 \registers_reg[17][23]  ( .D(n2989), .CK(n3891), .RN(n3303), .QN(
        n521) );
  DFFR_X1 \registers_reg[17][22]  ( .D(n2988), .CK(n3891), .RN(n3303), .QN(
        n522) );
  DFFR_X1 \registers_reg[17][21]  ( .D(n2987), .CK(n3891), .RN(n3303), .QN(
        n523) );
  DFFR_X1 \registers_reg[17][20]  ( .D(n2986), .CK(n3891), .RN(n3303), .QN(
        n524) );
  DFFR_X1 \registers_reg[17][19]  ( .D(n2985), .CK(n3891), .RN(n3303), .QN(
        n525) );
  DFFR_X1 \registers_reg[17][18]  ( .D(n2984), .CK(n3891), .RN(n3303), .QN(
        n526) );
  DFFR_X1 \registers_reg[17][17]  ( .D(n2983), .CK(n3891), .RN(n3303), .QN(
        n527) );
  DFFR_X1 \registers_reg[17][16]  ( .D(n2982), .CK(n3891), .RN(n3303), .QN(
        n528) );
  DFFR_X1 \registers_reg[17][15]  ( .D(n2981), .CK(n3891), .RN(n3303), .QN(
        n529) );
  DFFR_X1 \registers_reg[17][14]  ( .D(n2980), .CK(n3891), .RN(n3303), .QN(
        n530) );
  DFFR_X1 \registers_reg[17][13]  ( .D(n2979), .CK(n3891), .RN(n3302), .QN(
        n531) );
  DFFR_X1 \registers_reg[17][12]  ( .D(n2978), .CK(n3891), .RN(n3302), .QN(
        n532) );
  DFFR_X1 \registers_reg[17][11]  ( .D(n2977), .CK(n3891), .RN(n3302), .QN(
        n533) );
  DFFR_X1 \registers_reg[17][10]  ( .D(n2976), .CK(n3891), .RN(n3302), .QN(
        n534) );
  DFFR_X1 \registers_reg[17][9]  ( .D(n2975), .CK(n3891), .RN(n3302), .QN(n535) );
  DFFR_X1 \registers_reg[17][8]  ( .D(n2974), .CK(n3891), .RN(n3302), .QN(n536) );
  DFFR_X1 \registers_reg[17][7]  ( .D(n2973), .CK(n3891), .RN(n3302), .QN(n537) );
  DFFR_X1 \registers_reg[17][6]  ( .D(n2972), .CK(n3891), .RN(n3302), .QN(n538) );
  DFFR_X1 \registers_reg[17][5]  ( .D(n2971), .CK(n3891), .RN(n3302), .QN(n539) );
  DFFR_X1 \registers_reg[17][4]  ( .D(n2970), .CK(n3891), .RN(n3302), .QN(n540) );
  DFFR_X1 \registers_reg[17][3]  ( .D(n2969), .CK(n3891), .RN(n3302), .QN(n541) );
  DFFR_X1 \registers_reg[17][2]  ( .D(n2968), .CK(n3891), .RN(n3301), .QN(n542) );
  DFFR_X1 \registers_reg[17][1]  ( .D(n2967), .CK(n3891), .RN(n3301), .QN(n543) );
  DFFR_X1 \registers_reg[17][0]  ( .D(n2966), .CK(n3891), .RN(n3301), .QN(n544) );
  DFFR_X1 \registers_reg[18][31]  ( .D(n3624), .CK(n3891), .RN(n3301), .Q(
        \registers[18][31] ) );
  DFFR_X1 \registers_reg[18][30]  ( .D(n3623), .CK(n3891), .RN(n3301), .Q(
        \registers[18][30] ) );
  DFFR_X1 \registers_reg[18][29]  ( .D(n3622), .CK(n3891), .RN(n3301), .Q(
        \registers[18][29] ) );
  DFFR_X1 \registers_reg[18][28]  ( .D(n3621), .CK(n3891), .RN(n3301), .Q(
        \registers[18][28] ) );
  DFFR_X1 \registers_reg[18][27]  ( .D(n3620), .CK(n3891), .RN(n3301), .Q(
        \registers[18][27] ) );
  DFFR_X1 \registers_reg[18][26]  ( .D(n3619), .CK(n3891), .RN(n3301), .Q(
        \registers[18][26] ) );
  DFFR_X1 \registers_reg[18][25]  ( .D(n3618), .CK(n3891), .RN(n3301), .Q(
        \registers[18][25] ) );
  DFFR_X1 \registers_reg[18][24]  ( .D(n3617), .CK(n3891), .RN(n3301), .Q(
        \registers[18][24] ) );
  DFFR_X1 \registers_reg[18][23]  ( .D(n3616), .CK(n3891), .RN(n3300), .Q(
        \registers[18][23] ) );
  DFFR_X1 \registers_reg[18][22]  ( .D(n3615), .CK(n3891), .RN(n3300), .Q(
        \registers[18][22] ) );
  DFFR_X1 \registers_reg[18][21]  ( .D(n3614), .CK(n3891), .RN(n3300), .Q(
        \registers[18][21] ) );
  DFFR_X1 \registers_reg[18][20]  ( .D(n3613), .CK(n3891), .RN(n3300), .Q(
        \registers[18][20] ) );
  DFFR_X1 \registers_reg[18][19]  ( .D(n3612), .CK(n3891), .RN(n3300), .Q(
        \registers[18][19] ) );
  DFFR_X1 \registers_reg[18][18]  ( .D(n3611), .CK(n3891), .RN(n3300), .Q(
        \registers[18][18] ) );
  DFFR_X1 \registers_reg[18][17]  ( .D(n3610), .CK(n3891), .RN(n3300), .Q(
        \registers[18][17] ) );
  DFFR_X1 \registers_reg[18][16]  ( .D(n3609), .CK(n3891), .RN(n3300), .Q(
        \registers[18][16] ) );
  DFFR_X1 \registers_reg[18][15]  ( .D(n3608), .CK(n3891), .RN(n3300), .Q(
        \registers[18][15] ) );
  DFFR_X1 \registers_reg[18][14]  ( .D(n3607), .CK(n3891), .RN(n3300), .Q(
        \registers[18][14] ) );
  DFFR_X1 \registers_reg[18][13]  ( .D(n3606), .CK(n3891), .RN(n3300), .Q(
        \registers[18][13] ) );
  DFFR_X1 \registers_reg[18][12]  ( .D(n3605), .CK(n3891), .RN(n3299), .Q(
        \registers[18][12] ) );
  DFFR_X1 \registers_reg[18][11]  ( .D(n3604), .CK(n3891), .RN(n3299), .Q(
        \registers[18][11] ) );
  DFFR_X1 \registers_reg[18][10]  ( .D(n3603), .CK(n3891), .RN(n3299), .Q(
        \registers[18][10] ) );
  DFFR_X1 \registers_reg[18][9]  ( .D(n3602), .CK(n3891), .RN(n3299), .Q(
        \registers[18][9] ) );
  DFFR_X1 \registers_reg[18][8]  ( .D(n3601), .CK(n3891), .RN(n3299), .Q(
        \registers[18][8] ) );
  DFFR_X1 \registers_reg[18][7]  ( .D(n3600), .CK(n3891), .RN(n3299), .Q(
        \registers[18][7] ) );
  DFFR_X1 \registers_reg[18][6]  ( .D(n3599), .CK(n3891), .RN(n3299), .Q(
        \registers[18][6] ) );
  DFFR_X1 \registers_reg[18][5]  ( .D(n3598), .CK(n3891), .RN(n3299), .Q(
        \registers[18][5] ) );
  DFFR_X1 \registers_reg[18][4]  ( .D(n3597), .CK(n3891), .RN(n3299), .Q(
        \registers[18][4] ) );
  DFFR_X1 \registers_reg[18][3]  ( .D(n3596), .CK(n3891), .RN(n3299), .Q(
        \registers[18][3] ) );
  DFFR_X1 \registers_reg[18][2]  ( .D(n3595), .CK(n3891), .RN(n3299), .Q(
        \registers[18][2] ) );
  DFFR_X1 \registers_reg[18][1]  ( .D(n3594), .CK(n3891), .RN(n3298), .Q(
        \registers[18][1] ) );
  DFFR_X1 \registers_reg[18][0]  ( .D(n3593), .CK(n3891), .RN(n3298), .Q(
        \registers[18][0] ) );
  DFFR_X1 \registers_reg[19][31]  ( .D(n3656), .CK(n3891), .RN(n3298), .Q(
        \registers[19][31] ) );
  DFFR_X1 \registers_reg[19][30]  ( .D(n3655), .CK(n3891), .RN(n3298), .Q(
        \registers[19][30] ) );
  DFFR_X1 \registers_reg[19][29]  ( .D(n3654), .CK(n3891), .RN(n3298), .Q(
        \registers[19][29] ) );
  DFFR_X1 \registers_reg[19][28]  ( .D(n3653), .CK(n3891), .RN(n3298), .Q(
        \registers[19][28] ) );
  DFFR_X1 \registers_reg[19][27]  ( .D(n3652), .CK(n3891), .RN(n3298), .Q(
        \registers[19][27] ) );
  DFFR_X1 \registers_reg[19][26]  ( .D(n3651), .CK(n3891), .RN(n3298), .Q(
        \registers[19][26] ) );
  DFFR_X1 \registers_reg[19][25]  ( .D(n3650), .CK(n3891), .RN(n3298), .Q(
        \registers[19][25] ) );
  DFFR_X1 \registers_reg[19][24]  ( .D(n3649), .CK(n3891), .RN(n3298), .Q(
        \registers[19][24] ) );
  DFFR_X1 \registers_reg[19][23]  ( .D(n3648), .CK(n3891), .RN(n3298), .Q(
        \registers[19][23] ) );
  DFFR_X1 \registers_reg[19][22]  ( .D(n3647), .CK(n3891), .RN(n3297), .Q(
        \registers[19][22] ) );
  DFFR_X1 \registers_reg[19][21]  ( .D(n3646), .CK(n3891), .RN(n3297), .Q(
        \registers[19][21] ) );
  DFFR_X1 \registers_reg[19][20]  ( .D(n3645), .CK(n3891), .RN(n3297), .Q(
        \registers[19][20] ) );
  DFFR_X1 \registers_reg[19][19]  ( .D(n3644), .CK(n3891), .RN(n3297), .Q(
        \registers[19][19] ) );
  DFFR_X1 \registers_reg[19][18]  ( .D(n3643), .CK(n3891), .RN(n3297), .Q(
        \registers[19][18] ) );
  DFFR_X1 \registers_reg[19][17]  ( .D(n3642), .CK(n3891), .RN(n3297), .Q(
        \registers[19][17] ) );
  DFFR_X1 \registers_reg[19][16]  ( .D(n3641), .CK(n3891), .RN(n3297), .Q(
        \registers[19][16] ) );
  DFFR_X1 \registers_reg[19][15]  ( .D(n3640), .CK(n3891), .RN(n3297), .Q(
        \registers[19][15] ) );
  DFFR_X1 \registers_reg[19][14]  ( .D(n3639), .CK(n3891), .RN(n3297), .Q(
        \registers[19][14] ) );
  DFFR_X1 \registers_reg[19][13]  ( .D(n3638), .CK(n3891), .RN(n3297), .Q(
        \registers[19][13] ) );
  DFFR_X1 \registers_reg[19][12]  ( .D(n3637), .CK(n3891), .RN(n3297), .Q(
        \registers[19][12] ) );
  DFFR_X1 \registers_reg[19][11]  ( .D(n3636), .CK(n3891), .RN(n3296), .Q(
        \registers[19][11] ) );
  DFFR_X1 \registers_reg[19][10]  ( .D(n3635), .CK(n3891), .RN(n3296), .Q(
        \registers[19][10] ) );
  DFFR_X1 \registers_reg[19][9]  ( .D(n3634), .CK(n3891), .RN(n3296), .Q(
        \registers[19][9] ) );
  DFFR_X1 \registers_reg[19][8]  ( .D(n3633), .CK(n3891), .RN(n3296), .Q(
        \registers[19][8] ) );
  DFFR_X1 \registers_reg[19][7]  ( .D(n3632), .CK(n3891), .RN(n3296), .Q(
        \registers[19][7] ) );
  DFFR_X1 \registers_reg[19][6]  ( .D(n3631), .CK(n3891), .RN(n3296), .Q(
        \registers[19][6] ) );
  DFFR_X1 \registers_reg[19][5]  ( .D(n3630), .CK(n3891), .RN(n3296), .Q(
        \registers[19][5] ) );
  DFFR_X1 \registers_reg[19][4]  ( .D(n3629), .CK(n3891), .RN(n3296), .Q(
        \registers[19][4] ) );
  DFFR_X1 \registers_reg[19][3]  ( .D(n3628), .CK(n3891), .RN(n3296), .Q(
        \registers[19][3] ) );
  DFFR_X1 \registers_reg[19][2]  ( .D(n3627), .CK(n3891), .RN(n3296), .Q(
        \registers[19][2] ) );
  DFFR_X1 \registers_reg[19][1]  ( .D(n3626), .CK(n3891), .RN(n3296), .Q(
        \registers[19][1] ) );
  DFFR_X1 \registers_reg[19][0]  ( .D(n3625), .CK(n3891), .RN(n3295), .Q(
        \registers[19][0] ) );
  DFFR_X1 \registers_reg[20][31]  ( .D(n2965), .CK(n3891), .RN(n3295), .QN(
        n609) );
  DFFR_X1 \registers_reg[20][30]  ( .D(n2964), .CK(n3891), .RN(n3295), .QN(
        n610) );
  DFFR_X1 \registers_reg[20][29]  ( .D(n2963), .CK(n3891), .RN(n3295), .QN(
        n611) );
  DFFR_X1 \registers_reg[20][28]  ( .D(n2962), .CK(n3891), .RN(n3295), .QN(
        n612) );
  DFFR_X1 \registers_reg[20][27]  ( .D(n2961), .CK(n3891), .RN(n3295), .QN(
        n613) );
  DFFR_X1 \registers_reg[20][26]  ( .D(n2960), .CK(n3891), .RN(n3295), .QN(
        n614) );
  DFFR_X1 \registers_reg[20][25]  ( .D(n2959), .CK(n3891), .RN(n3295), .QN(
        n615) );
  DFFR_X1 \registers_reg[20][24]  ( .D(n2958), .CK(n3891), .RN(n3295), .QN(
        n616) );
  DFFR_X1 \registers_reg[20][23]  ( .D(n2957), .CK(n3891), .RN(n3295), .QN(
        n617) );
  DFFR_X1 \registers_reg[20][22]  ( .D(n2956), .CK(n3891), .RN(n3295), .QN(
        n618) );
  DFFR_X1 \registers_reg[20][21]  ( .D(n2955), .CK(n3891), .RN(n3294), .QN(
        n619) );
  DFFR_X1 \registers_reg[20][20]  ( .D(n2954), .CK(n3891), .RN(n3294), .QN(
        n620) );
  DFFR_X1 \registers_reg[20][19]  ( .D(n2953), .CK(n3891), .RN(n3294), .QN(
        n621) );
  DFFR_X1 \registers_reg[20][18]  ( .D(n2952), .CK(n3891), .RN(n3294), .QN(
        n622) );
  DFFR_X1 \registers_reg[20][17]  ( .D(n2951), .CK(n3891), .RN(n3294), .QN(
        n623) );
  DFFR_X1 \registers_reg[20][16]  ( .D(n2950), .CK(n3891), .RN(n3294), .QN(
        n624) );
  DFFR_X1 \registers_reg[20][15]  ( .D(n2949), .CK(n3891), .RN(n3294), .QN(
        n625) );
  DFFR_X1 \registers_reg[20][14]  ( .D(n2948), .CK(n3891), .RN(n3294), .QN(
        n626) );
  DFFR_X1 \registers_reg[20][13]  ( .D(n2947), .CK(n3891), .RN(n3294), .QN(
        n627) );
  DFFR_X1 \registers_reg[20][12]  ( .D(n2946), .CK(n3891), .RN(n3294), .QN(
        n628) );
  DFFR_X1 \registers_reg[20][11]  ( .D(n2945), .CK(n3891), .RN(n3294), .QN(
        n629) );
  DFFR_X1 \registers_reg[20][10]  ( .D(n2944), .CK(n3891), .RN(n3293), .QN(
        n630) );
  DFFR_X1 \registers_reg[20][9]  ( .D(n2943), .CK(n3891), .RN(n3293), .QN(n631) );
  DFFR_X1 \registers_reg[20][8]  ( .D(n2942), .CK(n3891), .RN(n3293), .QN(n632) );
  DFFR_X1 \registers_reg[20][7]  ( .D(n2941), .CK(n3891), .RN(n3293), .QN(n633) );
  DFFR_X1 \registers_reg[20][6]  ( .D(n2940), .CK(n3891), .RN(n3293), .QN(n634) );
  DFFR_X1 \registers_reg[20][5]  ( .D(n2939), .CK(n3891), .RN(n3293), .QN(n635) );
  DFFR_X1 \registers_reg[20][4]  ( .D(n2938), .CK(n3891), .RN(n3293), .QN(n636) );
  DFFR_X1 \registers_reg[20][3]  ( .D(n2937), .CK(n3891), .RN(n3293), .QN(n637) );
  DFFR_X1 \registers_reg[20][2]  ( .D(n2936), .CK(n3891), .RN(n3293), .QN(n638) );
  DFFR_X1 \registers_reg[20][1]  ( .D(n2935), .CK(n3891), .RN(n3293), .QN(n639) );
  DFFR_X1 \registers_reg[20][0]  ( .D(n2934), .CK(n3891), .RN(n3293), .QN(n640) );
  DFFR_X1 \registers_reg[21][31]  ( .D(n2933), .CK(n3891), .RN(n3292), .QN(
        n641) );
  DFFR_X1 \registers_reg[21][30]  ( .D(n2932), .CK(n3891), .RN(n3292), .QN(
        n642) );
  DFFR_X1 \registers_reg[21][29]  ( .D(n2931), .CK(n3891), .RN(n3292), .QN(
        n643) );
  DFFR_X1 \registers_reg[21][28]  ( .D(n2930), .CK(n3891), .RN(n3292), .QN(
        n644) );
  DFFR_X1 \registers_reg[21][27]  ( .D(n2929), .CK(n3891), .RN(n3292), .QN(
        n645) );
  DFFR_X1 \registers_reg[21][26]  ( .D(n2928), .CK(n3891), .RN(n3292), .QN(
        n646) );
  DFFR_X1 \registers_reg[21][25]  ( .D(n2927), .CK(n3891), .RN(n3292), .QN(
        n647) );
  DFFR_X1 \registers_reg[21][24]  ( .D(n2926), .CK(n3891), .RN(n3292), .QN(
        n648) );
  DFFR_X1 \registers_reg[21][23]  ( .D(n2925), .CK(n3891), .RN(n3292), .QN(
        n649) );
  DFFR_X1 \registers_reg[21][22]  ( .D(n2924), .CK(n3891), .RN(n3292), .QN(
        n650) );
  DFFR_X1 \registers_reg[21][21]  ( .D(n2923), .CK(n3891), .RN(n3292), .QN(
        n651) );
  DFFR_X1 \registers_reg[21][20]  ( .D(n2922), .CK(n3891), .RN(n3291), .QN(
        n652) );
  DFFR_X1 \registers_reg[21][19]  ( .D(n2921), .CK(n3891), .RN(n3291), .QN(
        n653) );
  DFFR_X1 \registers_reg[21][18]  ( .D(n2920), .CK(n3891), .RN(n3291), .QN(
        n654) );
  DFFR_X1 \registers_reg[21][17]  ( .D(n2919), .CK(n3891), .RN(n3291), .QN(
        n655) );
  DFFR_X1 \registers_reg[21][16]  ( .D(n2918), .CK(n3891), .RN(n3291), .QN(
        n656) );
  DFFR_X1 \registers_reg[21][15]  ( .D(n2917), .CK(n3891), .RN(n3291), .QN(
        n657) );
  DFFR_X1 \registers_reg[21][14]  ( .D(n2916), .CK(n3891), .RN(n3291), .QN(
        n658) );
  DFFR_X1 \registers_reg[21][13]  ( .D(n2915), .CK(n3891), .RN(n3291), .QN(
        n659) );
  DFFR_X1 \registers_reg[21][12]  ( .D(n2914), .CK(n3891), .RN(n3291), .QN(
        n660) );
  DFFR_X1 \registers_reg[21][11]  ( .D(n2913), .CK(n3891), .RN(n3291), .QN(
        n661) );
  DFFR_X1 \registers_reg[21][10]  ( .D(n2912), .CK(n3891), .RN(n3291), .QN(
        n662) );
  DFFR_X1 \registers_reg[21][9]  ( .D(n2911), .CK(n3891), .RN(n3290), .QN(n663) );
  DFFR_X1 \registers_reg[21][8]  ( .D(n2910), .CK(n3891), .RN(n3290), .QN(n664) );
  DFFR_X1 \registers_reg[21][7]  ( .D(n2909), .CK(n3891), .RN(n3290), .QN(n665) );
  DFFR_X1 \registers_reg[21][6]  ( .D(n2908), .CK(n3891), .RN(n3290), .QN(n666) );
  DFFR_X1 \registers_reg[21][5]  ( .D(n2907), .CK(n3891), .RN(n3290), .QN(n667) );
  DFFR_X1 \registers_reg[21][4]  ( .D(n2906), .CK(n3891), .RN(n3290), .QN(n668) );
  DFFR_X1 \registers_reg[21][3]  ( .D(n2905), .CK(n3891), .RN(n3290), .QN(n669) );
  DFFR_X1 \registers_reg[21][2]  ( .D(n2904), .CK(n3891), .RN(n3290), .QN(n670) );
  DFFR_X1 \registers_reg[21][1]  ( .D(n2903), .CK(n3891), .RN(n3290), .QN(n671) );
  DFFR_X1 \registers_reg[21][0]  ( .D(n2902), .CK(n3891), .RN(n3290), .QN(n672) );
  DFFR_X1 \registers_reg[22][31]  ( .D(n3688), .CK(n3891), .RN(n3290), .Q(
        \registers[22][31] ) );
  DFFR_X1 \registers_reg[22][30]  ( .D(n3687), .CK(n3891), .RN(n3289), .Q(
        \registers[22][30] ) );
  DFFR_X1 \registers_reg[22][29]  ( .D(n3686), .CK(n3891), .RN(n3289), .Q(
        \registers[22][29] ) );
  DFFR_X1 \registers_reg[22][28]  ( .D(n3685), .CK(n3891), .RN(n3289), .Q(
        \registers[22][28] ) );
  DFFR_X1 \registers_reg[22][27]  ( .D(n3684), .CK(n3891), .RN(n3289), .Q(
        \registers[22][27] ) );
  DFFR_X1 \registers_reg[22][26]  ( .D(n3683), .CK(n3891), .RN(n3289), .Q(
        \registers[22][26] ) );
  DFFR_X1 \registers_reg[22][25]  ( .D(n3682), .CK(n3891), .RN(n3289), .Q(
        \registers[22][25] ) );
  DFFR_X1 \registers_reg[22][24]  ( .D(n3681), .CK(n3891), .RN(n3289), .Q(
        \registers[22][24] ) );
  DFFR_X1 \registers_reg[22][23]  ( .D(n3680), .CK(n3891), .RN(n3289), .Q(
        \registers[22][23] ) );
  DFFR_X1 \registers_reg[22][22]  ( .D(n3679), .CK(n3891), .RN(n3289), .Q(
        \registers[22][22] ) );
  DFFR_X1 \registers_reg[22][21]  ( .D(n3678), .CK(n3891), .RN(n3289), .Q(
        \registers[22][21] ) );
  DFFR_X1 \registers_reg[22][20]  ( .D(n3677), .CK(n3891), .RN(n3289), .Q(
        \registers[22][20] ) );
  DFFR_X1 \registers_reg[22][19]  ( .D(n3676), .CK(n3891), .RN(n3288), .Q(
        \registers[22][19] ) );
  DFFR_X1 \registers_reg[22][18]  ( .D(n3675), .CK(n3891), .RN(n3288), .Q(
        \registers[22][18] ) );
  DFFR_X1 \registers_reg[22][17]  ( .D(n3674), .CK(n3891), .RN(n3288), .Q(
        \registers[22][17] ) );
  DFFR_X1 \registers_reg[22][16]  ( .D(n3673), .CK(n3891), .RN(n3288), .Q(
        \registers[22][16] ) );
  DFFR_X1 \registers_reg[22][15]  ( .D(n3672), .CK(n3891), .RN(n3288), .Q(
        \registers[22][15] ) );
  DFFR_X1 \registers_reg[22][14]  ( .D(n3671), .CK(n3891), .RN(n3288), .Q(
        \registers[22][14] ) );
  DFFR_X1 \registers_reg[22][13]  ( .D(n3670), .CK(n3891), .RN(n3288), .Q(
        \registers[22][13] ) );
  DFFR_X1 \registers_reg[22][12]  ( .D(n3669), .CK(n3891), .RN(n3288), .Q(
        \registers[22][12] ) );
  DFFR_X1 \registers_reg[22][11]  ( .D(n3668), .CK(n3891), .RN(n3288), .Q(
        \registers[22][11] ) );
  DFFR_X1 \registers_reg[22][10]  ( .D(n3667), .CK(n3891), .RN(n3288), .Q(
        \registers[22][10] ) );
  DFFR_X1 \registers_reg[22][9]  ( .D(n3666), .CK(n3891), .RN(n3288), .Q(
        \registers[22][9] ) );
  DFFR_X1 \registers_reg[22][8]  ( .D(n3665), .CK(n3891), .RN(n3287), .Q(
        \registers[22][8] ) );
  DFFR_X1 \registers_reg[22][7]  ( .D(n3664), .CK(n3891), .RN(n3287), .Q(
        \registers[22][7] ) );
  DFFR_X1 \registers_reg[22][6]  ( .D(n3663), .CK(n3891), .RN(n3287), .Q(
        \registers[22][6] ) );
  DFFR_X1 \registers_reg[22][5]  ( .D(n3662), .CK(n3891), .RN(n3287), .Q(
        \registers[22][5] ) );
  DFFR_X1 \registers_reg[22][4]  ( .D(n3661), .CK(n3891), .RN(n3287), .Q(
        \registers[22][4] ) );
  DFFR_X1 \registers_reg[22][3]  ( .D(n3660), .CK(n3891), .RN(n3287), .Q(
        \registers[22][3] ) );
  DFFR_X1 \registers_reg[22][2]  ( .D(n3659), .CK(n3891), .RN(n3287), .Q(
        \registers[22][2] ) );
  DFFR_X1 \registers_reg[22][1]  ( .D(n3658), .CK(n3891), .RN(n3287), .Q(
        \registers[22][1] ) );
  DFFR_X1 \registers_reg[22][0]  ( .D(n3657), .CK(n3891), .RN(n3287), .Q(
        \registers[22][0] ) );
  DFFR_X1 \registers_reg[23][31]  ( .D(n3720), .CK(n3891), .RN(n3287), .Q(
        \registers[23][31] ) );
  DFFR_X1 \registers_reg[23][30]  ( .D(n3719), .CK(n3891), .RN(n3287), .Q(
        \registers[23][30] ) );
  DFFR_X1 \registers_reg[23][29]  ( .D(n3718), .CK(n3891), .RN(n3286), .Q(
        \registers[23][29] ) );
  DFFR_X1 \registers_reg[23][28]  ( .D(n3717), .CK(n3891), .RN(n3286), .Q(
        \registers[23][28] ) );
  DFFR_X1 \registers_reg[23][27]  ( .D(n3716), .CK(n3891), .RN(n3286), .Q(
        \registers[23][27] ) );
  DFFR_X1 \registers_reg[23][26]  ( .D(n3715), .CK(n3891), .RN(n3286), .Q(
        \registers[23][26] ) );
  DFFR_X1 \registers_reg[23][25]  ( .D(n3714), .CK(n3891), .RN(n3286), .Q(
        \registers[23][25] ) );
  DFFR_X1 \registers_reg[23][24]  ( .D(n3713), .CK(n3891), .RN(n3286), .Q(
        \registers[23][24] ) );
  DFFR_X1 \registers_reg[23][23]  ( .D(n3712), .CK(n3891), .RN(n3286), .Q(
        \registers[23][23] ) );
  DFFR_X1 \registers_reg[23][22]  ( .D(n3711), .CK(n3891), .RN(n3286), .Q(
        \registers[23][22] ) );
  DFFR_X1 \registers_reg[23][21]  ( .D(n3710), .CK(n3891), .RN(n3286), .Q(
        \registers[23][21] ) );
  DFFR_X1 \registers_reg[23][20]  ( .D(n3709), .CK(n3891), .RN(n3286), .Q(
        \registers[23][20] ) );
  DFFR_X1 \registers_reg[23][19]  ( .D(n3708), .CK(n3891), .RN(n3286), .Q(
        \registers[23][19] ) );
  DFFR_X1 \registers_reg[23][18]  ( .D(n3707), .CK(n3891), .RN(n1067), .Q(
        \registers[23][18] ) );
  DFFR_X1 \registers_reg[23][17]  ( .D(n3706), .CK(n3891), .RN(n1067), .Q(
        \registers[23][17] ) );
  DFFR_X1 \registers_reg[23][16]  ( .D(n3705), .CK(n3891), .RN(n1067), .Q(
        \registers[23][16] ) );
  DFFR_X1 \registers_reg[23][15]  ( .D(n3704), .CK(n3891), .RN(n1067), .Q(
        \registers[23][15] ) );
  DFFR_X1 \registers_reg[23][14]  ( .D(n3703), .CK(n3891), .RN(n1067), .Q(
        \registers[23][14] ) );
  DFFR_X1 \registers_reg[23][13]  ( .D(n3702), .CK(n3891), .RN(n1067), .Q(
        \registers[23][13] ) );
  DFFR_X1 \registers_reg[23][12]  ( .D(n3701), .CK(n3891), .RN(n1067), .Q(
        \registers[23][12] ) );
  DFFR_X1 \registers_reg[23][11]  ( .D(n3700), .CK(n3891), .RN(n1067), .Q(
        \registers[23][11] ) );
  DFFR_X1 \registers_reg[23][10]  ( .D(n3699), .CK(n3891), .RN(n1067), .Q(
        \registers[23][10] ) );
  DFFR_X1 \registers_reg[23][9]  ( .D(n3698), .CK(n3891), .RN(n1067), .Q(
        \registers[23][9] ) );
  DFFR_X1 \registers_reg[23][8]  ( .D(n3697), .CK(n3891), .RN(n1067), .Q(
        \registers[23][8] ) );
  DFFR_X1 \registers_reg[23][7]  ( .D(n3696), .CK(n3891), .RN(n1066), .Q(
        \registers[23][7] ) );
  DFFR_X1 \registers_reg[23][6]  ( .D(n3695), .CK(n3891), .RN(n1066), .Q(
        \registers[23][6] ) );
  DFFR_X1 \registers_reg[23][5]  ( .D(n3694), .CK(n3891), .RN(n1066), .Q(
        \registers[23][5] ) );
  DFFR_X1 \registers_reg[23][4]  ( .D(n3693), .CK(n3891), .RN(n1066), .Q(
        \registers[23][4] ) );
  DFFR_X1 \registers_reg[23][3]  ( .D(n3692), .CK(n3891), .RN(n1066), .Q(
        \registers[23][3] ) );
  DFFR_X1 \registers_reg[23][2]  ( .D(n3691), .CK(n3891), .RN(n1066), .Q(
        \registers[23][2] ) );
  DFFR_X1 \registers_reg[23][1]  ( .D(n3690), .CK(n3891), .RN(n1066), .Q(
        \registers[23][1] ) );
  DFFR_X1 \registers_reg[23][0]  ( .D(n3689), .CK(n3891), .RN(n1066), .Q(
        \registers[23][0] ) );
  DFFR_X1 \registers_reg[24][31]  ( .D(n3752), .CK(n3891), .RN(n1066), .Q(
        \registers[24][31] ) );
  DFFR_X1 \registers_reg[24][30]  ( .D(n3751), .CK(n3891), .RN(n1066), .Q(
        \registers[24][30] ) );
  DFFR_X1 \registers_reg[24][29]  ( .D(n3750), .CK(n3891), .RN(n1066), .Q(
        \registers[24][29] ) );
  DFFR_X1 \registers_reg[24][28]  ( .D(n3749), .CK(n3891), .RN(n1065), .Q(
        \registers[24][28] ) );
  DFFR_X1 \registers_reg[24][27]  ( .D(n3748), .CK(n3891), .RN(n1065), .Q(
        \registers[24][27] ) );
  DFFR_X1 \registers_reg[24][26]  ( .D(n3747), .CK(n3891), .RN(n1065), .Q(
        \registers[24][26] ) );
  DFFR_X1 \registers_reg[24][25]  ( .D(n3746), .CK(n3891), .RN(n1065), .Q(
        \registers[24][25] ) );
  DFFR_X1 \registers_reg[24][24]  ( .D(n3745), .CK(n3891), .RN(n1065), .Q(
        \registers[24][24] ) );
  DFFR_X1 \registers_reg[24][23]  ( .D(n3744), .CK(n3891), .RN(n1065), .Q(
        \registers[24][23] ) );
  DFFR_X1 \registers_reg[24][22]  ( .D(n3743), .CK(n3891), .RN(n1065), .Q(
        \registers[24][22] ) );
  DFFR_X1 \registers_reg[24][21]  ( .D(n3742), .CK(n3891), .RN(n1065), .Q(
        \registers[24][21] ) );
  DFFR_X1 \registers_reg[24][20]  ( .D(n3741), .CK(n3891), .RN(n1065), .Q(
        \registers[24][20] ) );
  DFFR_X1 \registers_reg[24][19]  ( .D(n3740), .CK(n3891), .RN(n1065), .Q(
        \registers[24][19] ) );
  DFFR_X1 \registers_reg[24][18]  ( .D(n3739), .CK(n3891), .RN(n1065), .Q(
        \registers[24][18] ) );
  DFFR_X1 \registers_reg[24][17]  ( .D(n3738), .CK(n3891), .RN(n1064), .Q(
        \registers[24][17] ) );
  DFFR_X1 \registers_reg[24][16]  ( .D(n3737), .CK(n3891), .RN(n1064), .Q(
        \registers[24][16] ) );
  DFFR_X1 \registers_reg[24][15]  ( .D(n3736), .CK(n3891), .RN(n1064), .Q(
        \registers[24][15] ) );
  DFFR_X1 \registers_reg[24][14]  ( .D(n3735), .CK(n3891), .RN(n1064), .Q(
        \registers[24][14] ) );
  DFFR_X1 \registers_reg[24][13]  ( .D(n3734), .CK(n3891), .RN(n1064), .Q(
        \registers[24][13] ) );
  DFFR_X1 \registers_reg[24][12]  ( .D(n3733), .CK(n3891), .RN(n1064), .Q(
        \registers[24][12] ) );
  DFFR_X1 \registers_reg[24][11]  ( .D(n3732), .CK(n3891), .RN(n1064), .Q(
        \registers[24][11] ) );
  DFFR_X1 \registers_reg[24][10]  ( .D(n3731), .CK(n3891), .RN(n1064), .Q(
        \registers[24][10] ) );
  DFFR_X1 \registers_reg[24][9]  ( .D(n3730), .CK(n3891), .RN(n1064), .Q(
        \registers[24][9] ) );
  DFFR_X1 \registers_reg[24][8]  ( .D(n3729), .CK(n3891), .RN(n1064), .Q(
        \registers[24][8] ) );
  DFFR_X1 \registers_reg[24][7]  ( .D(n3728), .CK(n3891), .RN(n1064), .Q(
        \registers[24][7] ) );
  DFFR_X1 \registers_reg[24][6]  ( .D(n3727), .CK(n3891), .RN(n1063), .Q(
        \registers[24][6] ) );
  DFFR_X1 \registers_reg[24][5]  ( .D(n3726), .CK(n3891), .RN(n1063), .Q(
        \registers[24][5] ) );
  DFFR_X1 \registers_reg[24][4]  ( .D(n3725), .CK(n3891), .RN(n1063), .Q(
        \registers[24][4] ) );
  DFFR_X1 \registers_reg[24][3]  ( .D(n3724), .CK(n3891), .RN(n1063), .Q(
        \registers[24][3] ) );
  DFFR_X1 \registers_reg[24][2]  ( .D(n3723), .CK(n3891), .RN(n1063), .Q(
        \registers[24][2] ) );
  DFFR_X1 \registers_reg[24][1]  ( .D(n3722), .CK(n3891), .RN(n1063), .Q(
        \registers[24][1] ) );
  DFFR_X1 \registers_reg[24][0]  ( .D(n3721), .CK(n3891), .RN(n1063), .Q(
        \registers[24][0] ) );
  DFFR_X1 \registers_reg[25][31]  ( .D(n3784), .CK(n3891), .RN(n1063), .Q(
        \registers[25][31] ) );
  DFFR_X1 \registers_reg[25][30]  ( .D(n3783), .CK(n3891), .RN(n1063), .Q(
        \registers[25][30] ) );
  DFFR_X1 \registers_reg[25][29]  ( .D(n3782), .CK(n3891), .RN(n1063), .Q(
        \registers[25][29] ) );
  DFFR_X1 \registers_reg[25][28]  ( .D(n3781), .CK(n3891), .RN(n1063), .Q(
        \registers[25][28] ) );
  DFFR_X1 \registers_reg[25][27]  ( .D(n3780), .CK(n3891), .RN(n1062), .Q(
        \registers[25][27] ) );
  DFFR_X1 \registers_reg[25][26]  ( .D(n3779), .CK(n3891), .RN(n1062), .Q(
        \registers[25][26] ) );
  DFFR_X1 \registers_reg[25][25]  ( .D(n3778), .CK(n3891), .RN(n1062), .Q(
        \registers[25][25] ) );
  DFFR_X1 \registers_reg[25][24]  ( .D(n3777), .CK(n3891), .RN(n1062), .Q(
        \registers[25][24] ) );
  DFFR_X1 \registers_reg[25][23]  ( .D(n3776), .CK(n3891), .RN(n1062), .Q(
        \registers[25][23] ) );
  DFFR_X1 \registers_reg[25][22]  ( .D(n3775), .CK(n3891), .RN(n1062), .Q(
        \registers[25][22] ) );
  DFFR_X1 \registers_reg[25][21]  ( .D(n3774), .CK(n3891), .RN(n1062), .Q(
        \registers[25][21] ) );
  DFFR_X1 \registers_reg[25][20]  ( .D(n3773), .CK(n3891), .RN(n1062), .Q(
        \registers[25][20] ) );
  DFFR_X1 \registers_reg[25][19]  ( .D(n3772), .CK(n3891), .RN(n1062), .Q(
        \registers[25][19] ) );
  DFFR_X1 \registers_reg[25][18]  ( .D(n3771), .CK(n3891), .RN(n1062), .Q(
        \registers[25][18] ) );
  DFFR_X1 \registers_reg[25][17]  ( .D(n3770), .CK(n3891), .RN(n1062), .Q(
        \registers[25][17] ) );
  DFFR_X1 \registers_reg[25][16]  ( .D(n3769), .CK(n3891), .RN(n1061), .Q(
        \registers[25][16] ) );
  DFFR_X1 \registers_reg[25][15]  ( .D(n3768), .CK(n3891), .RN(n1061), .Q(
        \registers[25][15] ) );
  DFFR_X1 \registers_reg[25][14]  ( .D(n3767), .CK(n3891), .RN(n1061), .Q(
        \registers[25][14] ) );
  DFFR_X1 \registers_reg[25][13]  ( .D(n3766), .CK(n3891), .RN(n1061), .Q(
        \registers[25][13] ) );
  DFFR_X1 \registers_reg[25][12]  ( .D(n3765), .CK(n3891), .RN(n1061), .Q(
        \registers[25][12] ) );
  DFFR_X1 \registers_reg[25][11]  ( .D(n3764), .CK(n3891), .RN(n1061), .Q(
        \registers[25][11] ) );
  DFFR_X1 \registers_reg[25][10]  ( .D(n3763), .CK(n3891), .RN(n1061), .Q(
        \registers[25][10] ) );
  DFFR_X1 \registers_reg[25][9]  ( .D(n3762), .CK(n3891), .RN(n1061), .Q(
        \registers[25][9] ) );
  DFFR_X1 \registers_reg[25][8]  ( .D(n3761), .CK(n3891), .RN(n1061), .Q(
        \registers[25][8] ) );
  DFFR_X1 \registers_reg[25][7]  ( .D(n3760), .CK(n3891), .RN(n1061), .Q(
        \registers[25][7] ) );
  DFFR_X1 \registers_reg[25][6]  ( .D(n3759), .CK(n3891), .RN(n1061), .Q(
        \registers[25][6] ) );
  DFFR_X1 \registers_reg[25][5]  ( .D(n3758), .CK(n3891), .RN(n1060), .Q(
        \registers[25][5] ) );
  DFFR_X1 \registers_reg[25][4]  ( .D(n3757), .CK(n3891), .RN(n1060), .Q(
        \registers[25][4] ) );
  DFFR_X1 \registers_reg[25][3]  ( .D(n3756), .CK(n3891), .RN(n1060), .Q(
        \registers[25][3] ) );
  DFFR_X1 \registers_reg[25][2]  ( .D(n3755), .CK(n3891), .RN(n1060), .Q(
        \registers[25][2] ) );
  DFFR_X1 \registers_reg[25][1]  ( .D(n3754), .CK(n3891), .RN(n1060), .Q(
        \registers[25][1] ) );
  DFFR_X1 \registers_reg[25][0]  ( .D(n3753), .CK(n3891), .RN(n1060), .Q(
        \registers[25][0] ) );
  DFFR_X1 \registers_reg[26][31]  ( .D(n2901), .CK(n3891), .RN(n1060), .QN(
        n801) );
  DFFR_X1 \registers_reg[26][30]  ( .D(n2900), .CK(n3891), .RN(n1060), .QN(
        n802) );
  DFFR_X1 \registers_reg[26][29]  ( .D(n2899), .CK(n3891), .RN(n1060), .QN(
        n803) );
  DFFR_X1 \registers_reg[26][28]  ( .D(n2898), .CK(n3891), .RN(n1060), .QN(
        n804) );
  DFFR_X1 \registers_reg[26][27]  ( .D(n2897), .CK(n3891), .RN(n1060), .QN(
        n805) );
  DFFR_X1 \registers_reg[26][26]  ( .D(n2896), .CK(n3891), .RN(n1059), .QN(
        n806) );
  DFFR_X1 \registers_reg[26][25]  ( .D(n2895), .CK(n3891), .RN(n1059), .QN(
        n807) );
  DFFR_X1 \registers_reg[26][24]  ( .D(n2894), .CK(n3891), .RN(n1059), .QN(
        n808) );
  DFFR_X1 \registers_reg[26][23]  ( .D(n2893), .CK(n3891), .RN(n1059), .QN(
        n809) );
  DFFR_X1 \registers_reg[26][22]  ( .D(n2892), .CK(n3891), .RN(n1059), .QN(
        n810) );
  DFFR_X1 \registers_reg[26][21]  ( .D(n2891), .CK(n3891), .RN(n1059), .QN(
        n811) );
  DFFR_X1 \registers_reg[26][20]  ( .D(n2890), .CK(n3891), .RN(n1059), .QN(
        n812) );
  DFFR_X1 \registers_reg[26][19]  ( .D(n2889), .CK(n3891), .RN(n1059), .QN(
        n813) );
  DFFR_X1 \registers_reg[26][18]  ( .D(n2888), .CK(n3891), .RN(n1059), .QN(
        n814) );
  DFFR_X1 \registers_reg[26][17]  ( .D(n2887), .CK(n3891), .RN(n1059), .QN(
        n815) );
  DFFR_X1 \registers_reg[26][16]  ( .D(n2886), .CK(n3891), .RN(n1059), .QN(
        n816) );
  DFFR_X1 \registers_reg[26][15]  ( .D(n2885), .CK(n3891), .RN(n1058), .QN(
        n817) );
  DFFR_X1 \registers_reg[26][14]  ( .D(n2884), .CK(n3891), .RN(n1058), .QN(
        n818) );
  DFFR_X1 \registers_reg[26][13]  ( .D(n2883), .CK(n3891), .RN(n1058), .QN(
        n819) );
  DFFR_X1 \registers_reg[26][12]  ( .D(n2882), .CK(n3891), .RN(n1058), .QN(
        n820) );
  DFFR_X1 \registers_reg[26][11]  ( .D(n2881), .CK(n3891), .RN(n1058), .QN(
        n821) );
  DFFR_X1 \registers_reg[26][10]  ( .D(n2880), .CK(n3891), .RN(n1058), .QN(
        n822) );
  DFFR_X1 \registers_reg[26][9]  ( .D(n2879), .CK(n3891), .RN(n1058), .QN(n823) );
  DFFR_X1 \registers_reg[26][8]  ( .D(n2878), .CK(n3891), .RN(n1058), .QN(n824) );
  DFFR_X1 \registers_reg[26][7]  ( .D(n2877), .CK(n3891), .RN(n1058), .QN(n825) );
  DFFR_X1 \registers_reg[26][6]  ( .D(n2876), .CK(n3891), .RN(n1058), .QN(n826) );
  DFFR_X1 \registers_reg[26][5]  ( .D(n2875), .CK(n3891), .RN(n1058), .QN(n827) );
  DFFR_X1 \registers_reg[26][4]  ( .D(n2874), .CK(n3891), .RN(n1057), .QN(n828) );
  DFFR_X1 \registers_reg[26][3]  ( .D(n2873), .CK(n3891), .RN(n1057), .QN(n829) );
  DFFR_X1 \registers_reg[26][2]  ( .D(n2872), .CK(n3891), .RN(n1057), .QN(n830) );
  DFFR_X1 \registers_reg[26][1]  ( .D(n2871), .CK(n3891), .RN(n1057), .QN(n831) );
  DFFR_X1 \registers_reg[26][0]  ( .D(n2870), .CK(n3891), .RN(n1057), .QN(n832) );
  DFFR_X1 \registers_reg[27][31]  ( .D(n2869), .CK(n3891), .RN(n1057), .QN(
        n833) );
  DFFR_X1 \registers_reg[27][30]  ( .D(n2868), .CK(n3891), .RN(n1057), .QN(
        n834) );
  DFFR_X1 \registers_reg[27][29]  ( .D(n2867), .CK(n3891), .RN(n1057), .QN(
        n835) );
  DFFR_X1 \registers_reg[27][28]  ( .D(n2866), .CK(n3891), .RN(n1057), .QN(
        n836) );
  DFFR_X1 \registers_reg[27][27]  ( .D(n2865), .CK(n3891), .RN(n1057), .QN(
        n837) );
  DFFR_X1 \registers_reg[27][26]  ( .D(n2864), .CK(n3891), .RN(n1057), .QN(
        n838) );
  DFFR_X1 \registers_reg[27][25]  ( .D(n2863), .CK(n3891), .RN(n1056), .QN(
        n839) );
  DFFR_X1 \registers_reg[27][24]  ( .D(n2862), .CK(n3891), .RN(n1056), .QN(
        n840) );
  DFFR_X1 \registers_reg[27][23]  ( .D(n2861), .CK(n3891), .RN(n1056), .QN(
        n841) );
  DFFR_X1 \registers_reg[27][22]  ( .D(n2860), .CK(n3891), .RN(n1056), .QN(
        n842) );
  DFFR_X1 \registers_reg[27][21]  ( .D(n2859), .CK(n3891), .RN(n1056), .QN(
        n843) );
  DFFR_X1 \registers_reg[27][20]  ( .D(n2858), .CK(n3891), .RN(n1056), .QN(
        n844) );
  DFFR_X1 \registers_reg[27][19]  ( .D(n2857), .CK(n3891), .RN(n1056), .QN(
        n845) );
  DFFR_X1 \registers_reg[27][18]  ( .D(n2856), .CK(n3891), .RN(n1056), .QN(
        n846) );
  DFFR_X1 \registers_reg[27][17]  ( .D(n2855), .CK(n3891), .RN(n1056), .QN(
        n847) );
  DFFR_X1 \registers_reg[27][16]  ( .D(n2854), .CK(n3891), .RN(n1056), .QN(
        n848) );
  DFFR_X1 \registers_reg[27][15]  ( .D(n2853), .CK(n3891), .RN(n1056), .QN(
        n849) );
  DFFR_X1 \registers_reg[27][14]  ( .D(n2852), .CK(n3891), .RN(n1055), .QN(
        n850) );
  DFFR_X1 \registers_reg[27][13]  ( .D(n2851), .CK(n3891), .RN(n1055), .QN(
        n851) );
  DFFR_X1 \registers_reg[27][12]  ( .D(n2850), .CK(n3891), .RN(n1055), .QN(
        n852) );
  DFFR_X1 \registers_reg[27][11]  ( .D(n2849), .CK(n3891), .RN(n1055), .QN(
        n853) );
  DFFR_X1 \registers_reg[27][10]  ( .D(n2848), .CK(n3891), .RN(n1055), .QN(
        n854) );
  DFFR_X1 \registers_reg[27][9]  ( .D(n2847), .CK(n3891), .RN(n1055), .QN(n855) );
  DFFR_X1 \registers_reg[27][8]  ( .D(n2846), .CK(n3891), .RN(n1055), .QN(n856) );
  DFFR_X1 \registers_reg[27][7]  ( .D(n2845), .CK(n3891), .RN(n1055), .QN(n857) );
  DFFR_X1 \registers_reg[27][6]  ( .D(n2844), .CK(n3891), .RN(n1055), .QN(n858) );
  DFFR_X1 \registers_reg[27][5]  ( .D(n2843), .CK(n3891), .RN(n1055), .QN(n859) );
  DFFR_X1 \registers_reg[27][4]  ( .D(n2842), .CK(n3891), .RN(n1055), .QN(n860) );
  DFFR_X1 \registers_reg[27][3]  ( .D(n2841), .CK(n3891), .RN(n1054), .QN(n861) );
  DFFR_X1 \registers_reg[27][2]  ( .D(n2840), .CK(n3891), .RN(n1054), .QN(n862) );
  DFFR_X1 \registers_reg[27][1]  ( .D(n2839), .CK(n3891), .RN(n1054), .QN(n863) );
  DFFR_X1 \registers_reg[27][0]  ( .D(n2838), .CK(n3891), .RN(n1054), .QN(n864) );
  DFFR_X1 \registers_reg[28][31]  ( .D(n3816), .CK(n3891), .RN(n1054), .Q(
        \registers[28][31] ) );
  DFFR_X1 \registers_reg[28][30]  ( .D(n3815), .CK(n3891), .RN(n1054), .Q(
        \registers[28][30] ) );
  DFFR_X1 \registers_reg[28][29]  ( .D(n3814), .CK(n3891), .RN(n1054), .Q(
        \registers[28][29] ) );
  DFFR_X1 \registers_reg[28][28]  ( .D(n3813), .CK(n3891), .RN(n1054), .Q(
        \registers[28][28] ) );
  DFFR_X1 \registers_reg[28][27]  ( .D(n3812), .CK(n3891), .RN(n1054), .Q(
        \registers[28][27] ) );
  DFFR_X1 \registers_reg[28][26]  ( .D(n3811), .CK(n3891), .RN(n1054), .Q(
        \registers[28][26] ) );
  DFFR_X1 \registers_reg[28][25]  ( .D(n3810), .CK(n3891), .RN(n1054), .Q(
        \registers[28][25] ) );
  DFFR_X1 \registers_reg[28][24]  ( .D(n3809), .CK(n3891), .RN(n1053), .Q(
        \registers[28][24] ) );
  DFFR_X1 \registers_reg[28][23]  ( .D(n3808), .CK(n3891), .RN(n1053), .Q(
        \registers[28][23] ) );
  DFFR_X1 \registers_reg[28][22]  ( .D(n3807), .CK(n3891), .RN(n1053), .Q(
        \registers[28][22] ) );
  DFFR_X1 \registers_reg[28][21]  ( .D(n3806), .CK(n3891), .RN(n1053), .Q(
        \registers[28][21] ) );
  DFFR_X1 \registers_reg[28][20]  ( .D(n3805), .CK(n3891), .RN(n1053), .Q(
        \registers[28][20] ) );
  DFFR_X1 \registers_reg[28][19]  ( .D(n3804), .CK(n3891), .RN(n1053), .Q(
        \registers[28][19] ) );
  DFFR_X1 \registers_reg[28][18]  ( .D(n3803), .CK(n3891), .RN(n1053), .Q(
        \registers[28][18] ) );
  DFFR_X1 \registers_reg[28][17]  ( .D(n3802), .CK(n3891), .RN(n1053), .Q(
        \registers[28][17] ) );
  DFFR_X1 \registers_reg[28][16]  ( .D(n3801), .CK(n3891), .RN(n1053), .Q(
        \registers[28][16] ) );
  DFFR_X1 \registers_reg[28][15]  ( .D(n3800), .CK(n3891), .RN(n1053), .Q(
        \registers[28][15] ) );
  DFFR_X1 \registers_reg[28][14]  ( .D(n3799), .CK(n3891), .RN(n1053), .Q(
        \registers[28][14] ) );
  DFFR_X1 \registers_reg[28][13]  ( .D(n3798), .CK(n3891), .RN(n1052), .Q(
        \registers[28][13] ) );
  DFFR_X1 \registers_reg[28][12]  ( .D(n3797), .CK(n3891), .RN(n1052), .Q(
        \registers[28][12] ) );
  DFFR_X1 \registers_reg[28][11]  ( .D(n3796), .CK(n3891), .RN(n1052), .Q(
        \registers[28][11] ) );
  DFFR_X1 \registers_reg[28][10]  ( .D(n3795), .CK(n3891), .RN(n1052), .Q(
        \registers[28][10] ) );
  DFFR_X1 \registers_reg[28][9]  ( .D(n3794), .CK(n3891), .RN(n1052), .Q(
        \registers[28][9] ) );
  DFFR_X1 \registers_reg[28][8]  ( .D(n3793), .CK(n3891), .RN(n1052), .Q(
        \registers[28][8] ) );
  DFFR_X1 \registers_reg[28][7]  ( .D(n3792), .CK(n3891), .RN(n1052), .Q(
        \registers[28][7] ) );
  DFFR_X1 \registers_reg[28][6]  ( .D(n3791), .CK(n3891), .RN(n1052), .Q(
        \registers[28][6] ) );
  DFFR_X1 \registers_reg[28][5]  ( .D(n3790), .CK(n3891), .RN(n1052), .Q(
        \registers[28][5] ) );
  DFFR_X1 \registers_reg[28][4]  ( .D(n3789), .CK(n3891), .RN(n1052), .Q(
        \registers[28][4] ) );
  DFFR_X1 \registers_reg[28][3]  ( .D(n3788), .CK(n3891), .RN(n1052), .Q(
        \registers[28][3] ) );
  DFFR_X1 \registers_reg[28][2]  ( .D(n3787), .CK(n3891), .RN(n1051), .Q(
        \registers[28][2] ) );
  DFFR_X1 \registers_reg[28][1]  ( .D(n3786), .CK(n3891), .RN(n1051), .Q(
        \registers[28][1] ) );
  DFFR_X1 \registers_reg[28][0]  ( .D(n3785), .CK(n3891), .RN(n1051), .Q(
        \registers[28][0] ) );
  DFFR_X1 \registers_reg[29][31]  ( .D(n3848), .CK(n3891), .RN(n1051), .Q(
        \registers[29][31] ) );
  DFFR_X1 \registers_reg[29][30]  ( .D(n3847), .CK(n3891), .RN(n1051), .Q(
        \registers[29][30] ) );
  DFFR_X1 \registers_reg[29][29]  ( .D(n3846), .CK(n3891), .RN(n1051), .Q(
        \registers[29][29] ) );
  DFFR_X1 \registers_reg[29][28]  ( .D(n3845), .CK(n3891), .RN(n1051), .Q(
        \registers[29][28] ) );
  DFFR_X1 \registers_reg[29][27]  ( .D(n3844), .CK(n3891), .RN(n1051), .Q(
        \registers[29][27] ) );
  DFFR_X1 \registers_reg[29][26]  ( .D(n3843), .CK(n3891), .RN(n1051), .Q(
        \registers[29][26] ) );
  DFFR_X1 \registers_reg[29][25]  ( .D(n3842), .CK(n3891), .RN(n1051), .Q(
        \registers[29][25] ) );
  DFFR_X1 \registers_reg[29][24]  ( .D(n3841), .CK(n3891), .RN(n1051), .Q(
        \registers[29][24] ) );
  DFFR_X1 \registers_reg[29][23]  ( .D(n3840), .CK(n3891), .RN(n1050), .Q(
        \registers[29][23] ) );
  DFFR_X1 \registers_reg[29][22]  ( .D(n3839), .CK(n3891), .RN(n1050), .Q(
        \registers[29][22] ) );
  DFFR_X1 \registers_reg[29][21]  ( .D(n3838), .CK(n3891), .RN(n1050), .Q(
        \registers[29][21] ) );
  DFFR_X1 \registers_reg[29][20]  ( .D(n3837), .CK(n3891), .RN(n1050), .Q(
        \registers[29][20] ) );
  DFFR_X1 \registers_reg[29][19]  ( .D(n3836), .CK(n3891), .RN(n1050), .Q(
        \registers[29][19] ) );
  DFFR_X1 \registers_reg[29][18]  ( .D(n3835), .CK(n3891), .RN(n1050), .Q(
        \registers[29][18] ) );
  DFFR_X1 \registers_reg[29][17]  ( .D(n3834), .CK(n3891), .RN(n1050), .Q(
        \registers[29][17] ) );
  DFFR_X1 \registers_reg[29][16]  ( .D(n3833), .CK(n3891), .RN(n1050), .Q(
        \registers[29][16] ) );
  DFFR_X1 \registers_reg[29][15]  ( .D(n3832), .CK(n3891), .RN(n1050), .Q(
        \registers[29][15] ) );
  DFFR_X1 \registers_reg[29][14]  ( .D(n3831), .CK(n3891), .RN(n1050), .Q(
        \registers[29][14] ) );
  DFFR_X1 \registers_reg[29][13]  ( .D(n3830), .CK(n3891), .RN(n1050), .Q(
        \registers[29][13] ) );
  DFFR_X1 \registers_reg[29][12]  ( .D(n3829), .CK(n3891), .RN(n1049), .Q(
        \registers[29][12] ) );
  DFFR_X1 \registers_reg[29][11]  ( .D(n3828), .CK(n3891), .RN(n1049), .Q(
        \registers[29][11] ) );
  DFFR_X1 \registers_reg[29][10]  ( .D(n3827), .CK(n3891), .RN(n1049), .Q(
        \registers[29][10] ) );
  DFFR_X1 \registers_reg[29][9]  ( .D(n3826), .CK(n3891), .RN(n1049), .Q(
        \registers[29][9] ) );
  DFFR_X1 \registers_reg[29][8]  ( .D(n3825), .CK(n3891), .RN(n1049), .Q(
        \registers[29][8] ) );
  DFFR_X1 \registers_reg[29][7]  ( .D(n3824), .CK(n3891), .RN(n1049), .Q(
        \registers[29][7] ) );
  DFFR_X1 \registers_reg[29][6]  ( .D(n3823), .CK(n3891), .RN(n1049), .Q(
        \registers[29][6] ) );
  DFFR_X1 \registers_reg[29][5]  ( .D(n3822), .CK(n3891), .RN(n1049), .Q(
        \registers[29][5] ) );
  DFFR_X1 \registers_reg[29][4]  ( .D(n3821), .CK(n3891), .RN(n1049), .Q(
        \registers[29][4] ) );
  DFFR_X1 \registers_reg[29][3]  ( .D(n3820), .CK(n3891), .RN(n1049), .Q(
        \registers[29][3] ) );
  DFFR_X1 \registers_reg[29][2]  ( .D(n3819), .CK(n3891), .RN(n1049), .Q(
        \registers[29][2] ) );
  DFFR_X1 \registers_reg[29][1]  ( .D(n3818), .CK(n3891), .RN(n1048), .Q(
        \registers[29][1] ) );
  DFFR_X1 \registers_reg[29][0]  ( .D(n3817), .CK(n3891), .RN(n1048), .Q(
        \registers[29][0] ) );
  DFFR_X1 \registers_reg[30][31]  ( .D(n2837), .CK(n3891), .RN(n1048), .QN(
        n929) );
  DFFR_X1 \registers_reg[30][30]  ( .D(n2836), .CK(n3891), .RN(n1048), .QN(
        n930) );
  DFFR_X1 \registers_reg[30][29]  ( .D(n2835), .CK(n3891), .RN(n1048), .QN(
        n931) );
  DFFR_X1 \registers_reg[30][28]  ( .D(n2834), .CK(n3891), .RN(n1048), .QN(
        n932) );
  DFFR_X1 \registers_reg[30][27]  ( .D(n2833), .CK(n3891), .RN(n1048), .QN(
        n933) );
  DFFR_X1 \registers_reg[30][26]  ( .D(n2832), .CK(n3891), .RN(n1048), .QN(
        n934) );
  DFFR_X1 \registers_reg[30][25]  ( .D(n2831), .CK(n3891), .RN(n1048), .QN(
        n935) );
  DFFR_X1 \registers_reg[30][24]  ( .D(n2830), .CK(n3891), .RN(n1048), .QN(
        n936) );
  DFFR_X1 \registers_reg[30][23]  ( .D(n2829), .CK(n3891), .RN(n1048), .QN(
        n937) );
  DFFR_X1 \registers_reg[30][22]  ( .D(n2828), .CK(n3891), .RN(n1047), .QN(
        n938) );
  DFFR_X1 \registers_reg[30][21]  ( .D(n2827), .CK(n3891), .RN(n1047), .QN(
        n939) );
  DFFR_X1 \registers_reg[30][20]  ( .D(n2826), .CK(n3891), .RN(n1047), .QN(
        n940) );
  DFFR_X1 \registers_reg[30][19]  ( .D(n2825), .CK(n3891), .RN(n1047), .QN(
        n941) );
  DFFR_X1 \registers_reg[30][18]  ( .D(n2824), .CK(n3891), .RN(n1047), .QN(
        n942) );
  DFFR_X1 \registers_reg[30][17]  ( .D(n2823), .CK(n3891), .RN(n1047), .QN(
        n943) );
  DFFR_X1 \registers_reg[30][16]  ( .D(n2822), .CK(n3891), .RN(n1047), .QN(
        n944) );
  DFFR_X1 \registers_reg[30][15]  ( .D(n2821), .CK(n3891), .RN(n1047), .QN(
        n945) );
  DFFR_X1 \registers_reg[30][14]  ( .D(n2820), .CK(n3891), .RN(n1047), .QN(
        n946) );
  DFFR_X1 \registers_reg[30][13]  ( .D(n2819), .CK(n3891), .RN(n1047), .QN(
        n947) );
  DFFR_X1 \registers_reg[30][12]  ( .D(n2818), .CK(n3891), .RN(n1047), .QN(
        n948) );
  DFFR_X1 \registers_reg[30][11]  ( .D(n2817), .CK(n3891), .RN(n1046), .QN(
        n949) );
  DFFR_X1 \registers_reg[30][10]  ( .D(n2816), .CK(n3891), .RN(n1046), .QN(
        n950) );
  DFFR_X1 \registers_reg[30][9]  ( .D(n2815), .CK(n3891), .RN(n1046), .QN(n951) );
  DFFR_X1 \registers_reg[30][8]  ( .D(n2814), .CK(n3891), .RN(n1046), .QN(n952) );
  DFFR_X1 \registers_reg[30][7]  ( .D(n2813), .CK(n3891), .RN(n1046), .QN(n953) );
  DFFR_X1 \registers_reg[30][6]  ( .D(n2812), .CK(n3891), .RN(n1046), .QN(n954) );
  DFFR_X1 \registers_reg[30][5]  ( .D(n2811), .CK(n3891), .RN(n1046), .QN(n955) );
  DFFR_X1 \registers_reg[30][4]  ( .D(n2810), .CK(n3891), .RN(n1046), .QN(n956) );
  DFFR_X1 \registers_reg[30][3]  ( .D(n2809), .CK(n3891), .RN(n1046), .QN(n957) );
  DFFR_X1 \registers_reg[30][2]  ( .D(n2808), .CK(n3891), .RN(n1046), .QN(n958) );
  DFFR_X1 \registers_reg[30][1]  ( .D(n2807), .CK(n3891), .RN(n1046), .QN(n959) );
  DFFR_X1 \registers_reg[30][0]  ( .D(n2806), .CK(n3891), .RN(n1045), .QN(n960) );
  DFFR_X1 \registers_reg[31][31]  ( .D(n2805), .CK(n3891), .RN(n1045), .QN(
        n961) );
  DFFR_X1 \registers_reg[31][30]  ( .D(n2804), .CK(n3891), .RN(n1045), .QN(
        n962) );
  DFFR_X1 \registers_reg[31][29]  ( .D(n2803), .CK(n3891), .RN(n1045), .QN(
        n963) );
  DFFR_X1 \registers_reg[31][28]  ( .D(n2802), .CK(n3891), .RN(n1045), .QN(
        n964) );
  DFFR_X1 \registers_reg[31][27]  ( .D(n2801), .CK(n3891), .RN(n1045), .QN(
        n965) );
  DFFR_X1 \registers_reg[31][26]  ( .D(n2800), .CK(n3891), .RN(n1045), .QN(
        n966) );
  DFFR_X1 \registers_reg[31][25]  ( .D(n2799), .CK(n3891), .RN(n1045), .QN(
        n967) );
  DFFR_X1 \registers_reg[31][24]  ( .D(n2798), .CK(n3891), .RN(n1045), .QN(
        n968) );
  DFFR_X1 \registers_reg[31][23]  ( .D(n2797), .CK(n3891), .RN(n1045), .QN(
        n969) );
  DFFR_X1 \registers_reg[31][22]  ( .D(n2796), .CK(n3891), .RN(n1045), .QN(
        n970) );
  DFFR_X1 \registers_reg[31][21]  ( .D(n2795), .CK(n3891), .RN(n1044), .QN(
        n971) );
  DFFR_X1 \registers_reg[31][20]  ( .D(n2794), .CK(n3891), .RN(n1044), .QN(
        n972) );
  DFFR_X1 \registers_reg[31][19]  ( .D(n2793), .CK(n3891), .RN(n1044), .QN(
        n973) );
  DFFR_X1 \registers_reg[31][18]  ( .D(n2792), .CK(n3891), .RN(n1044), .QN(
        n974) );
  DFFR_X1 \registers_reg[31][17]  ( .D(n2791), .CK(n3891), .RN(n1044), .QN(
        n975) );
  DFFR_X1 \registers_reg[31][16]  ( .D(n2790), .CK(n3891), .RN(n1044), .QN(
        n976) );
  DFFR_X1 \registers_reg[31][15]  ( .D(n2789), .CK(n3891), .RN(n1044), .QN(
        n977) );
  DFFR_X1 \registers_reg[31][14]  ( .D(n2788), .CK(n3891), .RN(n1044), .QN(
        n978) );
  DFFR_X1 \registers_reg[31][13]  ( .D(n2787), .CK(n3891), .RN(n1044), .QN(
        n979) );
  DFFR_X1 \registers_reg[31][12]  ( .D(n2786), .CK(n3891), .RN(n1044), .QN(
        n980) );
  DFFR_X1 \registers_reg[31][11]  ( .D(n2785), .CK(n3891), .RN(n1044), .QN(
        n981) );
  DFFR_X1 \registers_reg[31][10]  ( .D(n2784), .CK(n3891), .RN(n1043), .QN(
        n982) );
  DFFR_X1 \registers_reg[31][9]  ( .D(n2783), .CK(n3891), .RN(n1043), .QN(n983) );
  DFFR_X1 \registers_reg[31][8]  ( .D(n2782), .CK(n3891), .RN(n1043), .QN(n984) );
  DFFR_X1 \registers_reg[31][7]  ( .D(n2781), .CK(n3891), .RN(n1043), .QN(n985) );
  DFFR_X1 \registers_reg[31][6]  ( .D(n2780), .CK(n3891), .RN(n1043), .QN(n986) );
  DFFR_X1 \registers_reg[31][5]  ( .D(n2779), .CK(n3891), .RN(n1043), .QN(n987) );
  DFFR_X1 \registers_reg[31][4]  ( .D(n2778), .CK(n3891), .RN(n1043), .QN(n988) );
  DFFR_X1 \registers_reg[31][3]  ( .D(n2777), .CK(n3891), .RN(n1043), .QN(n989) );
  DFFR_X1 \registers_reg[31][2]  ( .D(n2776), .CK(n3891), .RN(n1043), .QN(n990) );
  DFFR_X1 \registers_reg[31][1]  ( .D(n2775), .CK(n3891), .RN(n1043), .QN(n991) );
  DFFR_X1 \registers_reg[31][0]  ( .D(n2774), .CK(n3891), .RN(n1043), .QN(n992) );
  DLH_X1 \OUT1_reg[31]  ( .G(n1028), .D(N217), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n1028), .D(N216), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n1028), .D(N215), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n1028), .D(N214), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n1028), .D(N213), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n1028), .D(N212), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n1028), .D(N211), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n1028), .D(N210), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n1028), .D(N209), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n1028), .D(N208), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n1029), .D(N207), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n1029), .D(N206), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n1029), .D(N205), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n1029), .D(N204), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n1029), .D(N203), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n1029), .D(N202), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n1029), .D(N201), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n1029), .D(N200), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n1029), .D(N199), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n1029), .D(N198), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n1030), .D(N197), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n1030), .D(N196), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n1030), .D(N195), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n1030), .D(N194), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n1030), .D(N193), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n1030), .D(N192), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n1030), .D(N191), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n1030), .D(N190), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n1030), .D(N189), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n1030), .D(N188), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n1031), .D(N187), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n1031), .D(N186), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(n1024), .D(N352), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n1024), .D(N351), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n1024), .D(N350), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n1024), .D(N349), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n1024), .D(N348), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n1024), .D(N347), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n1024), .D(N346), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n1024), .D(N345), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n1024), .D(N344), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n1024), .D(N343), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n1025), .D(N342), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n1025), .D(N341), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n1025), .D(N340), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n1025), .D(N339), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n1025), .D(N338), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n1025), .D(N337), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n1025), .D(N336), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n1025), .D(N335), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n1025), .D(N334), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n1025), .D(N333), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n1026), .D(N332), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n1026), .D(N331), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n1026), .D(N330), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n1026), .D(N329), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n1026), .D(N328), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n1026), .D(N327), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n1026), .D(N326), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n1026), .D(N325), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n1026), .D(N324), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n1026), .D(N323), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n1027), .D(N322), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n1027), .D(N321), .Q(OUT2[0]) );
  OAI22_X2 U2 ( .A1(n1017), .A2(n3890), .B1(n1016), .B2(n992), .ZN(n2774) );
  OAI22_X2 U3 ( .A1(n1017), .A2(n3889), .B1(n1016), .B2(n991), .ZN(n2775) );
  OAI22_X2 U4 ( .A1(n1017), .A2(n3888), .B1(n1016), .B2(n990), .ZN(n2776) );
  OAI22_X2 U5 ( .A1(n1017), .A2(n3887), .B1(n1016), .B2(n989), .ZN(n2777) );
  OAI22_X2 U6 ( .A1(n1017), .A2(n3886), .B1(n1016), .B2(n988), .ZN(n2778) );
  OAI22_X2 U7 ( .A1(n1018), .A2(n3885), .B1(n1016), .B2(n987), .ZN(n2779) );
  OAI22_X2 U8 ( .A1(n1018), .A2(n3884), .B1(n1016), .B2(n986), .ZN(n2780) );
  OAI22_X2 U9 ( .A1(n1018), .A2(n3883), .B1(n1016), .B2(n985), .ZN(n2781) );
  OAI22_X2 U10 ( .A1(n1018), .A2(n3882), .B1(n1016), .B2(n984), .ZN(n2782) );
  OAI22_X2 U11 ( .A1(n1018), .A2(n3881), .B1(n1016), .B2(n983), .ZN(n2783) );
  OAI22_X2 U12 ( .A1(n1019), .A2(n3880), .B1(n1015), .B2(n982), .ZN(n2784) );
  OAI22_X2 U13 ( .A1(n1019), .A2(n3879), .B1(n1015), .B2(n981), .ZN(n2785) );
  OAI22_X2 U14 ( .A1(n1019), .A2(n3878), .B1(n1015), .B2(n980), .ZN(n2786) );
  OAI22_X2 U15 ( .A1(n1019), .A2(n3877), .B1(n1015), .B2(n979), .ZN(n2787) );
  OAI22_X2 U16 ( .A1(n1019), .A2(n3876), .B1(n1015), .B2(n978), .ZN(n2788) );
  OAI22_X2 U17 ( .A1(n1020), .A2(n3875), .B1(n1015), .B2(n977), .ZN(n2789) );
  OAI22_X2 U18 ( .A1(n1020), .A2(n3874), .B1(n1015), .B2(n976), .ZN(n2790) );
  OAI22_X2 U19 ( .A1(n1020), .A2(n3873), .B1(n1015), .B2(n975), .ZN(n2791) );
  OAI22_X2 U20 ( .A1(n1020), .A2(n3872), .B1(n1015), .B2(n974), .ZN(n2792) );
  OAI22_X2 U21 ( .A1(n1020), .A2(n3871), .B1(n1015), .B2(n973), .ZN(n2793) );
  OAI22_X2 U22 ( .A1(n1021), .A2(n3870), .B1(n1015), .B2(n972), .ZN(n2794) );
  OAI22_X2 U23 ( .A1(n1021), .A2(n3869), .B1(n1014), .B2(n971), .ZN(n2795) );
  OAI22_X2 U24 ( .A1(n1021), .A2(n3868), .B1(n1014), .B2(n970), .ZN(n2796) );
  OAI22_X2 U25 ( .A1(n1021), .A2(n3867), .B1(n1014), .B2(n969), .ZN(n2797) );
  OAI22_X2 U26 ( .A1(n1021), .A2(n3866), .B1(n1014), .B2(n968), .ZN(n2798) );
  OAI22_X2 U27 ( .A1(n1022), .A2(n3865), .B1(n1014), .B2(n967), .ZN(n2799) );
  OAI22_X2 U28 ( .A1(n1022), .A2(n3864), .B1(n1014), .B2(n966), .ZN(n2800) );
  OAI22_X2 U29 ( .A1(n1022), .A2(n3863), .B1(n1014), .B2(n965), .ZN(n2801) );
  OAI22_X2 U30 ( .A1(n1022), .A2(n3862), .B1(n1014), .B2(n964), .ZN(n2802) );
  OAI22_X2 U31 ( .A1(n1022), .A2(n3861), .B1(n1014), .B2(n963), .ZN(n2803) );
  OAI22_X2 U32 ( .A1(n1023), .A2(n3860), .B1(n1014), .B2(n962), .ZN(n2804) );
  OAI22_X2 U33 ( .A1(n1023), .A2(n3859), .B1(n1014), .B2(n961), .ZN(n2805) );
  NAND2_X2 U34 ( .A1(n1069), .A2(n1070), .ZN(n1068) );
  OAI22_X2 U35 ( .A1(n3890), .A2(n1005), .B1(n1006), .B2(n960), .ZN(n2806) );
  OAI22_X2 U36 ( .A1(n3889), .A2(n1005), .B1(n1006), .B2(n959), .ZN(n2807) );
  OAI22_X2 U37 ( .A1(n3888), .A2(n1005), .B1(n1006), .B2(n958), .ZN(n2808) );
  OAI22_X2 U38 ( .A1(n3887), .A2(n1005), .B1(n1006), .B2(n957), .ZN(n2809) );
  OAI22_X2 U39 ( .A1(n3886), .A2(n1005), .B1(n1006), .B2(n956), .ZN(n2810) );
  OAI22_X2 U40 ( .A1(n3885), .A2(n1005), .B1(n1007), .B2(n955), .ZN(n2811) );
  OAI22_X2 U41 ( .A1(n3884), .A2(n1005), .B1(n1007), .B2(n954), .ZN(n2812) );
  OAI22_X2 U42 ( .A1(n3883), .A2(n1005), .B1(n1007), .B2(n953), .ZN(n2813) );
  OAI22_X2 U43 ( .A1(n3882), .A2(n1004), .B1(n1007), .B2(n952), .ZN(n2814) );
  OAI22_X2 U44 ( .A1(n3881), .A2(n1004), .B1(n1007), .B2(n951), .ZN(n2815) );
  OAI22_X2 U45 ( .A1(n3880), .A2(n1004), .B1(n1008), .B2(n950), .ZN(n2816) );
  OAI22_X2 U46 ( .A1(n3879), .A2(n1004), .B1(n1008), .B2(n949), .ZN(n2817) );
  OAI22_X2 U47 ( .A1(n3878), .A2(n1004), .B1(n1008), .B2(n948), .ZN(n2818) );
  OAI22_X2 U48 ( .A1(n3877), .A2(n1004), .B1(n1008), .B2(n947), .ZN(n2819) );
  OAI22_X2 U49 ( .A1(n3876), .A2(n1004), .B1(n1008), .B2(n946), .ZN(n2820) );
  OAI22_X2 U50 ( .A1(n3875), .A2(n1004), .B1(n1009), .B2(n945), .ZN(n2821) );
  OAI22_X2 U51 ( .A1(n3874), .A2(n1004), .B1(n1009), .B2(n944), .ZN(n2822) );
  OAI22_X2 U52 ( .A1(n3873), .A2(n1004), .B1(n1009), .B2(n943), .ZN(n2823) );
  OAI22_X2 U53 ( .A1(n3872), .A2(n1004), .B1(n1009), .B2(n942), .ZN(n2824) );
  OAI22_X2 U54 ( .A1(n3871), .A2(n1004), .B1(n1009), .B2(n941), .ZN(n2825) );
  OAI22_X2 U55 ( .A1(n3870), .A2(n1003), .B1(n1010), .B2(n940), .ZN(n2826) );
  OAI22_X2 U56 ( .A1(n3869), .A2(n1003), .B1(n1010), .B2(n939), .ZN(n2827) );
  OAI22_X2 U57 ( .A1(n3868), .A2(n1003), .B1(n1010), .B2(n938), .ZN(n2828) );
  OAI22_X2 U58 ( .A1(n3867), .A2(n1003), .B1(n1010), .B2(n937), .ZN(n2829) );
  OAI22_X2 U59 ( .A1(n3866), .A2(n1003), .B1(n1010), .B2(n936), .ZN(n2830) );
  OAI22_X2 U60 ( .A1(n3865), .A2(n1003), .B1(n1011), .B2(n935), .ZN(n2831) );
  OAI22_X2 U61 ( .A1(n3864), .A2(n1003), .B1(n1011), .B2(n934), .ZN(n2832) );
  OAI22_X2 U62 ( .A1(n3863), .A2(n1003), .B1(n1011), .B2(n933), .ZN(n2833) );
  OAI22_X2 U63 ( .A1(n3862), .A2(n1003), .B1(n1011), .B2(n932), .ZN(n2834) );
  OAI22_X2 U64 ( .A1(n3861), .A2(n1003), .B1(n1011), .B2(n931), .ZN(n2835) );
  OAI22_X2 U65 ( .A1(n3860), .A2(n1003), .B1(n1012), .B2(n930), .ZN(n2836) );
  OAI22_X2 U66 ( .A1(n3859), .A2(n1003), .B1(n1012), .B2(n929), .ZN(n2837) );
  NAND2_X2 U67 ( .A1(n1072), .A2(n1070), .ZN(n1071) );
  AOI22_X2 U68 ( .A1(DATAIN[0]), .A2(n995), .B1(n996), .B2(\registers[29][0] ), 
        .ZN(n1073) );
  AOI22_X2 U69 ( .A1(DATAIN[1]), .A2(n995), .B1(n996), .B2(\registers[29][1] ), 
        .ZN(n1075) );
  AOI22_X2 U70 ( .A1(DATAIN[2]), .A2(n995), .B1(n996), .B2(\registers[29][2] ), 
        .ZN(n1076) );
  AOI22_X2 U71 ( .A1(DATAIN[3]), .A2(n995), .B1(n996), .B2(\registers[29][3] ), 
        .ZN(n1077) );
  AOI22_X2 U72 ( .A1(DATAIN[4]), .A2(n995), .B1(n996), .B2(\registers[29][4] ), 
        .ZN(n1078) );
  AOI22_X2 U73 ( .A1(DATAIN[5]), .A2(n995), .B1(n997), .B2(\registers[29][5] ), 
        .ZN(n1079) );
  AOI22_X2 U74 ( .A1(DATAIN[6]), .A2(n995), .B1(n997), .B2(\registers[29][6] ), 
        .ZN(n1080) );
  AOI22_X2 U75 ( .A1(DATAIN[7]), .A2(n995), .B1(n997), .B2(\registers[29][7] ), 
        .ZN(n1081) );
  AOI22_X2 U76 ( .A1(DATAIN[8]), .A2(n994), .B1(n997), .B2(\registers[29][8] ), 
        .ZN(n1082) );
  AOI22_X2 U77 ( .A1(DATAIN[9]), .A2(n994), .B1(n997), .B2(\registers[29][9] ), 
        .ZN(n1083) );
  AOI22_X2 U78 ( .A1(DATAIN[10]), .A2(n994), .B1(n998), .B2(
        \registers[29][10] ), .ZN(n1084) );
  AOI22_X2 U79 ( .A1(DATAIN[11]), .A2(n994), .B1(n998), .B2(
        \registers[29][11] ), .ZN(n1085) );
  AOI22_X2 U80 ( .A1(DATAIN[12]), .A2(n994), .B1(n998), .B2(
        \registers[29][12] ), .ZN(n1086) );
  AOI22_X2 U81 ( .A1(DATAIN[13]), .A2(n994), .B1(n998), .B2(
        \registers[29][13] ), .ZN(n1087) );
  AOI22_X2 U82 ( .A1(DATAIN[14]), .A2(n994), .B1(n998), .B2(
        \registers[29][14] ), .ZN(n1088) );
  AOI22_X2 U83 ( .A1(DATAIN[15]), .A2(n994), .B1(n999), .B2(
        \registers[29][15] ), .ZN(n1089) );
  AOI22_X2 U84 ( .A1(DATAIN[16]), .A2(n994), .B1(n999), .B2(
        \registers[29][16] ), .ZN(n1090) );
  AOI22_X2 U85 ( .A1(DATAIN[17]), .A2(n994), .B1(n999), .B2(
        \registers[29][17] ), .ZN(n1091) );
  AOI22_X2 U86 ( .A1(DATAIN[18]), .A2(n994), .B1(n999), .B2(
        \registers[29][18] ), .ZN(n1092) );
  AOI22_X2 U87 ( .A1(DATAIN[19]), .A2(n994), .B1(n999), .B2(
        \registers[29][19] ), .ZN(n1093) );
  AOI22_X2 U88 ( .A1(DATAIN[20]), .A2(n993), .B1(n1000), .B2(
        \registers[29][20] ), .ZN(n1094) );
  AOI22_X2 U89 ( .A1(DATAIN[21]), .A2(n993), .B1(n1000), .B2(
        \registers[29][21] ), .ZN(n1095) );
  AOI22_X2 U90 ( .A1(DATAIN[22]), .A2(n993), .B1(n1000), .B2(
        \registers[29][22] ), .ZN(n1096) );
  AOI22_X2 U91 ( .A1(DATAIN[23]), .A2(n993), .B1(n1000), .B2(
        \registers[29][23] ), .ZN(n1097) );
  AOI22_X2 U92 ( .A1(DATAIN[24]), .A2(n993), .B1(n1000), .B2(
        \registers[29][24] ), .ZN(n1098) );
  AOI22_X2 U93 ( .A1(DATAIN[25]), .A2(n993), .B1(n1001), .B2(
        \registers[29][25] ), .ZN(n1099) );
  AOI22_X2 U94 ( .A1(DATAIN[26]), .A2(n993), .B1(n1001), .B2(
        \registers[29][26] ), .ZN(n1100) );
  AOI22_X2 U95 ( .A1(DATAIN[27]), .A2(n993), .B1(n1001), .B2(
        \registers[29][27] ), .ZN(n1101) );
  AOI22_X2 U96 ( .A1(DATAIN[28]), .A2(n993), .B1(n1001), .B2(
        \registers[29][28] ), .ZN(n1102) );
  AOI22_X2 U97 ( .A1(DATAIN[29]), .A2(n993), .B1(n1001), .B2(
        \registers[29][29] ), .ZN(n1103) );
  AOI22_X2 U98 ( .A1(DATAIN[30]), .A2(n993), .B1(n1002), .B2(
        \registers[29][30] ), .ZN(n1104) );
  AOI22_X2 U99 ( .A1(DATAIN[31]), .A2(n993), .B1(n1002), .B2(
        \registers[29][31] ), .ZN(n1105) );
  NAND2_X2 U100 ( .A1(n1106), .A2(n1070), .ZN(n1074) );
  AOI22_X2 U101 ( .A1(DATAIN[0]), .A2(n921), .B1(n922), .B2(\registers[28][0] ), .ZN(n1107) );
  AOI22_X2 U102 ( .A1(DATAIN[1]), .A2(n921), .B1(n922), .B2(\registers[28][1] ), .ZN(n1109) );
  AOI22_X2 U103 ( .A1(DATAIN[2]), .A2(n921), .B1(n922), .B2(\registers[28][2] ), .ZN(n1110) );
  AOI22_X2 U104 ( .A1(DATAIN[3]), .A2(n921), .B1(n922), .B2(\registers[28][3] ), .ZN(n1111) );
  AOI22_X2 U105 ( .A1(DATAIN[4]), .A2(n921), .B1(n922), .B2(\registers[28][4] ), .ZN(n1112) );
  AOI22_X2 U106 ( .A1(DATAIN[5]), .A2(n921), .B1(n923), .B2(\registers[28][5] ), .ZN(n1113) );
  AOI22_X2 U107 ( .A1(DATAIN[6]), .A2(n921), .B1(n923), .B2(\registers[28][6] ), .ZN(n1114) );
  AOI22_X2 U108 ( .A1(DATAIN[7]), .A2(n921), .B1(n923), .B2(\registers[28][7] ), .ZN(n1115) );
  AOI22_X2 U109 ( .A1(DATAIN[8]), .A2(n920), .B1(n923), .B2(\registers[28][8] ), .ZN(n1116) );
  AOI22_X2 U110 ( .A1(DATAIN[9]), .A2(n920), .B1(n923), .B2(\registers[28][9] ), .ZN(n1117) );
  AOI22_X2 U111 ( .A1(DATAIN[10]), .A2(n920), .B1(n924), .B2(
        \registers[28][10] ), .ZN(n1118) );
  AOI22_X2 U112 ( .A1(DATAIN[11]), .A2(n920), .B1(n924), .B2(
        \registers[28][11] ), .ZN(n1119) );
  AOI22_X2 U113 ( .A1(DATAIN[12]), .A2(n920), .B1(n924), .B2(
        \registers[28][12] ), .ZN(n1120) );
  AOI22_X2 U114 ( .A1(DATAIN[13]), .A2(n920), .B1(n924), .B2(
        \registers[28][13] ), .ZN(n1121) );
  AOI22_X2 U115 ( .A1(DATAIN[14]), .A2(n920), .B1(n924), .B2(
        \registers[28][14] ), .ZN(n1122) );
  AOI22_X2 U116 ( .A1(DATAIN[15]), .A2(n920), .B1(n925), .B2(
        \registers[28][15] ), .ZN(n1123) );
  AOI22_X2 U117 ( .A1(DATAIN[16]), .A2(n920), .B1(n925), .B2(
        \registers[28][16] ), .ZN(n1124) );
  AOI22_X2 U118 ( .A1(DATAIN[17]), .A2(n920), .B1(n925), .B2(
        \registers[28][17] ), .ZN(n1125) );
  AOI22_X2 U119 ( .A1(DATAIN[18]), .A2(n920), .B1(n925), .B2(
        \registers[28][18] ), .ZN(n1126) );
  AOI22_X2 U120 ( .A1(DATAIN[19]), .A2(n920), .B1(n925), .B2(
        \registers[28][19] ), .ZN(n1127) );
  AOI22_X2 U121 ( .A1(DATAIN[20]), .A2(n919), .B1(n926), .B2(
        \registers[28][20] ), .ZN(n1128) );
  AOI22_X2 U122 ( .A1(DATAIN[21]), .A2(n919), .B1(n926), .B2(
        \registers[28][21] ), .ZN(n1129) );
  AOI22_X2 U123 ( .A1(DATAIN[22]), .A2(n919), .B1(n926), .B2(
        \registers[28][22] ), .ZN(n1130) );
  AOI22_X2 U124 ( .A1(DATAIN[23]), .A2(n919), .B1(n926), .B2(
        \registers[28][23] ), .ZN(n1131) );
  AOI22_X2 U125 ( .A1(DATAIN[24]), .A2(n919), .B1(n926), .B2(
        \registers[28][24] ), .ZN(n1132) );
  AOI22_X2 U126 ( .A1(DATAIN[25]), .A2(n919), .B1(n927), .B2(
        \registers[28][25] ), .ZN(n1133) );
  AOI22_X2 U127 ( .A1(DATAIN[26]), .A2(n919), .B1(n927), .B2(
        \registers[28][26] ), .ZN(n1134) );
  AOI22_X2 U128 ( .A1(DATAIN[27]), .A2(n919), .B1(n927), .B2(
        \registers[28][27] ), .ZN(n1135) );
  AOI22_X2 U129 ( .A1(DATAIN[28]), .A2(n919), .B1(n927), .B2(
        \registers[28][28] ), .ZN(n1136) );
  AOI22_X2 U130 ( .A1(DATAIN[29]), .A2(n919), .B1(n927), .B2(
        \registers[28][29] ), .ZN(n1137) );
  AOI22_X2 U131 ( .A1(DATAIN[30]), .A2(n919), .B1(n928), .B2(
        \registers[28][30] ), .ZN(n1138) );
  AOI22_X2 U132 ( .A1(DATAIN[31]), .A2(n919), .B1(n928), .B2(
        \registers[28][31] ), .ZN(n1139) );
  NAND2_X2 U133 ( .A1(n1140), .A2(n1070), .ZN(n1108) );
  OAI22_X2 U134 ( .A1(n3890), .A2(n910), .B1(n911), .B2(n864), .ZN(n2838) );
  OAI22_X2 U135 ( .A1(n3889), .A2(n910), .B1(n911), .B2(n863), .ZN(n2839) );
  OAI22_X2 U136 ( .A1(n3888), .A2(n910), .B1(n911), .B2(n862), .ZN(n2840) );
  OAI22_X2 U137 ( .A1(n3887), .A2(n910), .B1(n911), .B2(n861), .ZN(n2841) );
  OAI22_X2 U138 ( .A1(n3886), .A2(n910), .B1(n911), .B2(n860), .ZN(n2842) );
  OAI22_X2 U139 ( .A1(n3885), .A2(n910), .B1(n912), .B2(n859), .ZN(n2843) );
  OAI22_X2 U140 ( .A1(n3884), .A2(n910), .B1(n912), .B2(n858), .ZN(n2844) );
  OAI22_X2 U141 ( .A1(n3883), .A2(n910), .B1(n912), .B2(n857), .ZN(n2845) );
  OAI22_X2 U142 ( .A1(n3882), .A2(n909), .B1(n912), .B2(n856), .ZN(n2846) );
  OAI22_X2 U143 ( .A1(n3881), .A2(n909), .B1(n912), .B2(n855), .ZN(n2847) );
  OAI22_X2 U144 ( .A1(n3880), .A2(n909), .B1(n913), .B2(n854), .ZN(n2848) );
  OAI22_X2 U145 ( .A1(n3879), .A2(n909), .B1(n913), .B2(n853), .ZN(n2849) );
  OAI22_X2 U146 ( .A1(n3878), .A2(n909), .B1(n913), .B2(n852), .ZN(n2850) );
  OAI22_X2 U147 ( .A1(n3877), .A2(n909), .B1(n913), .B2(n851), .ZN(n2851) );
  OAI22_X2 U148 ( .A1(n3876), .A2(n909), .B1(n913), .B2(n850), .ZN(n2852) );
  OAI22_X2 U149 ( .A1(n3875), .A2(n909), .B1(n914), .B2(n849), .ZN(n2853) );
  OAI22_X2 U150 ( .A1(n3874), .A2(n909), .B1(n914), .B2(n848), .ZN(n2854) );
  OAI22_X2 U151 ( .A1(n3873), .A2(n909), .B1(n914), .B2(n847), .ZN(n2855) );
  OAI22_X2 U152 ( .A1(n3872), .A2(n909), .B1(n914), .B2(n846), .ZN(n2856) );
  OAI22_X2 U153 ( .A1(n3871), .A2(n909), .B1(n914), .B2(n845), .ZN(n2857) );
  OAI22_X2 U154 ( .A1(n3870), .A2(n908), .B1(n915), .B2(n844), .ZN(n2858) );
  OAI22_X2 U155 ( .A1(n3869), .A2(n908), .B1(n915), .B2(n843), .ZN(n2859) );
  OAI22_X2 U156 ( .A1(n3868), .A2(n908), .B1(n915), .B2(n842), .ZN(n2860) );
  OAI22_X2 U157 ( .A1(n3867), .A2(n908), .B1(n915), .B2(n841), .ZN(n2861) );
  OAI22_X2 U158 ( .A1(n3866), .A2(n908), .B1(n915), .B2(n840), .ZN(n2862) );
  OAI22_X2 U159 ( .A1(n3865), .A2(n908), .B1(n916), .B2(n839), .ZN(n2863) );
  OAI22_X2 U160 ( .A1(n3864), .A2(n908), .B1(n916), .B2(n838), .ZN(n2864) );
  OAI22_X2 U161 ( .A1(n3863), .A2(n908), .B1(n916), .B2(n837), .ZN(n2865) );
  OAI22_X2 U162 ( .A1(n3862), .A2(n908), .B1(n916), .B2(n836), .ZN(n2866) );
  OAI22_X2 U163 ( .A1(n3861), .A2(n908), .B1(n916), .B2(n835), .ZN(n2867) );
  OAI22_X2 U164 ( .A1(n3860), .A2(n908), .B1(n917), .B2(n834), .ZN(n2868) );
  OAI22_X2 U165 ( .A1(n3859), .A2(n908), .B1(n917), .B2(n833), .ZN(n2869) );
  NAND2_X2 U166 ( .A1(n1142), .A2(n1070), .ZN(n1141) );
  OAI22_X2 U167 ( .A1(n3890), .A2(n899), .B1(n900), .B2(n832), .ZN(n2870) );
  OAI22_X2 U168 ( .A1(n3889), .A2(n899), .B1(n900), .B2(n831), .ZN(n2871) );
  OAI22_X2 U169 ( .A1(n3888), .A2(n899), .B1(n900), .B2(n830), .ZN(n2872) );
  OAI22_X2 U170 ( .A1(n3887), .A2(n899), .B1(n900), .B2(n829), .ZN(n2873) );
  OAI22_X2 U171 ( .A1(n3886), .A2(n899), .B1(n900), .B2(n828), .ZN(n2874) );
  OAI22_X2 U172 ( .A1(n3885), .A2(n899), .B1(n901), .B2(n827), .ZN(n2875) );
  OAI22_X2 U173 ( .A1(n3884), .A2(n899), .B1(n901), .B2(n826), .ZN(n2876) );
  OAI22_X2 U174 ( .A1(n3883), .A2(n899), .B1(n901), .B2(n825), .ZN(n2877) );
  OAI22_X2 U175 ( .A1(n3882), .A2(n898), .B1(n901), .B2(n824), .ZN(n2878) );
  OAI22_X2 U176 ( .A1(n3881), .A2(n898), .B1(n901), .B2(n823), .ZN(n2879) );
  OAI22_X2 U177 ( .A1(n3880), .A2(n898), .B1(n902), .B2(n822), .ZN(n2880) );
  OAI22_X2 U178 ( .A1(n3879), .A2(n898), .B1(n902), .B2(n821), .ZN(n2881) );
  OAI22_X2 U179 ( .A1(n3878), .A2(n898), .B1(n902), .B2(n820), .ZN(n2882) );
  OAI22_X2 U180 ( .A1(n3877), .A2(n898), .B1(n902), .B2(n819), .ZN(n2883) );
  OAI22_X2 U181 ( .A1(n3876), .A2(n898), .B1(n902), .B2(n818), .ZN(n2884) );
  OAI22_X2 U182 ( .A1(n3875), .A2(n898), .B1(n903), .B2(n817), .ZN(n2885) );
  OAI22_X2 U183 ( .A1(n3874), .A2(n898), .B1(n903), .B2(n816), .ZN(n2886) );
  OAI22_X2 U184 ( .A1(n3873), .A2(n898), .B1(n903), .B2(n815), .ZN(n2887) );
  OAI22_X2 U185 ( .A1(n3872), .A2(n898), .B1(n903), .B2(n814), .ZN(n2888) );
  OAI22_X2 U186 ( .A1(n3871), .A2(n898), .B1(n903), .B2(n813), .ZN(n2889) );
  OAI22_X2 U187 ( .A1(n3870), .A2(n897), .B1(n904), .B2(n812), .ZN(n2890) );
  OAI22_X2 U188 ( .A1(n3869), .A2(n897), .B1(n904), .B2(n811), .ZN(n2891) );
  OAI22_X2 U189 ( .A1(n3868), .A2(n897), .B1(n904), .B2(n810), .ZN(n2892) );
  OAI22_X2 U190 ( .A1(n3867), .A2(n897), .B1(n904), .B2(n809), .ZN(n2893) );
  OAI22_X2 U191 ( .A1(n3866), .A2(n897), .B1(n904), .B2(n808), .ZN(n2894) );
  OAI22_X2 U192 ( .A1(n3865), .A2(n897), .B1(n905), .B2(n807), .ZN(n2895) );
  OAI22_X2 U193 ( .A1(n3864), .A2(n897), .B1(n905), .B2(n806), .ZN(n2896) );
  OAI22_X2 U194 ( .A1(n3863), .A2(n897), .B1(n905), .B2(n805), .ZN(n2897) );
  OAI22_X2 U195 ( .A1(n3862), .A2(n897), .B1(n905), .B2(n804), .ZN(n2898) );
  OAI22_X2 U196 ( .A1(n3861), .A2(n897), .B1(n905), .B2(n803), .ZN(n2899) );
  OAI22_X2 U197 ( .A1(n3860), .A2(n897), .B1(n906), .B2(n802), .ZN(n2900) );
  OAI22_X2 U198 ( .A1(n3859), .A2(n897), .B1(n906), .B2(n801), .ZN(n2901) );
  NAND2_X2 U199 ( .A1(n1144), .A2(n1070), .ZN(n1143) );
  AOI22_X2 U200 ( .A1(DATAIN[0]), .A2(n889), .B1(n890), .B2(\registers[25][0] ), .ZN(n1145) );
  AOI22_X2 U201 ( .A1(DATAIN[1]), .A2(n889), .B1(n890), .B2(\registers[25][1] ), .ZN(n1147) );
  AOI22_X2 U202 ( .A1(DATAIN[2]), .A2(n889), .B1(n890), .B2(\registers[25][2] ), .ZN(n1148) );
  AOI22_X2 U203 ( .A1(DATAIN[3]), .A2(n889), .B1(n890), .B2(\registers[25][3] ), .ZN(n1149) );
  AOI22_X2 U204 ( .A1(DATAIN[4]), .A2(n889), .B1(n890), .B2(\registers[25][4] ), .ZN(n1150) );
  AOI22_X2 U205 ( .A1(DATAIN[5]), .A2(n889), .B1(n891), .B2(\registers[25][5] ), .ZN(n1151) );
  AOI22_X2 U206 ( .A1(DATAIN[6]), .A2(n889), .B1(n891), .B2(\registers[25][6] ), .ZN(n1152) );
  AOI22_X2 U207 ( .A1(DATAIN[7]), .A2(n889), .B1(n891), .B2(\registers[25][7] ), .ZN(n1153) );
  AOI22_X2 U208 ( .A1(DATAIN[8]), .A2(n888), .B1(n891), .B2(\registers[25][8] ), .ZN(n1154) );
  AOI22_X2 U209 ( .A1(DATAIN[9]), .A2(n888), .B1(n891), .B2(\registers[25][9] ), .ZN(n1155) );
  AOI22_X2 U210 ( .A1(DATAIN[10]), .A2(n888), .B1(n892), .B2(
        \registers[25][10] ), .ZN(n1156) );
  AOI22_X2 U211 ( .A1(DATAIN[11]), .A2(n888), .B1(n892), .B2(
        \registers[25][11] ), .ZN(n1157) );
  AOI22_X2 U212 ( .A1(DATAIN[12]), .A2(n888), .B1(n892), .B2(
        \registers[25][12] ), .ZN(n1158) );
  AOI22_X2 U213 ( .A1(DATAIN[13]), .A2(n888), .B1(n892), .B2(
        \registers[25][13] ), .ZN(n1159) );
  AOI22_X2 U214 ( .A1(DATAIN[14]), .A2(n888), .B1(n892), .B2(
        \registers[25][14] ), .ZN(n1160) );
  AOI22_X2 U215 ( .A1(DATAIN[15]), .A2(n888), .B1(n893), .B2(
        \registers[25][15] ), .ZN(n1161) );
  AOI22_X2 U216 ( .A1(DATAIN[16]), .A2(n888), .B1(n893), .B2(
        \registers[25][16] ), .ZN(n1162) );
  AOI22_X2 U217 ( .A1(DATAIN[17]), .A2(n888), .B1(n893), .B2(
        \registers[25][17] ), .ZN(n1163) );
  AOI22_X2 U218 ( .A1(DATAIN[18]), .A2(n888), .B1(n893), .B2(
        \registers[25][18] ), .ZN(n1164) );
  AOI22_X2 U219 ( .A1(DATAIN[19]), .A2(n888), .B1(n893), .B2(
        \registers[25][19] ), .ZN(n1165) );
  AOI22_X2 U220 ( .A1(DATAIN[20]), .A2(n887), .B1(n894), .B2(
        \registers[25][20] ), .ZN(n1166) );
  AOI22_X2 U221 ( .A1(DATAIN[21]), .A2(n887), .B1(n894), .B2(
        \registers[25][21] ), .ZN(n1167) );
  AOI22_X2 U222 ( .A1(DATAIN[22]), .A2(n887), .B1(n894), .B2(
        \registers[25][22] ), .ZN(n1168) );
  AOI22_X2 U223 ( .A1(DATAIN[23]), .A2(n887), .B1(n894), .B2(
        \registers[25][23] ), .ZN(n1169) );
  AOI22_X2 U224 ( .A1(DATAIN[24]), .A2(n887), .B1(n894), .B2(
        \registers[25][24] ), .ZN(n1170) );
  AOI22_X2 U225 ( .A1(DATAIN[25]), .A2(n887), .B1(n895), .B2(
        \registers[25][25] ), .ZN(n1171) );
  AOI22_X2 U226 ( .A1(DATAIN[26]), .A2(n887), .B1(n895), .B2(
        \registers[25][26] ), .ZN(n1172) );
  AOI22_X2 U227 ( .A1(DATAIN[27]), .A2(n887), .B1(n895), .B2(
        \registers[25][27] ), .ZN(n1173) );
  AOI22_X2 U228 ( .A1(DATAIN[28]), .A2(n887), .B1(n895), .B2(
        \registers[25][28] ), .ZN(n1174) );
  AOI22_X2 U229 ( .A1(DATAIN[29]), .A2(n887), .B1(n895), .B2(
        \registers[25][29] ), .ZN(n1175) );
  AOI22_X2 U230 ( .A1(DATAIN[30]), .A2(n887), .B1(n896), .B2(
        \registers[25][30] ), .ZN(n1176) );
  AOI22_X2 U231 ( .A1(DATAIN[31]), .A2(n887), .B1(n896), .B2(
        \registers[25][31] ), .ZN(n1177) );
  NAND2_X2 U232 ( .A1(n1178), .A2(n1070), .ZN(n1146) );
  AOI22_X2 U233 ( .A1(DATAIN[0]), .A2(n879), .B1(n880), .B2(\registers[24][0] ), .ZN(n1179) );
  AOI22_X2 U234 ( .A1(DATAIN[1]), .A2(n879), .B1(n880), .B2(\registers[24][1] ), .ZN(n1181) );
  AOI22_X2 U235 ( .A1(DATAIN[2]), .A2(n879), .B1(n880), .B2(\registers[24][2] ), .ZN(n1182) );
  AOI22_X2 U236 ( .A1(DATAIN[3]), .A2(n879), .B1(n880), .B2(\registers[24][3] ), .ZN(n1183) );
  AOI22_X2 U237 ( .A1(DATAIN[4]), .A2(n879), .B1(n880), .B2(\registers[24][4] ), .ZN(n1184) );
  AOI22_X2 U238 ( .A1(DATAIN[5]), .A2(n879), .B1(n881), .B2(\registers[24][5] ), .ZN(n1185) );
  AOI22_X2 U239 ( .A1(DATAIN[6]), .A2(n879), .B1(n881), .B2(\registers[24][6] ), .ZN(n1186) );
  AOI22_X2 U240 ( .A1(DATAIN[7]), .A2(n879), .B1(n881), .B2(\registers[24][7] ), .ZN(n1187) );
  AOI22_X2 U241 ( .A1(DATAIN[8]), .A2(n878), .B1(n881), .B2(\registers[24][8] ), .ZN(n1188) );
  AOI22_X2 U242 ( .A1(DATAIN[9]), .A2(n878), .B1(n881), .B2(\registers[24][9] ), .ZN(n1189) );
  AOI22_X2 U243 ( .A1(DATAIN[10]), .A2(n878), .B1(n882), .B2(
        \registers[24][10] ), .ZN(n1190) );
  AOI22_X2 U244 ( .A1(DATAIN[11]), .A2(n878), .B1(n882), .B2(
        \registers[24][11] ), .ZN(n1191) );
  AOI22_X2 U245 ( .A1(DATAIN[12]), .A2(n878), .B1(n882), .B2(
        \registers[24][12] ), .ZN(n1192) );
  AOI22_X2 U246 ( .A1(DATAIN[13]), .A2(n878), .B1(n882), .B2(
        \registers[24][13] ), .ZN(n1193) );
  AOI22_X2 U247 ( .A1(DATAIN[14]), .A2(n878), .B1(n882), .B2(
        \registers[24][14] ), .ZN(n1194) );
  AOI22_X2 U248 ( .A1(DATAIN[15]), .A2(n878), .B1(n883), .B2(
        \registers[24][15] ), .ZN(n1195) );
  AOI22_X2 U249 ( .A1(DATAIN[16]), .A2(n878), .B1(n883), .B2(
        \registers[24][16] ), .ZN(n1196) );
  AOI22_X2 U250 ( .A1(DATAIN[17]), .A2(n878), .B1(n883), .B2(
        \registers[24][17] ), .ZN(n1197) );
  AOI22_X2 U251 ( .A1(DATAIN[18]), .A2(n878), .B1(n883), .B2(
        \registers[24][18] ), .ZN(n1198) );
  AOI22_X2 U252 ( .A1(DATAIN[19]), .A2(n878), .B1(n883), .B2(
        \registers[24][19] ), .ZN(n1199) );
  AOI22_X2 U253 ( .A1(DATAIN[20]), .A2(n877), .B1(n884), .B2(
        \registers[24][20] ), .ZN(n1200) );
  AOI22_X2 U254 ( .A1(DATAIN[21]), .A2(n877), .B1(n884), .B2(
        \registers[24][21] ), .ZN(n1201) );
  AOI22_X2 U255 ( .A1(DATAIN[22]), .A2(n877), .B1(n884), .B2(
        \registers[24][22] ), .ZN(n1202) );
  AOI22_X2 U256 ( .A1(DATAIN[23]), .A2(n877), .B1(n884), .B2(
        \registers[24][23] ), .ZN(n1203) );
  AOI22_X2 U257 ( .A1(DATAIN[24]), .A2(n877), .B1(n884), .B2(
        \registers[24][24] ), .ZN(n1204) );
  AOI22_X2 U258 ( .A1(DATAIN[25]), .A2(n877), .B1(n885), .B2(
        \registers[24][25] ), .ZN(n1205) );
  AOI22_X2 U259 ( .A1(DATAIN[26]), .A2(n877), .B1(n885), .B2(
        \registers[24][26] ), .ZN(n1206) );
  AOI22_X2 U260 ( .A1(DATAIN[27]), .A2(n877), .B1(n885), .B2(
        \registers[24][27] ), .ZN(n1207) );
  AOI22_X2 U261 ( .A1(DATAIN[28]), .A2(n877), .B1(n885), .B2(
        \registers[24][28] ), .ZN(n1208) );
  AOI22_X2 U262 ( .A1(DATAIN[29]), .A2(n877), .B1(n885), .B2(
        \registers[24][29] ), .ZN(n1209) );
  AOI22_X2 U263 ( .A1(DATAIN[30]), .A2(n877), .B1(n886), .B2(
        \registers[24][30] ), .ZN(n1210) );
  AOI22_X2 U264 ( .A1(DATAIN[31]), .A2(n877), .B1(n886), .B2(
        \registers[24][31] ), .ZN(n1211) );
  NAND2_X2 U265 ( .A1(n1212), .A2(n1070), .ZN(n1180) );
  AND3_X2 U266 ( .A1(ADD_WR[3]), .A2(n1213), .A3(ADD_WR[4]), .ZN(n1070) );
  AOI22_X2 U267 ( .A1(DATAIN[0]), .A2(n869), .B1(n870), .B2(\registers[23][0] ), .ZN(n1214) );
  AOI22_X2 U268 ( .A1(DATAIN[1]), .A2(n869), .B1(n870), .B2(\registers[23][1] ), .ZN(n1216) );
  AOI22_X2 U269 ( .A1(DATAIN[2]), .A2(n869), .B1(n870), .B2(\registers[23][2] ), .ZN(n1217) );
  AOI22_X2 U270 ( .A1(DATAIN[3]), .A2(n869), .B1(n870), .B2(\registers[23][3] ), .ZN(n1218) );
  AOI22_X2 U271 ( .A1(DATAIN[4]), .A2(n869), .B1(n870), .B2(\registers[23][4] ), .ZN(n1219) );
  AOI22_X2 U272 ( .A1(DATAIN[5]), .A2(n869), .B1(n871), .B2(\registers[23][5] ), .ZN(n1220) );
  AOI22_X2 U273 ( .A1(DATAIN[6]), .A2(n869), .B1(n871), .B2(\registers[23][6] ), .ZN(n1221) );
  AOI22_X2 U274 ( .A1(DATAIN[7]), .A2(n869), .B1(n871), .B2(\registers[23][7] ), .ZN(n1222) );
  AOI22_X2 U275 ( .A1(DATAIN[8]), .A2(n868), .B1(n871), .B2(\registers[23][8] ), .ZN(n1223) );
  AOI22_X2 U276 ( .A1(DATAIN[9]), .A2(n868), .B1(n871), .B2(\registers[23][9] ), .ZN(n1224) );
  AOI22_X2 U277 ( .A1(DATAIN[10]), .A2(n868), .B1(n872), .B2(
        \registers[23][10] ), .ZN(n1225) );
  AOI22_X2 U278 ( .A1(DATAIN[11]), .A2(n868), .B1(n872), .B2(
        \registers[23][11] ), .ZN(n1226) );
  AOI22_X2 U279 ( .A1(DATAIN[12]), .A2(n868), .B1(n872), .B2(
        \registers[23][12] ), .ZN(n1227) );
  AOI22_X2 U280 ( .A1(DATAIN[13]), .A2(n868), .B1(n872), .B2(
        \registers[23][13] ), .ZN(n1228) );
  AOI22_X2 U281 ( .A1(DATAIN[14]), .A2(n868), .B1(n872), .B2(
        \registers[23][14] ), .ZN(n1229) );
  AOI22_X2 U282 ( .A1(DATAIN[15]), .A2(n868), .B1(n873), .B2(
        \registers[23][15] ), .ZN(n1230) );
  AOI22_X2 U283 ( .A1(DATAIN[16]), .A2(n868), .B1(n873), .B2(
        \registers[23][16] ), .ZN(n1231) );
  AOI22_X2 U284 ( .A1(DATAIN[17]), .A2(n868), .B1(n873), .B2(
        \registers[23][17] ), .ZN(n1232) );
  AOI22_X2 U285 ( .A1(DATAIN[18]), .A2(n868), .B1(n873), .B2(
        \registers[23][18] ), .ZN(n1233) );
  AOI22_X2 U286 ( .A1(DATAIN[19]), .A2(n868), .B1(n873), .B2(
        \registers[23][19] ), .ZN(n1234) );
  AOI22_X2 U287 ( .A1(DATAIN[20]), .A2(n867), .B1(n874), .B2(
        \registers[23][20] ), .ZN(n1235) );
  AOI22_X2 U288 ( .A1(DATAIN[21]), .A2(n867), .B1(n874), .B2(
        \registers[23][21] ), .ZN(n1236) );
  AOI22_X2 U289 ( .A1(DATAIN[22]), .A2(n867), .B1(n874), .B2(
        \registers[23][22] ), .ZN(n1237) );
  AOI22_X2 U290 ( .A1(DATAIN[23]), .A2(n867), .B1(n874), .B2(
        \registers[23][23] ), .ZN(n1238) );
  AOI22_X2 U291 ( .A1(DATAIN[24]), .A2(n867), .B1(n874), .B2(
        \registers[23][24] ), .ZN(n1239) );
  AOI22_X2 U292 ( .A1(DATAIN[25]), .A2(n867), .B1(n875), .B2(
        \registers[23][25] ), .ZN(n1240) );
  AOI22_X2 U293 ( .A1(DATAIN[26]), .A2(n867), .B1(n875), .B2(
        \registers[23][26] ), .ZN(n1241) );
  AOI22_X2 U294 ( .A1(DATAIN[27]), .A2(n867), .B1(n875), .B2(
        \registers[23][27] ), .ZN(n1242) );
  AOI22_X2 U295 ( .A1(DATAIN[28]), .A2(n867), .B1(n875), .B2(
        \registers[23][28] ), .ZN(n1243) );
  AOI22_X2 U296 ( .A1(DATAIN[29]), .A2(n867), .B1(n875), .B2(
        \registers[23][29] ), .ZN(n1244) );
  AOI22_X2 U297 ( .A1(DATAIN[30]), .A2(n867), .B1(n876), .B2(
        \registers[23][30] ), .ZN(n1245) );
  AOI22_X2 U298 ( .A1(DATAIN[31]), .A2(n867), .B1(n876), .B2(
        \registers[23][31] ), .ZN(n1246) );
  NAND2_X2 U299 ( .A1(n1247), .A2(n1069), .ZN(n1215) );
  AOI22_X2 U300 ( .A1(DATAIN[0]), .A2(n795), .B1(n796), .B2(\registers[22][0] ), .ZN(n1248) );
  AOI22_X2 U301 ( .A1(DATAIN[1]), .A2(n795), .B1(n796), .B2(\registers[22][1] ), .ZN(n1250) );
  AOI22_X2 U302 ( .A1(DATAIN[2]), .A2(n795), .B1(n796), .B2(\registers[22][2] ), .ZN(n1251) );
  AOI22_X2 U303 ( .A1(DATAIN[3]), .A2(n795), .B1(n796), .B2(\registers[22][3] ), .ZN(n1252) );
  AOI22_X2 U304 ( .A1(DATAIN[4]), .A2(n795), .B1(n796), .B2(\registers[22][4] ), .ZN(n1253) );
  AOI22_X2 U305 ( .A1(DATAIN[5]), .A2(n795), .B1(n797), .B2(\registers[22][5] ), .ZN(n1254) );
  AOI22_X2 U306 ( .A1(DATAIN[6]), .A2(n795), .B1(n797), .B2(\registers[22][6] ), .ZN(n1255) );
  AOI22_X2 U307 ( .A1(DATAIN[7]), .A2(n795), .B1(n797), .B2(\registers[22][7] ), .ZN(n1256) );
  AOI22_X2 U308 ( .A1(DATAIN[8]), .A2(n794), .B1(n797), .B2(\registers[22][8] ), .ZN(n1257) );
  AOI22_X2 U309 ( .A1(DATAIN[9]), .A2(n794), .B1(n797), .B2(\registers[22][9] ), .ZN(n1258) );
  AOI22_X2 U310 ( .A1(DATAIN[10]), .A2(n794), .B1(n798), .B2(
        \registers[22][10] ), .ZN(n1259) );
  AOI22_X2 U311 ( .A1(DATAIN[11]), .A2(n794), .B1(n798), .B2(
        \registers[22][11] ), .ZN(n1260) );
  AOI22_X2 U312 ( .A1(DATAIN[12]), .A2(n794), .B1(n798), .B2(
        \registers[22][12] ), .ZN(n1261) );
  AOI22_X2 U313 ( .A1(DATAIN[13]), .A2(n794), .B1(n798), .B2(
        \registers[22][13] ), .ZN(n1262) );
  AOI22_X2 U314 ( .A1(DATAIN[14]), .A2(n794), .B1(n798), .B2(
        \registers[22][14] ), .ZN(n1263) );
  AOI22_X2 U315 ( .A1(DATAIN[15]), .A2(n794), .B1(n799), .B2(
        \registers[22][15] ), .ZN(n1264) );
  AOI22_X2 U316 ( .A1(DATAIN[16]), .A2(n794), .B1(n799), .B2(
        \registers[22][16] ), .ZN(n1265) );
  AOI22_X2 U317 ( .A1(DATAIN[17]), .A2(n794), .B1(n799), .B2(
        \registers[22][17] ), .ZN(n1266) );
  AOI22_X2 U318 ( .A1(DATAIN[18]), .A2(n794), .B1(n799), .B2(
        \registers[22][18] ), .ZN(n1267) );
  AOI22_X2 U319 ( .A1(DATAIN[19]), .A2(n794), .B1(n799), .B2(
        \registers[22][19] ), .ZN(n1268) );
  AOI22_X2 U320 ( .A1(DATAIN[20]), .A2(n793), .B1(n800), .B2(
        \registers[22][20] ), .ZN(n1269) );
  AOI22_X2 U321 ( .A1(DATAIN[21]), .A2(n793), .B1(n800), .B2(
        \registers[22][21] ), .ZN(n1270) );
  AOI22_X2 U322 ( .A1(DATAIN[22]), .A2(n793), .B1(n800), .B2(
        \registers[22][22] ), .ZN(n1271) );
  AOI22_X2 U323 ( .A1(DATAIN[23]), .A2(n793), .B1(n800), .B2(
        \registers[22][23] ), .ZN(n1272) );
  AOI22_X2 U324 ( .A1(DATAIN[24]), .A2(n793), .B1(n800), .B2(
        \registers[22][24] ), .ZN(n1273) );
  AOI22_X2 U325 ( .A1(DATAIN[25]), .A2(n793), .B1(n865), .B2(
        \registers[22][25] ), .ZN(n1274) );
  AOI22_X2 U326 ( .A1(DATAIN[26]), .A2(n793), .B1(n865), .B2(
        \registers[22][26] ), .ZN(n1275) );
  AOI22_X2 U327 ( .A1(DATAIN[27]), .A2(n793), .B1(n865), .B2(
        \registers[22][27] ), .ZN(n1276) );
  AOI22_X2 U328 ( .A1(DATAIN[28]), .A2(n793), .B1(n865), .B2(
        \registers[22][28] ), .ZN(n1277) );
  AOI22_X2 U329 ( .A1(DATAIN[29]), .A2(n793), .B1(n865), .B2(
        \registers[22][29] ), .ZN(n1278) );
  AOI22_X2 U330 ( .A1(DATAIN[30]), .A2(n793), .B1(n866), .B2(
        \registers[22][30] ), .ZN(n1279) );
  AOI22_X2 U331 ( .A1(DATAIN[31]), .A2(n793), .B1(n866), .B2(
        \registers[22][31] ), .ZN(n1280) );
  NAND2_X2 U332 ( .A1(n1247), .A2(n1072), .ZN(n1249) );
  OAI22_X2 U333 ( .A1(n3890), .A2(n784), .B1(n785), .B2(n672), .ZN(n2902) );
  OAI22_X2 U334 ( .A1(n3889), .A2(n784), .B1(n785), .B2(n671), .ZN(n2903) );
  OAI22_X2 U335 ( .A1(n3888), .A2(n784), .B1(n785), .B2(n670), .ZN(n2904) );
  OAI22_X2 U336 ( .A1(n3887), .A2(n784), .B1(n785), .B2(n669), .ZN(n2905) );
  OAI22_X2 U337 ( .A1(n3886), .A2(n784), .B1(n785), .B2(n668), .ZN(n2906) );
  OAI22_X2 U338 ( .A1(n3885), .A2(n784), .B1(n786), .B2(n667), .ZN(n2907) );
  OAI22_X2 U339 ( .A1(n3884), .A2(n784), .B1(n786), .B2(n666), .ZN(n2908) );
  OAI22_X2 U340 ( .A1(n3883), .A2(n784), .B1(n786), .B2(n665), .ZN(n2909) );
  OAI22_X2 U341 ( .A1(n3882), .A2(n783), .B1(n786), .B2(n664), .ZN(n2910) );
  OAI22_X2 U342 ( .A1(n3881), .A2(n783), .B1(n786), .B2(n663), .ZN(n2911) );
  OAI22_X2 U343 ( .A1(n3880), .A2(n783), .B1(n787), .B2(n662), .ZN(n2912) );
  OAI22_X2 U344 ( .A1(n3879), .A2(n783), .B1(n787), .B2(n661), .ZN(n2913) );
  OAI22_X2 U345 ( .A1(n3878), .A2(n783), .B1(n787), .B2(n660), .ZN(n2914) );
  OAI22_X2 U346 ( .A1(n3877), .A2(n783), .B1(n787), .B2(n659), .ZN(n2915) );
  OAI22_X2 U347 ( .A1(n3876), .A2(n783), .B1(n787), .B2(n658), .ZN(n2916) );
  OAI22_X2 U348 ( .A1(n3875), .A2(n783), .B1(n788), .B2(n657), .ZN(n2917) );
  OAI22_X2 U349 ( .A1(n3874), .A2(n783), .B1(n788), .B2(n656), .ZN(n2918) );
  OAI22_X2 U350 ( .A1(n3873), .A2(n783), .B1(n788), .B2(n655), .ZN(n2919) );
  OAI22_X2 U351 ( .A1(n3872), .A2(n783), .B1(n788), .B2(n654), .ZN(n2920) );
  OAI22_X2 U352 ( .A1(n3871), .A2(n783), .B1(n788), .B2(n653), .ZN(n2921) );
  OAI22_X2 U353 ( .A1(n3870), .A2(n782), .B1(n789), .B2(n652), .ZN(n2922) );
  OAI22_X2 U354 ( .A1(n3869), .A2(n782), .B1(n789), .B2(n651), .ZN(n2923) );
  OAI22_X2 U355 ( .A1(n3868), .A2(n782), .B1(n789), .B2(n650), .ZN(n2924) );
  OAI22_X2 U356 ( .A1(n3867), .A2(n782), .B1(n789), .B2(n649), .ZN(n2925) );
  OAI22_X2 U357 ( .A1(n3866), .A2(n782), .B1(n789), .B2(n648), .ZN(n2926) );
  OAI22_X2 U358 ( .A1(n3865), .A2(n782), .B1(n790), .B2(n647), .ZN(n2927) );
  OAI22_X2 U359 ( .A1(n3864), .A2(n782), .B1(n790), .B2(n646), .ZN(n2928) );
  OAI22_X2 U360 ( .A1(n3863), .A2(n782), .B1(n790), .B2(n645), .ZN(n2929) );
  OAI22_X2 U361 ( .A1(n3862), .A2(n782), .B1(n790), .B2(n644), .ZN(n2930) );
  OAI22_X2 U362 ( .A1(n3861), .A2(n782), .B1(n790), .B2(n643), .ZN(n2931) );
  OAI22_X2 U363 ( .A1(n3860), .A2(n782), .B1(n791), .B2(n642), .ZN(n2932) );
  OAI22_X2 U364 ( .A1(n3859), .A2(n782), .B1(n791), .B2(n641), .ZN(n2933) );
  NAND2_X2 U365 ( .A1(n1247), .A2(n1106), .ZN(n1281) );
  OAI22_X2 U366 ( .A1(n3890), .A2(n773), .B1(n774), .B2(n640), .ZN(n2934) );
  OAI22_X2 U367 ( .A1(n3889), .A2(n773), .B1(n774), .B2(n639), .ZN(n2935) );
  OAI22_X2 U368 ( .A1(n3888), .A2(n773), .B1(n774), .B2(n638), .ZN(n2936) );
  OAI22_X2 U369 ( .A1(n3887), .A2(n773), .B1(n774), .B2(n637), .ZN(n2937) );
  OAI22_X2 U370 ( .A1(n3886), .A2(n773), .B1(n774), .B2(n636), .ZN(n2938) );
  OAI22_X2 U371 ( .A1(n3885), .A2(n773), .B1(n775), .B2(n635), .ZN(n2939) );
  OAI22_X2 U372 ( .A1(n3884), .A2(n773), .B1(n775), .B2(n634), .ZN(n2940) );
  OAI22_X2 U373 ( .A1(n3883), .A2(n773), .B1(n775), .B2(n633), .ZN(n2941) );
  OAI22_X2 U374 ( .A1(n3882), .A2(n772), .B1(n775), .B2(n632), .ZN(n2942) );
  OAI22_X2 U375 ( .A1(n3881), .A2(n772), .B1(n775), .B2(n631), .ZN(n2943) );
  OAI22_X2 U376 ( .A1(n3880), .A2(n772), .B1(n776), .B2(n630), .ZN(n2944) );
  OAI22_X2 U377 ( .A1(n3879), .A2(n772), .B1(n776), .B2(n629), .ZN(n2945) );
  OAI22_X2 U378 ( .A1(n3878), .A2(n772), .B1(n776), .B2(n628), .ZN(n2946) );
  OAI22_X2 U379 ( .A1(n3877), .A2(n772), .B1(n776), .B2(n627), .ZN(n2947) );
  OAI22_X2 U380 ( .A1(n3876), .A2(n772), .B1(n776), .B2(n626), .ZN(n2948) );
  OAI22_X2 U381 ( .A1(n3875), .A2(n772), .B1(n777), .B2(n625), .ZN(n2949) );
  OAI22_X2 U382 ( .A1(n3874), .A2(n772), .B1(n777), .B2(n624), .ZN(n2950) );
  OAI22_X2 U383 ( .A1(n3873), .A2(n772), .B1(n777), .B2(n623), .ZN(n2951) );
  OAI22_X2 U384 ( .A1(n3872), .A2(n772), .B1(n777), .B2(n622), .ZN(n2952) );
  OAI22_X2 U385 ( .A1(n3871), .A2(n772), .B1(n777), .B2(n621), .ZN(n2953) );
  OAI22_X2 U386 ( .A1(n3870), .A2(n771), .B1(n778), .B2(n620), .ZN(n2954) );
  OAI22_X2 U387 ( .A1(n3869), .A2(n771), .B1(n778), .B2(n619), .ZN(n2955) );
  OAI22_X2 U388 ( .A1(n3868), .A2(n771), .B1(n778), .B2(n618), .ZN(n2956) );
  OAI22_X2 U389 ( .A1(n3867), .A2(n771), .B1(n778), .B2(n617), .ZN(n2957) );
  OAI22_X2 U390 ( .A1(n3866), .A2(n771), .B1(n778), .B2(n616), .ZN(n2958) );
  OAI22_X2 U391 ( .A1(n3865), .A2(n771), .B1(n779), .B2(n615), .ZN(n2959) );
  OAI22_X2 U392 ( .A1(n3864), .A2(n771), .B1(n779), .B2(n614), .ZN(n2960) );
  OAI22_X2 U393 ( .A1(n3863), .A2(n771), .B1(n779), .B2(n613), .ZN(n2961) );
  OAI22_X2 U394 ( .A1(n3862), .A2(n771), .B1(n779), .B2(n612), .ZN(n2962) );
  OAI22_X2 U395 ( .A1(n3861), .A2(n771), .B1(n779), .B2(n611), .ZN(n2963) );
  OAI22_X2 U396 ( .A1(n3860), .A2(n771), .B1(n780), .B2(n610), .ZN(n2964) );
  OAI22_X2 U397 ( .A1(n3859), .A2(n771), .B1(n780), .B2(n609), .ZN(n2965) );
  NAND2_X2 U398 ( .A1(n1247), .A2(n1140), .ZN(n1282) );
  AOI22_X2 U399 ( .A1(DATAIN[0]), .A2(n763), .B1(n764), .B2(\registers[19][0] ), .ZN(n1283) );
  AOI22_X2 U400 ( .A1(DATAIN[1]), .A2(n763), .B1(n764), .B2(\registers[19][1] ), .ZN(n1285) );
  AOI22_X2 U401 ( .A1(DATAIN[2]), .A2(n763), .B1(n764), .B2(\registers[19][2] ), .ZN(n1286) );
  AOI22_X2 U402 ( .A1(DATAIN[3]), .A2(n763), .B1(n764), .B2(\registers[19][3] ), .ZN(n1287) );
  AOI22_X2 U403 ( .A1(DATAIN[4]), .A2(n763), .B1(n764), .B2(\registers[19][4] ), .ZN(n1288) );
  AOI22_X2 U404 ( .A1(DATAIN[5]), .A2(n763), .B1(n765), .B2(\registers[19][5] ), .ZN(n1289) );
  AOI22_X2 U405 ( .A1(DATAIN[6]), .A2(n763), .B1(n765), .B2(\registers[19][6] ), .ZN(n1290) );
  AOI22_X2 U406 ( .A1(DATAIN[7]), .A2(n763), .B1(n765), .B2(\registers[19][7] ), .ZN(n1291) );
  AOI22_X2 U407 ( .A1(DATAIN[8]), .A2(n762), .B1(n765), .B2(\registers[19][8] ), .ZN(n1292) );
  AOI22_X2 U408 ( .A1(DATAIN[9]), .A2(n762), .B1(n765), .B2(\registers[19][9] ), .ZN(n1293) );
  AOI22_X2 U409 ( .A1(DATAIN[10]), .A2(n762), .B1(n766), .B2(
        \registers[19][10] ), .ZN(n1294) );
  AOI22_X2 U410 ( .A1(DATAIN[11]), .A2(n762), .B1(n766), .B2(
        \registers[19][11] ), .ZN(n1295) );
  AOI22_X2 U411 ( .A1(DATAIN[12]), .A2(n762), .B1(n766), .B2(
        \registers[19][12] ), .ZN(n1296) );
  AOI22_X2 U412 ( .A1(DATAIN[13]), .A2(n762), .B1(n766), .B2(
        \registers[19][13] ), .ZN(n1297) );
  AOI22_X2 U413 ( .A1(DATAIN[14]), .A2(n762), .B1(n766), .B2(
        \registers[19][14] ), .ZN(n1298) );
  AOI22_X2 U414 ( .A1(DATAIN[15]), .A2(n762), .B1(n767), .B2(
        \registers[19][15] ), .ZN(n1299) );
  AOI22_X2 U415 ( .A1(DATAIN[16]), .A2(n762), .B1(n767), .B2(
        \registers[19][16] ), .ZN(n1300) );
  AOI22_X2 U416 ( .A1(DATAIN[17]), .A2(n762), .B1(n767), .B2(
        \registers[19][17] ), .ZN(n1301) );
  AOI22_X2 U417 ( .A1(DATAIN[18]), .A2(n762), .B1(n767), .B2(
        \registers[19][18] ), .ZN(n1302) );
  AOI22_X2 U418 ( .A1(DATAIN[19]), .A2(n762), .B1(n767), .B2(
        \registers[19][19] ), .ZN(n1303) );
  AOI22_X2 U419 ( .A1(DATAIN[20]), .A2(n761), .B1(n768), .B2(
        \registers[19][20] ), .ZN(n1304) );
  AOI22_X2 U420 ( .A1(DATAIN[21]), .A2(n761), .B1(n768), .B2(
        \registers[19][21] ), .ZN(n1305) );
  AOI22_X2 U421 ( .A1(DATAIN[22]), .A2(n761), .B1(n768), .B2(
        \registers[19][22] ), .ZN(n1306) );
  AOI22_X2 U422 ( .A1(DATAIN[23]), .A2(n761), .B1(n768), .B2(
        \registers[19][23] ), .ZN(n1307) );
  AOI22_X2 U423 ( .A1(DATAIN[24]), .A2(n761), .B1(n768), .B2(
        \registers[19][24] ), .ZN(n1308) );
  AOI22_X2 U424 ( .A1(DATAIN[25]), .A2(n761), .B1(n769), .B2(
        \registers[19][25] ), .ZN(n1309) );
  AOI22_X2 U425 ( .A1(DATAIN[26]), .A2(n761), .B1(n769), .B2(
        \registers[19][26] ), .ZN(n1310) );
  AOI22_X2 U426 ( .A1(DATAIN[27]), .A2(n761), .B1(n769), .B2(
        \registers[19][27] ), .ZN(n1311) );
  AOI22_X2 U427 ( .A1(DATAIN[28]), .A2(n761), .B1(n769), .B2(
        \registers[19][28] ), .ZN(n1312) );
  AOI22_X2 U428 ( .A1(DATAIN[29]), .A2(n761), .B1(n769), .B2(
        \registers[19][29] ), .ZN(n1313) );
  AOI22_X2 U429 ( .A1(DATAIN[30]), .A2(n761), .B1(n770), .B2(
        \registers[19][30] ), .ZN(n1314) );
  AOI22_X2 U430 ( .A1(DATAIN[31]), .A2(n761), .B1(n770), .B2(
        \registers[19][31] ), .ZN(n1315) );
  NAND2_X2 U431 ( .A1(n1247), .A2(n1142), .ZN(n1284) );
  AOI22_X2 U432 ( .A1(DATAIN[0]), .A2(n753), .B1(n754), .B2(\registers[18][0] ), .ZN(n1316) );
  AOI22_X2 U433 ( .A1(DATAIN[1]), .A2(n753), .B1(n754), .B2(\registers[18][1] ), .ZN(n1318) );
  AOI22_X2 U434 ( .A1(DATAIN[2]), .A2(n753), .B1(n754), .B2(\registers[18][2] ), .ZN(n1319) );
  AOI22_X2 U435 ( .A1(DATAIN[3]), .A2(n753), .B1(n754), .B2(\registers[18][3] ), .ZN(n1320) );
  AOI22_X2 U436 ( .A1(DATAIN[4]), .A2(n753), .B1(n754), .B2(\registers[18][4] ), .ZN(n1321) );
  AOI22_X2 U437 ( .A1(DATAIN[5]), .A2(n753), .B1(n755), .B2(\registers[18][5] ), .ZN(n1322) );
  AOI22_X2 U438 ( .A1(DATAIN[6]), .A2(n753), .B1(n755), .B2(\registers[18][6] ), .ZN(n1323) );
  AOI22_X2 U439 ( .A1(DATAIN[7]), .A2(n753), .B1(n755), .B2(\registers[18][7] ), .ZN(n1324) );
  AOI22_X2 U440 ( .A1(DATAIN[8]), .A2(n752), .B1(n755), .B2(\registers[18][8] ), .ZN(n1325) );
  AOI22_X2 U441 ( .A1(DATAIN[9]), .A2(n752), .B1(n755), .B2(\registers[18][9] ), .ZN(n1326) );
  AOI22_X2 U442 ( .A1(DATAIN[10]), .A2(n752), .B1(n756), .B2(
        \registers[18][10] ), .ZN(n1327) );
  AOI22_X2 U443 ( .A1(DATAIN[11]), .A2(n752), .B1(n756), .B2(
        \registers[18][11] ), .ZN(n1328) );
  AOI22_X2 U444 ( .A1(DATAIN[12]), .A2(n752), .B1(n756), .B2(
        \registers[18][12] ), .ZN(n1329) );
  AOI22_X2 U445 ( .A1(DATAIN[13]), .A2(n752), .B1(n756), .B2(
        \registers[18][13] ), .ZN(n1330) );
  AOI22_X2 U446 ( .A1(DATAIN[14]), .A2(n752), .B1(n756), .B2(
        \registers[18][14] ), .ZN(n1331) );
  AOI22_X2 U447 ( .A1(DATAIN[15]), .A2(n752), .B1(n757), .B2(
        \registers[18][15] ), .ZN(n1332) );
  AOI22_X2 U448 ( .A1(DATAIN[16]), .A2(n752), .B1(n757), .B2(
        \registers[18][16] ), .ZN(n1333) );
  AOI22_X2 U449 ( .A1(DATAIN[17]), .A2(n752), .B1(n757), .B2(
        \registers[18][17] ), .ZN(n1334) );
  AOI22_X2 U450 ( .A1(DATAIN[18]), .A2(n752), .B1(n757), .B2(
        \registers[18][18] ), .ZN(n1335) );
  AOI22_X2 U451 ( .A1(DATAIN[19]), .A2(n752), .B1(n757), .B2(
        \registers[18][19] ), .ZN(n1336) );
  AOI22_X2 U452 ( .A1(DATAIN[20]), .A2(n751), .B1(n758), .B2(
        \registers[18][20] ), .ZN(n1337) );
  AOI22_X2 U453 ( .A1(DATAIN[21]), .A2(n751), .B1(n758), .B2(
        \registers[18][21] ), .ZN(n1338) );
  AOI22_X2 U454 ( .A1(DATAIN[22]), .A2(n751), .B1(n758), .B2(
        \registers[18][22] ), .ZN(n1339) );
  AOI22_X2 U455 ( .A1(DATAIN[23]), .A2(n751), .B1(n758), .B2(
        \registers[18][23] ), .ZN(n1340) );
  AOI22_X2 U456 ( .A1(DATAIN[24]), .A2(n751), .B1(n758), .B2(
        \registers[18][24] ), .ZN(n1341) );
  AOI22_X2 U457 ( .A1(DATAIN[25]), .A2(n751), .B1(n759), .B2(
        \registers[18][25] ), .ZN(n1342) );
  AOI22_X2 U458 ( .A1(DATAIN[26]), .A2(n751), .B1(n759), .B2(
        \registers[18][26] ), .ZN(n1343) );
  AOI22_X2 U459 ( .A1(DATAIN[27]), .A2(n751), .B1(n759), .B2(
        \registers[18][27] ), .ZN(n1344) );
  AOI22_X2 U460 ( .A1(DATAIN[28]), .A2(n751), .B1(n759), .B2(
        \registers[18][28] ), .ZN(n1345) );
  AOI22_X2 U461 ( .A1(DATAIN[29]), .A2(n751), .B1(n759), .B2(
        \registers[18][29] ), .ZN(n1346) );
  AOI22_X2 U462 ( .A1(DATAIN[30]), .A2(n751), .B1(n760), .B2(
        \registers[18][30] ), .ZN(n1347) );
  AOI22_X2 U463 ( .A1(DATAIN[31]), .A2(n751), .B1(n760), .B2(
        \registers[18][31] ), .ZN(n1348) );
  NAND2_X2 U464 ( .A1(n1247), .A2(n1144), .ZN(n1317) );
  OAI22_X2 U465 ( .A1(n3890), .A2(n742), .B1(n743), .B2(n544), .ZN(n2966) );
  OAI22_X2 U466 ( .A1(n3889), .A2(n742), .B1(n743), .B2(n543), .ZN(n2967) );
  OAI22_X2 U467 ( .A1(n3888), .A2(n742), .B1(n743), .B2(n542), .ZN(n2968) );
  OAI22_X2 U468 ( .A1(n3887), .A2(n742), .B1(n743), .B2(n541), .ZN(n2969) );
  OAI22_X2 U469 ( .A1(n3886), .A2(n742), .B1(n743), .B2(n540), .ZN(n2970) );
  OAI22_X2 U470 ( .A1(n3885), .A2(n742), .B1(n744), .B2(n539), .ZN(n2971) );
  OAI22_X2 U471 ( .A1(n3884), .A2(n742), .B1(n744), .B2(n538), .ZN(n2972) );
  OAI22_X2 U472 ( .A1(n3883), .A2(n742), .B1(n744), .B2(n537), .ZN(n2973) );
  OAI22_X2 U473 ( .A1(n3882), .A2(n741), .B1(n744), .B2(n536), .ZN(n2974) );
  OAI22_X2 U474 ( .A1(n3881), .A2(n741), .B1(n744), .B2(n535), .ZN(n2975) );
  OAI22_X2 U475 ( .A1(n3880), .A2(n741), .B1(n745), .B2(n534), .ZN(n2976) );
  OAI22_X2 U476 ( .A1(n3879), .A2(n741), .B1(n745), .B2(n533), .ZN(n2977) );
  OAI22_X2 U477 ( .A1(n3878), .A2(n741), .B1(n745), .B2(n532), .ZN(n2978) );
  OAI22_X2 U478 ( .A1(n3877), .A2(n741), .B1(n745), .B2(n531), .ZN(n2979) );
  OAI22_X2 U479 ( .A1(n3876), .A2(n741), .B1(n745), .B2(n530), .ZN(n2980) );
  OAI22_X2 U480 ( .A1(n3875), .A2(n741), .B1(n746), .B2(n529), .ZN(n2981) );
  OAI22_X2 U481 ( .A1(n3874), .A2(n741), .B1(n746), .B2(n528), .ZN(n2982) );
  OAI22_X2 U482 ( .A1(n3873), .A2(n741), .B1(n746), .B2(n527), .ZN(n2983) );
  OAI22_X2 U483 ( .A1(n3872), .A2(n741), .B1(n746), .B2(n526), .ZN(n2984) );
  OAI22_X2 U484 ( .A1(n3871), .A2(n741), .B1(n746), .B2(n525), .ZN(n2985) );
  OAI22_X2 U485 ( .A1(n3870), .A2(n740), .B1(n747), .B2(n524), .ZN(n2986) );
  OAI22_X2 U486 ( .A1(n3869), .A2(n740), .B1(n747), .B2(n523), .ZN(n2987) );
  OAI22_X2 U487 ( .A1(n3868), .A2(n740), .B1(n747), .B2(n522), .ZN(n2988) );
  OAI22_X2 U488 ( .A1(n3867), .A2(n740), .B1(n747), .B2(n521), .ZN(n2989) );
  OAI22_X2 U489 ( .A1(n3866), .A2(n740), .B1(n747), .B2(n520), .ZN(n2990) );
  OAI22_X2 U490 ( .A1(n3865), .A2(n740), .B1(n748), .B2(n519), .ZN(n2991) );
  OAI22_X2 U491 ( .A1(n3864), .A2(n740), .B1(n748), .B2(n518), .ZN(n2992) );
  OAI22_X2 U492 ( .A1(n3863), .A2(n740), .B1(n748), .B2(n517), .ZN(n2993) );
  OAI22_X2 U493 ( .A1(n3862), .A2(n740), .B1(n748), .B2(n516), .ZN(n2994) );
  OAI22_X2 U494 ( .A1(n3861), .A2(n740), .B1(n748), .B2(n515), .ZN(n2995) );
  OAI22_X2 U495 ( .A1(n3860), .A2(n740), .B1(n749), .B2(n514), .ZN(n2996) );
  OAI22_X2 U496 ( .A1(n3859), .A2(n740), .B1(n749), .B2(n513), .ZN(n2997) );
  NAND2_X2 U497 ( .A1(n1247), .A2(n1178), .ZN(n1349) );
  OAI22_X2 U498 ( .A1(n3890), .A2(n731), .B1(n732), .B2(n512), .ZN(n2998) );
  OAI22_X2 U499 ( .A1(n3889), .A2(n731), .B1(n732), .B2(n511), .ZN(n2999) );
  OAI22_X2 U500 ( .A1(n3888), .A2(n731), .B1(n732), .B2(n510), .ZN(n3000) );
  OAI22_X2 U501 ( .A1(n3887), .A2(n731), .B1(n732), .B2(n509), .ZN(n3001) );
  OAI22_X2 U502 ( .A1(n3886), .A2(n731), .B1(n732), .B2(n508), .ZN(n3002) );
  OAI22_X2 U503 ( .A1(n3885), .A2(n731), .B1(n733), .B2(n507), .ZN(n3003) );
  OAI22_X2 U504 ( .A1(n3884), .A2(n731), .B1(n733), .B2(n506), .ZN(n3004) );
  OAI22_X2 U505 ( .A1(n3883), .A2(n731), .B1(n733), .B2(n505), .ZN(n3005) );
  OAI22_X2 U506 ( .A1(n3882), .A2(n730), .B1(n733), .B2(n504), .ZN(n3006) );
  OAI22_X2 U507 ( .A1(n3881), .A2(n730), .B1(n733), .B2(n503), .ZN(n3007) );
  OAI22_X2 U508 ( .A1(n3880), .A2(n730), .B1(n734), .B2(n502), .ZN(n3008) );
  OAI22_X2 U509 ( .A1(n3879), .A2(n730), .B1(n734), .B2(n501), .ZN(n3009) );
  OAI22_X2 U510 ( .A1(n3878), .A2(n730), .B1(n734), .B2(n500), .ZN(n3010) );
  OAI22_X2 U511 ( .A1(n3877), .A2(n730), .B1(n734), .B2(n499), .ZN(n3011) );
  OAI22_X2 U512 ( .A1(n3876), .A2(n730), .B1(n734), .B2(n498), .ZN(n3012) );
  OAI22_X2 U513 ( .A1(n3875), .A2(n730), .B1(n735), .B2(n497), .ZN(n3013) );
  OAI22_X2 U514 ( .A1(n3874), .A2(n730), .B1(n735), .B2(n496), .ZN(n3014) );
  OAI22_X2 U515 ( .A1(n3873), .A2(n730), .B1(n735), .B2(n495), .ZN(n3015) );
  OAI22_X2 U516 ( .A1(n3872), .A2(n730), .B1(n735), .B2(n494), .ZN(n3016) );
  OAI22_X2 U517 ( .A1(n3871), .A2(n730), .B1(n735), .B2(n493), .ZN(n3017) );
  OAI22_X2 U518 ( .A1(n3870), .A2(n729), .B1(n736), .B2(n492), .ZN(n3018) );
  OAI22_X2 U519 ( .A1(n3869), .A2(n729), .B1(n736), .B2(n491), .ZN(n3019) );
  OAI22_X2 U520 ( .A1(n3868), .A2(n729), .B1(n736), .B2(n490), .ZN(n3020) );
  OAI22_X2 U521 ( .A1(n3867), .A2(n729), .B1(n736), .B2(n489), .ZN(n3021) );
  OAI22_X2 U522 ( .A1(n3866), .A2(n729), .B1(n736), .B2(n488), .ZN(n3022) );
  OAI22_X2 U523 ( .A1(n3865), .A2(n729), .B1(n737), .B2(n487), .ZN(n3023) );
  OAI22_X2 U524 ( .A1(n3864), .A2(n729), .B1(n737), .B2(n486), .ZN(n3024) );
  OAI22_X2 U525 ( .A1(n3863), .A2(n729), .B1(n737), .B2(n485), .ZN(n3025) );
  OAI22_X2 U526 ( .A1(n3862), .A2(n729), .B1(n737), .B2(n484), .ZN(n3026) );
  OAI22_X2 U527 ( .A1(n3861), .A2(n729), .B1(n737), .B2(n483), .ZN(n3027) );
  OAI22_X2 U528 ( .A1(n3860), .A2(n729), .B1(n738), .B2(n482), .ZN(n3028) );
  OAI22_X2 U529 ( .A1(n3859), .A2(n729), .B1(n738), .B2(n481), .ZN(n3029) );
  NAND2_X2 U530 ( .A1(n1247), .A2(n1212), .ZN(n1350) );
  AND3_X2 U531 ( .A1(n1213), .A2(n3849), .A3(ADD_WR[4]), .ZN(n1247) );
  OAI22_X2 U532 ( .A1(n3890), .A2(n720), .B1(n721), .B2(n480), .ZN(n3030) );
  OAI22_X2 U533 ( .A1(n3889), .A2(n720), .B1(n721), .B2(n479), .ZN(n3031) );
  OAI22_X2 U534 ( .A1(n3888), .A2(n720), .B1(n721), .B2(n478), .ZN(n3032) );
  OAI22_X2 U535 ( .A1(n3887), .A2(n720), .B1(n721), .B2(n477), .ZN(n3033) );
  OAI22_X2 U536 ( .A1(n3886), .A2(n720), .B1(n721), .B2(n476), .ZN(n3034) );
  OAI22_X2 U537 ( .A1(n3885), .A2(n720), .B1(n722), .B2(n475), .ZN(n3035) );
  OAI22_X2 U538 ( .A1(n3884), .A2(n720), .B1(n722), .B2(n474), .ZN(n3036) );
  OAI22_X2 U539 ( .A1(n3883), .A2(n720), .B1(n722), .B2(n473), .ZN(n3037) );
  OAI22_X2 U540 ( .A1(n3882), .A2(n719), .B1(n722), .B2(n472), .ZN(n3038) );
  OAI22_X2 U541 ( .A1(n3881), .A2(n719), .B1(n722), .B2(n471), .ZN(n3039) );
  OAI22_X2 U542 ( .A1(n3880), .A2(n719), .B1(n723), .B2(n470), .ZN(n3040) );
  OAI22_X2 U543 ( .A1(n3879), .A2(n719), .B1(n723), .B2(n469), .ZN(n3041) );
  OAI22_X2 U544 ( .A1(n3878), .A2(n719), .B1(n723), .B2(n468), .ZN(n3042) );
  OAI22_X2 U545 ( .A1(n3877), .A2(n719), .B1(n723), .B2(n467), .ZN(n3043) );
  OAI22_X2 U546 ( .A1(n3876), .A2(n719), .B1(n723), .B2(n466), .ZN(n3044) );
  OAI22_X2 U547 ( .A1(n3875), .A2(n719), .B1(n724), .B2(n465), .ZN(n3045) );
  OAI22_X2 U548 ( .A1(n3874), .A2(n719), .B1(n724), .B2(n464), .ZN(n3046) );
  OAI22_X2 U549 ( .A1(n3873), .A2(n719), .B1(n724), .B2(n463), .ZN(n3047) );
  OAI22_X2 U550 ( .A1(n3872), .A2(n719), .B1(n724), .B2(n462), .ZN(n3048) );
  OAI22_X2 U551 ( .A1(n3871), .A2(n719), .B1(n724), .B2(n461), .ZN(n3049) );
  OAI22_X2 U552 ( .A1(n3870), .A2(n718), .B1(n725), .B2(n460), .ZN(n3050) );
  OAI22_X2 U553 ( .A1(n3869), .A2(n718), .B1(n725), .B2(n459), .ZN(n3051) );
  OAI22_X2 U554 ( .A1(n3868), .A2(n718), .B1(n725), .B2(n458), .ZN(n3052) );
  OAI22_X2 U555 ( .A1(n3867), .A2(n718), .B1(n725), .B2(n457), .ZN(n3053) );
  OAI22_X2 U556 ( .A1(n3866), .A2(n718), .B1(n725), .B2(n456), .ZN(n3054) );
  OAI22_X2 U557 ( .A1(n3865), .A2(n718), .B1(n726), .B2(n455), .ZN(n3055) );
  OAI22_X2 U558 ( .A1(n3864), .A2(n718), .B1(n726), .B2(n454), .ZN(n3056) );
  OAI22_X2 U559 ( .A1(n3863), .A2(n718), .B1(n726), .B2(n453), .ZN(n3057) );
  OAI22_X2 U560 ( .A1(n3862), .A2(n718), .B1(n726), .B2(n452), .ZN(n3058) );
  OAI22_X2 U561 ( .A1(n3861), .A2(n718), .B1(n726), .B2(n451), .ZN(n3059) );
  OAI22_X2 U562 ( .A1(n3860), .A2(n718), .B1(n727), .B2(n450), .ZN(n3060) );
  OAI22_X2 U563 ( .A1(n3859), .A2(n718), .B1(n727), .B2(n449), .ZN(n3061) );
  NAND2_X2 U564 ( .A1(n1352), .A2(n1069), .ZN(n1351) );
  OAI22_X2 U565 ( .A1(n3890), .A2(n709), .B1(n710), .B2(n448), .ZN(n3062) );
  OAI22_X2 U566 ( .A1(n3889), .A2(n709), .B1(n710), .B2(n447), .ZN(n3063) );
  OAI22_X2 U567 ( .A1(n3888), .A2(n709), .B1(n710), .B2(n446), .ZN(n3064) );
  OAI22_X2 U568 ( .A1(n3887), .A2(n709), .B1(n710), .B2(n445), .ZN(n3065) );
  OAI22_X2 U569 ( .A1(n3886), .A2(n709), .B1(n710), .B2(n444), .ZN(n3066) );
  OAI22_X2 U570 ( .A1(n3885), .A2(n709), .B1(n711), .B2(n443), .ZN(n3067) );
  OAI22_X2 U571 ( .A1(n3884), .A2(n709), .B1(n711), .B2(n442), .ZN(n3068) );
  OAI22_X2 U572 ( .A1(n3883), .A2(n709), .B1(n711), .B2(n441), .ZN(n3069) );
  OAI22_X2 U573 ( .A1(n3882), .A2(n708), .B1(n711), .B2(n440), .ZN(n3070) );
  OAI22_X2 U574 ( .A1(n3881), .A2(n708), .B1(n711), .B2(n439), .ZN(n3071) );
  OAI22_X2 U575 ( .A1(n3880), .A2(n708), .B1(n712), .B2(n438), .ZN(n3072) );
  OAI22_X2 U576 ( .A1(n3879), .A2(n708), .B1(n712), .B2(n437), .ZN(n3073) );
  OAI22_X2 U577 ( .A1(n3878), .A2(n708), .B1(n712), .B2(n436), .ZN(n3074) );
  OAI22_X2 U578 ( .A1(n3877), .A2(n708), .B1(n712), .B2(n435), .ZN(n3075) );
  OAI22_X2 U579 ( .A1(n3876), .A2(n708), .B1(n712), .B2(n434), .ZN(n3076) );
  OAI22_X2 U580 ( .A1(n3875), .A2(n708), .B1(n713), .B2(n433), .ZN(n3077) );
  OAI22_X2 U581 ( .A1(n3874), .A2(n708), .B1(n713), .B2(n432), .ZN(n3078) );
  OAI22_X2 U582 ( .A1(n3873), .A2(n708), .B1(n713), .B2(n431), .ZN(n3079) );
  OAI22_X2 U583 ( .A1(n3872), .A2(n708), .B1(n713), .B2(n430), .ZN(n3080) );
  OAI22_X2 U584 ( .A1(n3871), .A2(n708), .B1(n713), .B2(n429), .ZN(n3081) );
  OAI22_X2 U585 ( .A1(n3870), .A2(n707), .B1(n714), .B2(n428), .ZN(n3082) );
  OAI22_X2 U586 ( .A1(n3869), .A2(n707), .B1(n714), .B2(n427), .ZN(n3083) );
  OAI22_X2 U587 ( .A1(n3868), .A2(n707), .B1(n714), .B2(n426), .ZN(n3084) );
  OAI22_X2 U588 ( .A1(n3867), .A2(n707), .B1(n714), .B2(n425), .ZN(n3085) );
  OAI22_X2 U589 ( .A1(n3866), .A2(n707), .B1(n714), .B2(n424), .ZN(n3086) );
  OAI22_X2 U590 ( .A1(n3865), .A2(n707), .B1(n715), .B2(n423), .ZN(n3087) );
  OAI22_X2 U591 ( .A1(n3864), .A2(n707), .B1(n715), .B2(n422), .ZN(n3088) );
  OAI22_X2 U592 ( .A1(n3863), .A2(n707), .B1(n715), .B2(n421), .ZN(n3089) );
  OAI22_X2 U593 ( .A1(n3862), .A2(n707), .B1(n715), .B2(n420), .ZN(n3090) );
  OAI22_X2 U594 ( .A1(n3861), .A2(n707), .B1(n715), .B2(n419), .ZN(n3091) );
  OAI22_X2 U595 ( .A1(n3860), .A2(n707), .B1(n716), .B2(n418), .ZN(n3092) );
  OAI22_X2 U596 ( .A1(n3859), .A2(n707), .B1(n716), .B2(n417), .ZN(n3093) );
  NAND2_X2 U597 ( .A1(n1352), .A2(n1072), .ZN(n1353) );
  AOI22_X2 U598 ( .A1(DATAIN[0]), .A2(n699), .B1(n700), .B2(\registers[13][0] ), .ZN(n1354) );
  AOI22_X2 U599 ( .A1(DATAIN[1]), .A2(n699), .B1(n700), .B2(\registers[13][1] ), .ZN(n1356) );
  AOI22_X2 U600 ( .A1(DATAIN[2]), .A2(n699), .B1(n700), .B2(\registers[13][2] ), .ZN(n1357) );
  AOI22_X2 U601 ( .A1(DATAIN[3]), .A2(n699), .B1(n700), .B2(\registers[13][3] ), .ZN(n1358) );
  AOI22_X2 U602 ( .A1(DATAIN[4]), .A2(n699), .B1(n700), .B2(\registers[13][4] ), .ZN(n1359) );
  AOI22_X2 U603 ( .A1(DATAIN[5]), .A2(n699), .B1(n701), .B2(\registers[13][5] ), .ZN(n1360) );
  AOI22_X2 U604 ( .A1(DATAIN[6]), .A2(n699), .B1(n701), .B2(\registers[13][6] ), .ZN(n1361) );
  AOI22_X2 U605 ( .A1(DATAIN[7]), .A2(n699), .B1(n701), .B2(\registers[13][7] ), .ZN(n1362) );
  AOI22_X2 U606 ( .A1(DATAIN[8]), .A2(n698), .B1(n701), .B2(\registers[13][8] ), .ZN(n1363) );
  AOI22_X2 U607 ( .A1(DATAIN[9]), .A2(n698), .B1(n701), .B2(\registers[13][9] ), .ZN(n1364) );
  AOI22_X2 U608 ( .A1(DATAIN[10]), .A2(n698), .B1(n702), .B2(
        \registers[13][10] ), .ZN(n1365) );
  AOI22_X2 U609 ( .A1(DATAIN[11]), .A2(n698), .B1(n702), .B2(
        \registers[13][11] ), .ZN(n1366) );
  AOI22_X2 U610 ( .A1(DATAIN[12]), .A2(n698), .B1(n702), .B2(
        \registers[13][12] ), .ZN(n1367) );
  AOI22_X2 U611 ( .A1(DATAIN[13]), .A2(n698), .B1(n702), .B2(
        \registers[13][13] ), .ZN(n1368) );
  AOI22_X2 U612 ( .A1(DATAIN[14]), .A2(n698), .B1(n702), .B2(
        \registers[13][14] ), .ZN(n1369) );
  AOI22_X2 U613 ( .A1(DATAIN[15]), .A2(n698), .B1(n703), .B2(
        \registers[13][15] ), .ZN(n1370) );
  AOI22_X2 U614 ( .A1(DATAIN[16]), .A2(n698), .B1(n703), .B2(
        \registers[13][16] ), .ZN(n1371) );
  AOI22_X2 U615 ( .A1(DATAIN[17]), .A2(n698), .B1(n703), .B2(
        \registers[13][17] ), .ZN(n1372) );
  AOI22_X2 U616 ( .A1(DATAIN[18]), .A2(n698), .B1(n703), .B2(
        \registers[13][18] ), .ZN(n1373) );
  AOI22_X2 U617 ( .A1(DATAIN[19]), .A2(n698), .B1(n703), .B2(
        \registers[13][19] ), .ZN(n1374) );
  AOI22_X2 U618 ( .A1(DATAIN[20]), .A2(n697), .B1(n704), .B2(
        \registers[13][20] ), .ZN(n1375) );
  AOI22_X2 U619 ( .A1(DATAIN[21]), .A2(n697), .B1(n704), .B2(
        \registers[13][21] ), .ZN(n1376) );
  AOI22_X2 U620 ( .A1(DATAIN[22]), .A2(n697), .B1(n704), .B2(
        \registers[13][22] ), .ZN(n1377) );
  AOI22_X2 U621 ( .A1(DATAIN[23]), .A2(n697), .B1(n704), .B2(
        \registers[13][23] ), .ZN(n1378) );
  AOI22_X2 U622 ( .A1(DATAIN[24]), .A2(n697), .B1(n704), .B2(
        \registers[13][24] ), .ZN(n1379) );
  AOI22_X2 U623 ( .A1(DATAIN[25]), .A2(n697), .B1(n705), .B2(
        \registers[13][25] ), .ZN(n1380) );
  AOI22_X2 U624 ( .A1(DATAIN[26]), .A2(n697), .B1(n705), .B2(
        \registers[13][26] ), .ZN(n1381) );
  AOI22_X2 U625 ( .A1(DATAIN[27]), .A2(n697), .B1(n705), .B2(
        \registers[13][27] ), .ZN(n1382) );
  AOI22_X2 U626 ( .A1(DATAIN[28]), .A2(n697), .B1(n705), .B2(
        \registers[13][28] ), .ZN(n1383) );
  AOI22_X2 U627 ( .A1(DATAIN[29]), .A2(n697), .B1(n705), .B2(
        \registers[13][29] ), .ZN(n1384) );
  AOI22_X2 U628 ( .A1(DATAIN[30]), .A2(n697), .B1(n706), .B2(
        \registers[13][30] ), .ZN(n1385) );
  AOI22_X2 U629 ( .A1(DATAIN[31]), .A2(n697), .B1(n706), .B2(
        \registers[13][31] ), .ZN(n1386) );
  NAND2_X2 U630 ( .A1(n1352), .A2(n1106), .ZN(n1355) );
  AOI22_X2 U631 ( .A1(DATAIN[0]), .A2(n689), .B1(n690), .B2(\registers[12][0] ), .ZN(n1387) );
  AOI22_X2 U632 ( .A1(DATAIN[1]), .A2(n689), .B1(n690), .B2(\registers[12][1] ), .ZN(n1389) );
  AOI22_X2 U633 ( .A1(DATAIN[2]), .A2(n689), .B1(n690), .B2(\registers[12][2] ), .ZN(n1390) );
  AOI22_X2 U634 ( .A1(DATAIN[3]), .A2(n689), .B1(n690), .B2(\registers[12][3] ), .ZN(n1391) );
  AOI22_X2 U635 ( .A1(DATAIN[4]), .A2(n689), .B1(n690), .B2(\registers[12][4] ), .ZN(n1392) );
  AOI22_X2 U636 ( .A1(DATAIN[5]), .A2(n689), .B1(n691), .B2(\registers[12][5] ), .ZN(n1393) );
  AOI22_X2 U637 ( .A1(DATAIN[6]), .A2(n689), .B1(n691), .B2(\registers[12][6] ), .ZN(n1394) );
  AOI22_X2 U638 ( .A1(DATAIN[7]), .A2(n689), .B1(n691), .B2(\registers[12][7] ), .ZN(n1395) );
  AOI22_X2 U639 ( .A1(DATAIN[8]), .A2(n688), .B1(n691), .B2(\registers[12][8] ), .ZN(n1396) );
  AOI22_X2 U640 ( .A1(DATAIN[9]), .A2(n688), .B1(n691), .B2(\registers[12][9] ), .ZN(n1397) );
  AOI22_X2 U641 ( .A1(DATAIN[10]), .A2(n688), .B1(n692), .B2(
        \registers[12][10] ), .ZN(n1398) );
  AOI22_X2 U642 ( .A1(DATAIN[11]), .A2(n688), .B1(n692), .B2(
        \registers[12][11] ), .ZN(n1399) );
  AOI22_X2 U643 ( .A1(DATAIN[12]), .A2(n688), .B1(n692), .B2(
        \registers[12][12] ), .ZN(n1400) );
  AOI22_X2 U644 ( .A1(DATAIN[13]), .A2(n688), .B1(n692), .B2(
        \registers[12][13] ), .ZN(n1401) );
  AOI22_X2 U645 ( .A1(DATAIN[14]), .A2(n688), .B1(n692), .B2(
        \registers[12][14] ), .ZN(n1402) );
  AOI22_X2 U646 ( .A1(DATAIN[15]), .A2(n688), .B1(n693), .B2(
        \registers[12][15] ), .ZN(n1403) );
  AOI22_X2 U647 ( .A1(DATAIN[16]), .A2(n688), .B1(n693), .B2(
        \registers[12][16] ), .ZN(n1404) );
  AOI22_X2 U648 ( .A1(DATAIN[17]), .A2(n688), .B1(n693), .B2(
        \registers[12][17] ), .ZN(n1405) );
  AOI22_X2 U649 ( .A1(DATAIN[18]), .A2(n688), .B1(n693), .B2(
        \registers[12][18] ), .ZN(n1406) );
  AOI22_X2 U650 ( .A1(DATAIN[19]), .A2(n688), .B1(n693), .B2(
        \registers[12][19] ), .ZN(n1407) );
  AOI22_X2 U651 ( .A1(DATAIN[20]), .A2(n687), .B1(n694), .B2(
        \registers[12][20] ), .ZN(n1408) );
  AOI22_X2 U652 ( .A1(DATAIN[21]), .A2(n687), .B1(n694), .B2(
        \registers[12][21] ), .ZN(n1409) );
  AOI22_X2 U653 ( .A1(DATAIN[22]), .A2(n687), .B1(n694), .B2(
        \registers[12][22] ), .ZN(n1410) );
  AOI22_X2 U654 ( .A1(DATAIN[23]), .A2(n687), .B1(n694), .B2(
        \registers[12][23] ), .ZN(n1411) );
  AOI22_X2 U655 ( .A1(DATAIN[24]), .A2(n687), .B1(n694), .B2(
        \registers[12][24] ), .ZN(n1412) );
  AOI22_X2 U656 ( .A1(DATAIN[25]), .A2(n687), .B1(n695), .B2(
        \registers[12][25] ), .ZN(n1413) );
  AOI22_X2 U657 ( .A1(DATAIN[26]), .A2(n687), .B1(n695), .B2(
        \registers[12][26] ), .ZN(n1414) );
  AOI22_X2 U658 ( .A1(DATAIN[27]), .A2(n687), .B1(n695), .B2(
        \registers[12][27] ), .ZN(n1415) );
  AOI22_X2 U659 ( .A1(DATAIN[28]), .A2(n687), .B1(n695), .B2(
        \registers[12][28] ), .ZN(n1416) );
  AOI22_X2 U660 ( .A1(DATAIN[29]), .A2(n687), .B1(n695), .B2(
        \registers[12][29] ), .ZN(n1417) );
  AOI22_X2 U661 ( .A1(DATAIN[30]), .A2(n687), .B1(n696), .B2(
        \registers[12][30] ), .ZN(n1418) );
  AOI22_X2 U662 ( .A1(DATAIN[31]), .A2(n687), .B1(n696), .B2(
        \registers[12][31] ), .ZN(n1419) );
  NAND2_X2 U663 ( .A1(n1352), .A2(n1140), .ZN(n1388) );
  OAI22_X2 U664 ( .A1(n3890), .A2(n678), .B1(n679), .B2(n352), .ZN(n3094) );
  OAI22_X2 U665 ( .A1(n3889), .A2(n678), .B1(n679), .B2(n351), .ZN(n3095) );
  OAI22_X2 U666 ( .A1(n3888), .A2(n678), .B1(n679), .B2(n350), .ZN(n3096) );
  OAI22_X2 U667 ( .A1(n3887), .A2(n678), .B1(n679), .B2(n349), .ZN(n3097) );
  OAI22_X2 U668 ( .A1(n3886), .A2(n678), .B1(n679), .B2(n348), .ZN(n3098) );
  OAI22_X2 U669 ( .A1(n3885), .A2(n678), .B1(n680), .B2(n347), .ZN(n3099) );
  OAI22_X2 U670 ( .A1(n3884), .A2(n678), .B1(n680), .B2(n346), .ZN(n3100) );
  OAI22_X2 U671 ( .A1(n3883), .A2(n678), .B1(n680), .B2(n345), .ZN(n3101) );
  OAI22_X2 U672 ( .A1(n3882), .A2(n677), .B1(n680), .B2(n344), .ZN(n3102) );
  OAI22_X2 U673 ( .A1(n3881), .A2(n677), .B1(n680), .B2(n343), .ZN(n3103) );
  OAI22_X2 U674 ( .A1(n3880), .A2(n677), .B1(n681), .B2(n342), .ZN(n3104) );
  OAI22_X2 U675 ( .A1(n3879), .A2(n677), .B1(n681), .B2(n341), .ZN(n3105) );
  OAI22_X2 U676 ( .A1(n3878), .A2(n677), .B1(n681), .B2(n340), .ZN(n3106) );
  OAI22_X2 U677 ( .A1(n3877), .A2(n677), .B1(n681), .B2(n339), .ZN(n3107) );
  OAI22_X2 U678 ( .A1(n3876), .A2(n677), .B1(n681), .B2(n338), .ZN(n3108) );
  OAI22_X2 U679 ( .A1(n3875), .A2(n677), .B1(n682), .B2(n337), .ZN(n3109) );
  OAI22_X2 U680 ( .A1(n3874), .A2(n677), .B1(n682), .B2(n336), .ZN(n3110) );
  OAI22_X2 U681 ( .A1(n3873), .A2(n677), .B1(n682), .B2(n335), .ZN(n3111) );
  OAI22_X2 U682 ( .A1(n3872), .A2(n677), .B1(n682), .B2(n334), .ZN(n3112) );
  OAI22_X2 U683 ( .A1(n3871), .A2(n677), .B1(n682), .B2(n333), .ZN(n3113) );
  OAI22_X2 U684 ( .A1(n3870), .A2(n676), .B1(n683), .B2(n332), .ZN(n3114) );
  OAI22_X2 U685 ( .A1(n3869), .A2(n676), .B1(n683), .B2(n331), .ZN(n3115) );
  OAI22_X2 U686 ( .A1(n3868), .A2(n676), .B1(n683), .B2(n330), .ZN(n3116) );
  OAI22_X2 U687 ( .A1(n3867), .A2(n676), .B1(n683), .B2(n329), .ZN(n3117) );
  OAI22_X2 U688 ( .A1(n3866), .A2(n676), .B1(n683), .B2(n328), .ZN(n3118) );
  OAI22_X2 U689 ( .A1(n3865), .A2(n676), .B1(n684), .B2(n327), .ZN(n3119) );
  OAI22_X2 U690 ( .A1(n3864), .A2(n676), .B1(n684), .B2(n326), .ZN(n3120) );
  OAI22_X2 U691 ( .A1(n3863), .A2(n676), .B1(n684), .B2(n325), .ZN(n3121) );
  OAI22_X2 U692 ( .A1(n3862), .A2(n676), .B1(n684), .B2(n324), .ZN(n3122) );
  OAI22_X2 U693 ( .A1(n3861), .A2(n676), .B1(n684), .B2(n323), .ZN(n3123) );
  OAI22_X2 U694 ( .A1(n3860), .A2(n676), .B1(n685), .B2(n322), .ZN(n3124) );
  OAI22_X2 U695 ( .A1(n3859), .A2(n676), .B1(n685), .B2(n321), .ZN(n3125) );
  NAND2_X2 U696 ( .A1(n1352), .A2(n1142), .ZN(n1420) );
  OAI22_X2 U697 ( .A1(n3890), .A2(n603), .B1(n604), .B2(n320), .ZN(n3126) );
  OAI22_X2 U698 ( .A1(n3889), .A2(n603), .B1(n604), .B2(n319), .ZN(n3127) );
  OAI22_X2 U699 ( .A1(n3888), .A2(n603), .B1(n604), .B2(n318), .ZN(n3128) );
  OAI22_X2 U700 ( .A1(n3887), .A2(n603), .B1(n604), .B2(n317), .ZN(n3129) );
  OAI22_X2 U701 ( .A1(n3886), .A2(n603), .B1(n604), .B2(n316), .ZN(n3130) );
  OAI22_X2 U702 ( .A1(n3885), .A2(n603), .B1(n605), .B2(n315), .ZN(n3131) );
  OAI22_X2 U703 ( .A1(n3884), .A2(n603), .B1(n605), .B2(n314), .ZN(n3132) );
  OAI22_X2 U704 ( .A1(n3883), .A2(n603), .B1(n605), .B2(n313), .ZN(n3133) );
  OAI22_X2 U705 ( .A1(n3882), .A2(n602), .B1(n605), .B2(n312), .ZN(n3134) );
  OAI22_X2 U706 ( .A1(n3881), .A2(n602), .B1(n605), .B2(n311), .ZN(n3135) );
  OAI22_X2 U707 ( .A1(n3880), .A2(n602), .B1(n606), .B2(n310), .ZN(n3136) );
  OAI22_X2 U708 ( .A1(n3879), .A2(n602), .B1(n606), .B2(n309), .ZN(n3137) );
  OAI22_X2 U709 ( .A1(n3878), .A2(n602), .B1(n606), .B2(n308), .ZN(n3138) );
  OAI22_X2 U710 ( .A1(n3877), .A2(n602), .B1(n606), .B2(n307), .ZN(n3139) );
  OAI22_X2 U711 ( .A1(n3876), .A2(n602), .B1(n606), .B2(n306), .ZN(n3140) );
  OAI22_X2 U712 ( .A1(n3875), .A2(n602), .B1(n607), .B2(n305), .ZN(n3141) );
  OAI22_X2 U713 ( .A1(n3874), .A2(n602), .B1(n607), .B2(n304), .ZN(n3142) );
  OAI22_X2 U714 ( .A1(n3873), .A2(n602), .B1(n607), .B2(n303), .ZN(n3143) );
  OAI22_X2 U715 ( .A1(n3872), .A2(n602), .B1(n607), .B2(n302), .ZN(n3144) );
  OAI22_X2 U716 ( .A1(n3871), .A2(n602), .B1(n607), .B2(n301), .ZN(n3145) );
  OAI22_X2 U717 ( .A1(n3870), .A2(n601), .B1(n608), .B2(n300), .ZN(n3146) );
  OAI22_X2 U718 ( .A1(n3869), .A2(n601), .B1(n608), .B2(n299), .ZN(n3147) );
  OAI22_X2 U719 ( .A1(n3868), .A2(n601), .B1(n608), .B2(n298), .ZN(n3148) );
  OAI22_X2 U720 ( .A1(n3867), .A2(n601), .B1(n608), .B2(n297), .ZN(n3149) );
  OAI22_X2 U721 ( .A1(n3866), .A2(n601), .B1(n608), .B2(n296), .ZN(n3150) );
  OAI22_X2 U722 ( .A1(n3865), .A2(n601), .B1(n673), .B2(n295), .ZN(n3151) );
  OAI22_X2 U723 ( .A1(n3864), .A2(n601), .B1(n673), .B2(n294), .ZN(n3152) );
  OAI22_X2 U724 ( .A1(n3863), .A2(n601), .B1(n673), .B2(n293), .ZN(n3153) );
  OAI22_X2 U725 ( .A1(n3862), .A2(n601), .B1(n673), .B2(n292), .ZN(n3154) );
  OAI22_X2 U726 ( .A1(n3861), .A2(n601), .B1(n673), .B2(n291), .ZN(n3155) );
  OAI22_X2 U727 ( .A1(n3860), .A2(n601), .B1(n674), .B2(n290), .ZN(n3156) );
  OAI22_X2 U728 ( .A1(n3859), .A2(n601), .B1(n674), .B2(n289), .ZN(n3157) );
  NAND2_X2 U729 ( .A1(n1352), .A2(n1144), .ZN(n1421) );
  AOI22_X2 U730 ( .A1(DATAIN[0]), .A2(n593), .B1(n594), .B2(\registers[9][0] ), 
        .ZN(n1422) );
  AOI22_X2 U731 ( .A1(DATAIN[1]), .A2(n593), .B1(n594), .B2(\registers[9][1] ), 
        .ZN(n1424) );
  AOI22_X2 U732 ( .A1(DATAIN[2]), .A2(n593), .B1(n594), .B2(\registers[9][2] ), 
        .ZN(n1425) );
  AOI22_X2 U733 ( .A1(DATAIN[3]), .A2(n593), .B1(n594), .B2(\registers[9][3] ), 
        .ZN(n1426) );
  AOI22_X2 U734 ( .A1(DATAIN[4]), .A2(n593), .B1(n594), .B2(\registers[9][4] ), 
        .ZN(n1427) );
  AOI22_X2 U735 ( .A1(DATAIN[5]), .A2(n593), .B1(n595), .B2(\registers[9][5] ), 
        .ZN(n1428) );
  AOI22_X2 U736 ( .A1(DATAIN[6]), .A2(n593), .B1(n595), .B2(\registers[9][6] ), 
        .ZN(n1429) );
  AOI22_X2 U737 ( .A1(DATAIN[7]), .A2(n593), .B1(n595), .B2(\registers[9][7] ), 
        .ZN(n1430) );
  AOI22_X2 U738 ( .A1(DATAIN[8]), .A2(n592), .B1(n595), .B2(\registers[9][8] ), 
        .ZN(n1431) );
  AOI22_X2 U739 ( .A1(DATAIN[9]), .A2(n592), .B1(n595), .B2(\registers[9][9] ), 
        .ZN(n1432) );
  AOI22_X2 U740 ( .A1(DATAIN[10]), .A2(n592), .B1(n596), .B2(
        \registers[9][10] ), .ZN(n1433) );
  AOI22_X2 U741 ( .A1(DATAIN[11]), .A2(n592), .B1(n596), .B2(
        \registers[9][11] ), .ZN(n1434) );
  AOI22_X2 U742 ( .A1(DATAIN[12]), .A2(n592), .B1(n596), .B2(
        \registers[9][12] ), .ZN(n1435) );
  AOI22_X2 U743 ( .A1(DATAIN[13]), .A2(n592), .B1(n596), .B2(
        \registers[9][13] ), .ZN(n1436) );
  AOI22_X2 U744 ( .A1(DATAIN[14]), .A2(n592), .B1(n596), .B2(
        \registers[9][14] ), .ZN(n1437) );
  AOI22_X2 U745 ( .A1(DATAIN[15]), .A2(n592), .B1(n597), .B2(
        \registers[9][15] ), .ZN(n1438) );
  AOI22_X2 U746 ( .A1(DATAIN[16]), .A2(n592), .B1(n597), .B2(
        \registers[9][16] ), .ZN(n1439) );
  AOI22_X2 U747 ( .A1(DATAIN[17]), .A2(n592), .B1(n597), .B2(
        \registers[9][17] ), .ZN(n1440) );
  AOI22_X2 U748 ( .A1(DATAIN[18]), .A2(n592), .B1(n597), .B2(
        \registers[9][18] ), .ZN(n1441) );
  AOI22_X2 U749 ( .A1(DATAIN[19]), .A2(n592), .B1(n597), .B2(
        \registers[9][19] ), .ZN(n1442) );
  AOI22_X2 U750 ( .A1(DATAIN[20]), .A2(n591), .B1(n598), .B2(
        \registers[9][20] ), .ZN(n1443) );
  AOI22_X2 U751 ( .A1(DATAIN[21]), .A2(n591), .B1(n598), .B2(
        \registers[9][21] ), .ZN(n1444) );
  AOI22_X2 U752 ( .A1(DATAIN[22]), .A2(n591), .B1(n598), .B2(
        \registers[9][22] ), .ZN(n1445) );
  AOI22_X2 U753 ( .A1(DATAIN[23]), .A2(n591), .B1(n598), .B2(
        \registers[9][23] ), .ZN(n1446) );
  AOI22_X2 U754 ( .A1(DATAIN[24]), .A2(n591), .B1(n598), .B2(
        \registers[9][24] ), .ZN(n1447) );
  AOI22_X2 U755 ( .A1(DATAIN[25]), .A2(n591), .B1(n599), .B2(
        \registers[9][25] ), .ZN(n1448) );
  AOI22_X2 U756 ( .A1(DATAIN[26]), .A2(n591), .B1(n599), .B2(
        \registers[9][26] ), .ZN(n1449) );
  AOI22_X2 U757 ( .A1(DATAIN[27]), .A2(n591), .B1(n599), .B2(
        \registers[9][27] ), .ZN(n1450) );
  AOI22_X2 U758 ( .A1(DATAIN[28]), .A2(n591), .B1(n599), .B2(
        \registers[9][28] ), .ZN(n1451) );
  AOI22_X2 U759 ( .A1(DATAIN[29]), .A2(n591), .B1(n599), .B2(
        \registers[9][29] ), .ZN(n1452) );
  AOI22_X2 U760 ( .A1(DATAIN[30]), .A2(n591), .B1(n600), .B2(
        \registers[9][30] ), .ZN(n1453) );
  AOI22_X2 U761 ( .A1(DATAIN[31]), .A2(n591), .B1(n600), .B2(
        \registers[9][31] ), .ZN(n1454) );
  NAND2_X2 U762 ( .A1(n1352), .A2(n1178), .ZN(n1423) );
  AOI22_X2 U763 ( .A1(DATAIN[0]), .A2(n583), .B1(n584), .B2(\registers[8][0] ), 
        .ZN(n1455) );
  AOI22_X2 U764 ( .A1(DATAIN[1]), .A2(n583), .B1(n584), .B2(\registers[8][1] ), 
        .ZN(n1457) );
  AOI22_X2 U765 ( .A1(DATAIN[2]), .A2(n583), .B1(n584), .B2(\registers[8][2] ), 
        .ZN(n1458) );
  AOI22_X2 U766 ( .A1(DATAIN[3]), .A2(n583), .B1(n584), .B2(\registers[8][3] ), 
        .ZN(n1459) );
  AOI22_X2 U767 ( .A1(DATAIN[4]), .A2(n583), .B1(n584), .B2(\registers[8][4] ), 
        .ZN(n1460) );
  AOI22_X2 U768 ( .A1(DATAIN[5]), .A2(n583), .B1(n585), .B2(\registers[8][5] ), 
        .ZN(n1461) );
  AOI22_X2 U769 ( .A1(DATAIN[6]), .A2(n583), .B1(n585), .B2(\registers[8][6] ), 
        .ZN(n1462) );
  AOI22_X2 U770 ( .A1(DATAIN[7]), .A2(n583), .B1(n585), .B2(\registers[8][7] ), 
        .ZN(n1463) );
  AOI22_X2 U771 ( .A1(DATAIN[8]), .A2(n582), .B1(n585), .B2(\registers[8][8] ), 
        .ZN(n1464) );
  AOI22_X2 U772 ( .A1(DATAIN[9]), .A2(n582), .B1(n585), .B2(\registers[8][9] ), 
        .ZN(n1465) );
  AOI22_X2 U773 ( .A1(DATAIN[10]), .A2(n582), .B1(n586), .B2(
        \registers[8][10] ), .ZN(n1466) );
  AOI22_X2 U774 ( .A1(DATAIN[11]), .A2(n582), .B1(n586), .B2(
        \registers[8][11] ), .ZN(n1467) );
  AOI22_X2 U775 ( .A1(DATAIN[12]), .A2(n582), .B1(n586), .B2(
        \registers[8][12] ), .ZN(n1468) );
  AOI22_X2 U776 ( .A1(DATAIN[13]), .A2(n582), .B1(n586), .B2(
        \registers[8][13] ), .ZN(n1469) );
  AOI22_X2 U777 ( .A1(DATAIN[14]), .A2(n582), .B1(n586), .B2(
        \registers[8][14] ), .ZN(n1470) );
  AOI22_X2 U778 ( .A1(DATAIN[15]), .A2(n582), .B1(n587), .B2(
        \registers[8][15] ), .ZN(n1471) );
  AOI22_X2 U779 ( .A1(DATAIN[16]), .A2(n582), .B1(n587), .B2(
        \registers[8][16] ), .ZN(n1472) );
  AOI22_X2 U780 ( .A1(DATAIN[17]), .A2(n582), .B1(n587), .B2(
        \registers[8][17] ), .ZN(n1473) );
  AOI22_X2 U781 ( .A1(DATAIN[18]), .A2(n582), .B1(n587), .B2(
        \registers[8][18] ), .ZN(n1474) );
  AOI22_X2 U782 ( .A1(DATAIN[19]), .A2(n582), .B1(n587), .B2(
        \registers[8][19] ), .ZN(n1475) );
  AOI22_X2 U783 ( .A1(DATAIN[20]), .A2(n581), .B1(n588), .B2(
        \registers[8][20] ), .ZN(n1476) );
  AOI22_X2 U784 ( .A1(DATAIN[21]), .A2(n581), .B1(n588), .B2(
        \registers[8][21] ), .ZN(n1477) );
  AOI22_X2 U785 ( .A1(DATAIN[22]), .A2(n581), .B1(n588), .B2(
        \registers[8][22] ), .ZN(n1478) );
  AOI22_X2 U786 ( .A1(DATAIN[23]), .A2(n581), .B1(n588), .B2(
        \registers[8][23] ), .ZN(n1479) );
  AOI22_X2 U787 ( .A1(DATAIN[24]), .A2(n581), .B1(n588), .B2(
        \registers[8][24] ), .ZN(n1480) );
  AOI22_X2 U788 ( .A1(DATAIN[25]), .A2(n581), .B1(n589), .B2(
        \registers[8][25] ), .ZN(n1481) );
  AOI22_X2 U789 ( .A1(DATAIN[26]), .A2(n581), .B1(n589), .B2(
        \registers[8][26] ), .ZN(n1482) );
  AOI22_X2 U790 ( .A1(DATAIN[27]), .A2(n581), .B1(n589), .B2(
        \registers[8][27] ), .ZN(n1483) );
  AOI22_X2 U791 ( .A1(DATAIN[28]), .A2(n581), .B1(n589), .B2(
        \registers[8][28] ), .ZN(n1484) );
  AOI22_X2 U792 ( .A1(DATAIN[29]), .A2(n581), .B1(n589), .B2(
        \registers[8][29] ), .ZN(n1485) );
  AOI22_X2 U793 ( .A1(DATAIN[30]), .A2(n581), .B1(n590), .B2(
        \registers[8][30] ), .ZN(n1486) );
  AOI22_X2 U794 ( .A1(DATAIN[31]), .A2(n581), .B1(n590), .B2(
        \registers[8][31] ), .ZN(n1487) );
  NAND2_X2 U795 ( .A1(n1352), .A2(n1212), .ZN(n1456) );
  AND3_X2 U796 ( .A1(n1213), .A2(n3592), .A3(ADD_WR[3]), .ZN(n1352) );
  AOI22_X2 U797 ( .A1(DATAIN[0]), .A2(n573), .B1(n574), .B2(\registers[7][0] ), 
        .ZN(n1488) );
  AOI22_X2 U798 ( .A1(DATAIN[1]), .A2(n573), .B1(n574), .B2(\registers[7][1] ), 
        .ZN(n1490) );
  AOI22_X2 U799 ( .A1(DATAIN[2]), .A2(n573), .B1(n574), .B2(\registers[7][2] ), 
        .ZN(n1491) );
  AOI22_X2 U800 ( .A1(DATAIN[3]), .A2(n573), .B1(n574), .B2(\registers[7][3] ), 
        .ZN(n1492) );
  AOI22_X2 U801 ( .A1(DATAIN[4]), .A2(n573), .B1(n574), .B2(\registers[7][4] ), 
        .ZN(n1493) );
  AOI22_X2 U802 ( .A1(DATAIN[5]), .A2(n573), .B1(n575), .B2(\registers[7][5] ), 
        .ZN(n1494) );
  AOI22_X2 U803 ( .A1(DATAIN[6]), .A2(n573), .B1(n575), .B2(\registers[7][6] ), 
        .ZN(n1495) );
  AOI22_X2 U804 ( .A1(DATAIN[7]), .A2(n573), .B1(n575), .B2(\registers[7][7] ), 
        .ZN(n1496) );
  AOI22_X2 U805 ( .A1(DATAIN[8]), .A2(n572), .B1(n575), .B2(\registers[7][8] ), 
        .ZN(n1497) );
  AOI22_X2 U806 ( .A1(DATAIN[9]), .A2(n572), .B1(n575), .B2(\registers[7][9] ), 
        .ZN(n1498) );
  AOI22_X2 U807 ( .A1(DATAIN[10]), .A2(n572), .B1(n576), .B2(
        \registers[7][10] ), .ZN(n1499) );
  AOI22_X2 U808 ( .A1(DATAIN[11]), .A2(n572), .B1(n576), .B2(
        \registers[7][11] ), .ZN(n1500) );
  AOI22_X2 U809 ( .A1(DATAIN[12]), .A2(n572), .B1(n576), .B2(
        \registers[7][12] ), .ZN(n1501) );
  AOI22_X2 U810 ( .A1(DATAIN[13]), .A2(n572), .B1(n576), .B2(
        \registers[7][13] ), .ZN(n1502) );
  AOI22_X2 U811 ( .A1(DATAIN[14]), .A2(n572), .B1(n576), .B2(
        \registers[7][14] ), .ZN(n1503) );
  AOI22_X2 U812 ( .A1(DATAIN[15]), .A2(n572), .B1(n577), .B2(
        \registers[7][15] ), .ZN(n1504) );
  AOI22_X2 U813 ( .A1(DATAIN[16]), .A2(n572), .B1(n577), .B2(
        \registers[7][16] ), .ZN(n1505) );
  AOI22_X2 U814 ( .A1(DATAIN[17]), .A2(n572), .B1(n577), .B2(
        \registers[7][17] ), .ZN(n1506) );
  AOI22_X2 U815 ( .A1(DATAIN[18]), .A2(n572), .B1(n577), .B2(
        \registers[7][18] ), .ZN(n1507) );
  AOI22_X2 U816 ( .A1(DATAIN[19]), .A2(n572), .B1(n577), .B2(
        \registers[7][19] ), .ZN(n1508) );
  AOI22_X2 U817 ( .A1(DATAIN[20]), .A2(n571), .B1(n578), .B2(
        \registers[7][20] ), .ZN(n1509) );
  AOI22_X2 U818 ( .A1(DATAIN[21]), .A2(n571), .B1(n578), .B2(
        \registers[7][21] ), .ZN(n1510) );
  AOI22_X2 U819 ( .A1(DATAIN[22]), .A2(n571), .B1(n578), .B2(
        \registers[7][22] ), .ZN(n1511) );
  AOI22_X2 U820 ( .A1(DATAIN[23]), .A2(n571), .B1(n578), .B2(
        \registers[7][23] ), .ZN(n1512) );
  AOI22_X2 U821 ( .A1(DATAIN[24]), .A2(n571), .B1(n578), .B2(
        \registers[7][24] ), .ZN(n1513) );
  AOI22_X2 U822 ( .A1(DATAIN[25]), .A2(n571), .B1(n579), .B2(
        \registers[7][25] ), .ZN(n1514) );
  AOI22_X2 U823 ( .A1(DATAIN[26]), .A2(n571), .B1(n579), .B2(
        \registers[7][26] ), .ZN(n1515) );
  AOI22_X2 U824 ( .A1(DATAIN[27]), .A2(n571), .B1(n579), .B2(
        \registers[7][27] ), .ZN(n1516) );
  AOI22_X2 U825 ( .A1(DATAIN[28]), .A2(n571), .B1(n579), .B2(
        \registers[7][28] ), .ZN(n1517) );
  AOI22_X2 U826 ( .A1(DATAIN[29]), .A2(n571), .B1(n579), .B2(
        \registers[7][29] ), .ZN(n1518) );
  AOI22_X2 U827 ( .A1(DATAIN[30]), .A2(n571), .B1(n580), .B2(
        \registers[7][30] ), .ZN(n1519) );
  AOI22_X2 U828 ( .A1(DATAIN[31]), .A2(n571), .B1(n580), .B2(
        \registers[7][31] ), .ZN(n1520) );
  NAND2_X2 U829 ( .A1(n1521), .A2(n1069), .ZN(n1489) );
  NOR3_X2 U830 ( .A1(n3851), .A2(n3852), .A3(n3850), .ZN(n1069) );
  AOI22_X2 U831 ( .A1(DATAIN[0]), .A2(n563), .B1(n564), .B2(\registers[6][0] ), 
        .ZN(n1522) );
  AOI22_X2 U832 ( .A1(DATAIN[1]), .A2(n563), .B1(n564), .B2(\registers[6][1] ), 
        .ZN(n1524) );
  AOI22_X2 U833 ( .A1(DATAIN[2]), .A2(n563), .B1(n564), .B2(\registers[6][2] ), 
        .ZN(n1525) );
  AOI22_X2 U834 ( .A1(DATAIN[3]), .A2(n563), .B1(n564), .B2(\registers[6][3] ), 
        .ZN(n1526) );
  AOI22_X2 U835 ( .A1(DATAIN[4]), .A2(n563), .B1(n564), .B2(\registers[6][4] ), 
        .ZN(n1527) );
  AOI22_X2 U836 ( .A1(DATAIN[5]), .A2(n563), .B1(n565), .B2(\registers[6][5] ), 
        .ZN(n1528) );
  AOI22_X2 U837 ( .A1(DATAIN[6]), .A2(n563), .B1(n565), .B2(\registers[6][6] ), 
        .ZN(n1529) );
  AOI22_X2 U838 ( .A1(DATAIN[7]), .A2(n563), .B1(n565), .B2(\registers[6][7] ), 
        .ZN(n1530) );
  AOI22_X2 U839 ( .A1(DATAIN[8]), .A2(n562), .B1(n565), .B2(\registers[6][8] ), 
        .ZN(n1531) );
  AOI22_X2 U840 ( .A1(DATAIN[9]), .A2(n562), .B1(n565), .B2(\registers[6][9] ), 
        .ZN(n1532) );
  AOI22_X2 U841 ( .A1(DATAIN[10]), .A2(n562), .B1(n566), .B2(
        \registers[6][10] ), .ZN(n1533) );
  AOI22_X2 U842 ( .A1(DATAIN[11]), .A2(n562), .B1(n566), .B2(
        \registers[6][11] ), .ZN(n1534) );
  AOI22_X2 U843 ( .A1(DATAIN[12]), .A2(n562), .B1(n566), .B2(
        \registers[6][12] ), .ZN(n1535) );
  AOI22_X2 U844 ( .A1(DATAIN[13]), .A2(n562), .B1(n566), .B2(
        \registers[6][13] ), .ZN(n1536) );
  AOI22_X2 U845 ( .A1(DATAIN[14]), .A2(n562), .B1(n566), .B2(
        \registers[6][14] ), .ZN(n1537) );
  AOI22_X2 U846 ( .A1(DATAIN[15]), .A2(n562), .B1(n567), .B2(
        \registers[6][15] ), .ZN(n1538) );
  AOI22_X2 U847 ( .A1(DATAIN[16]), .A2(n562), .B1(n567), .B2(
        \registers[6][16] ), .ZN(n1539) );
  AOI22_X2 U848 ( .A1(DATAIN[17]), .A2(n562), .B1(n567), .B2(
        \registers[6][17] ), .ZN(n1540) );
  AOI22_X2 U849 ( .A1(DATAIN[18]), .A2(n562), .B1(n567), .B2(
        \registers[6][18] ), .ZN(n1541) );
  AOI22_X2 U850 ( .A1(DATAIN[19]), .A2(n562), .B1(n567), .B2(
        \registers[6][19] ), .ZN(n1542) );
  AOI22_X2 U851 ( .A1(DATAIN[20]), .A2(n561), .B1(n568), .B2(
        \registers[6][20] ), .ZN(n1543) );
  AOI22_X2 U852 ( .A1(DATAIN[21]), .A2(n561), .B1(n568), .B2(
        \registers[6][21] ), .ZN(n1544) );
  AOI22_X2 U853 ( .A1(DATAIN[22]), .A2(n561), .B1(n568), .B2(
        \registers[6][22] ), .ZN(n1545) );
  AOI22_X2 U854 ( .A1(DATAIN[23]), .A2(n561), .B1(n568), .B2(
        \registers[6][23] ), .ZN(n1546) );
  AOI22_X2 U855 ( .A1(DATAIN[24]), .A2(n561), .B1(n568), .B2(
        \registers[6][24] ), .ZN(n1547) );
  AOI22_X2 U856 ( .A1(DATAIN[25]), .A2(n561), .B1(n569), .B2(
        \registers[6][25] ), .ZN(n1548) );
  AOI22_X2 U857 ( .A1(DATAIN[26]), .A2(n561), .B1(n569), .B2(
        \registers[6][26] ), .ZN(n1549) );
  AOI22_X2 U858 ( .A1(DATAIN[27]), .A2(n561), .B1(n569), .B2(
        \registers[6][27] ), .ZN(n1550) );
  AOI22_X2 U859 ( .A1(DATAIN[28]), .A2(n561), .B1(n569), .B2(
        \registers[6][28] ), .ZN(n1551) );
  AOI22_X2 U860 ( .A1(DATAIN[29]), .A2(n561), .B1(n569), .B2(
        \registers[6][29] ), .ZN(n1552) );
  AOI22_X2 U861 ( .A1(DATAIN[30]), .A2(n561), .B1(n570), .B2(
        \registers[6][30] ), .ZN(n1553) );
  AOI22_X2 U862 ( .A1(DATAIN[31]), .A2(n561), .B1(n570), .B2(
        \registers[6][31] ), .ZN(n1554) );
  NAND2_X2 U863 ( .A1(n1521), .A2(n1072), .ZN(n1523) );
  NOR3_X2 U864 ( .A1(n3851), .A2(ADD_WR[0]), .A3(n3850), .ZN(n1072) );
  OAI22_X2 U865 ( .A1(n3890), .A2(n552), .B1(n553), .B2(n160), .ZN(n3158) );
  OAI22_X2 U866 ( .A1(n3889), .A2(n552), .B1(n553), .B2(n159), .ZN(n3159) );
  OAI22_X2 U867 ( .A1(n3888), .A2(n552), .B1(n553), .B2(n158), .ZN(n3160) );
  OAI22_X2 U868 ( .A1(n3887), .A2(n552), .B1(n553), .B2(n157), .ZN(n3161) );
  OAI22_X2 U869 ( .A1(n3886), .A2(n552), .B1(n553), .B2(n156), .ZN(n3162) );
  OAI22_X2 U870 ( .A1(n3885), .A2(n552), .B1(n554), .B2(n155), .ZN(n3163) );
  OAI22_X2 U871 ( .A1(n3884), .A2(n552), .B1(n554), .B2(n154), .ZN(n3164) );
  OAI22_X2 U872 ( .A1(n3883), .A2(n552), .B1(n554), .B2(n153), .ZN(n3165) );
  OAI22_X2 U873 ( .A1(n3882), .A2(n551), .B1(n554), .B2(n152), .ZN(n3166) );
  OAI22_X2 U874 ( .A1(n3881), .A2(n551), .B1(n554), .B2(n151), .ZN(n3167) );
  OAI22_X2 U875 ( .A1(n3880), .A2(n551), .B1(n555), .B2(n150), .ZN(n3168) );
  OAI22_X2 U876 ( .A1(n3879), .A2(n551), .B1(n555), .B2(n149), .ZN(n3169) );
  OAI22_X2 U877 ( .A1(n3878), .A2(n551), .B1(n555), .B2(n148), .ZN(n3170) );
  OAI22_X2 U878 ( .A1(n3877), .A2(n551), .B1(n555), .B2(n147), .ZN(n3171) );
  OAI22_X2 U879 ( .A1(n3876), .A2(n551), .B1(n555), .B2(n146), .ZN(n3172) );
  OAI22_X2 U880 ( .A1(n3875), .A2(n551), .B1(n556), .B2(n145), .ZN(n3173) );
  OAI22_X2 U881 ( .A1(n3874), .A2(n551), .B1(n556), .B2(n144), .ZN(n3174) );
  OAI22_X2 U882 ( .A1(n3873), .A2(n551), .B1(n556), .B2(n143), .ZN(n3175) );
  OAI22_X2 U883 ( .A1(n3872), .A2(n551), .B1(n556), .B2(n142), .ZN(n3176) );
  OAI22_X2 U884 ( .A1(n3871), .A2(n551), .B1(n556), .B2(n141), .ZN(n3177) );
  OAI22_X2 U885 ( .A1(n3870), .A2(n550), .B1(n557), .B2(n140), .ZN(n3178) );
  OAI22_X2 U886 ( .A1(n3869), .A2(n550), .B1(n557), .B2(n139), .ZN(n3179) );
  OAI22_X2 U887 ( .A1(n3868), .A2(n550), .B1(n557), .B2(n138), .ZN(n3180) );
  OAI22_X2 U888 ( .A1(n3867), .A2(n550), .B1(n557), .B2(n137), .ZN(n3181) );
  OAI22_X2 U889 ( .A1(n3866), .A2(n550), .B1(n557), .B2(n136), .ZN(n3182) );
  OAI22_X2 U890 ( .A1(n3865), .A2(n550), .B1(n558), .B2(n135), .ZN(n3183) );
  OAI22_X2 U891 ( .A1(n3864), .A2(n550), .B1(n558), .B2(n134), .ZN(n3184) );
  OAI22_X2 U892 ( .A1(n3863), .A2(n550), .B1(n558), .B2(n133), .ZN(n3185) );
  OAI22_X2 U893 ( .A1(n3862), .A2(n550), .B1(n558), .B2(n132), .ZN(n3186) );
  OAI22_X2 U894 ( .A1(n3861), .A2(n550), .B1(n558), .B2(n131), .ZN(n3187) );
  OAI22_X2 U895 ( .A1(n3860), .A2(n550), .B1(n559), .B2(n130), .ZN(n3188) );
  OAI22_X2 U896 ( .A1(n3859), .A2(n550), .B1(n559), .B2(n129), .ZN(n3189) );
  NAND2_X2 U897 ( .A1(n1521), .A2(n1106), .ZN(n1555) );
  NOR3_X2 U898 ( .A1(n3852), .A2(ADD_WR[1]), .A3(n3850), .ZN(n1106) );
  OAI22_X2 U899 ( .A1(n3890), .A2(n413), .B1(n414), .B2(n128), .ZN(n3190) );
  OAI22_X2 U900 ( .A1(n3889), .A2(n413), .B1(n414), .B2(n127), .ZN(n3191) );
  OAI22_X2 U901 ( .A1(n3888), .A2(n413), .B1(n414), .B2(n126), .ZN(n3192) );
  OAI22_X2 U902 ( .A1(n3887), .A2(n413), .B1(n414), .B2(n125), .ZN(n3193) );
  OAI22_X2 U903 ( .A1(n3886), .A2(n413), .B1(n414), .B2(n124), .ZN(n3194) );
  OAI22_X2 U904 ( .A1(n3885), .A2(n413), .B1(n415), .B2(n123), .ZN(n3195) );
  OAI22_X2 U905 ( .A1(n3884), .A2(n413), .B1(n415), .B2(n122), .ZN(n3196) );
  OAI22_X2 U906 ( .A1(n3883), .A2(n413), .B1(n415), .B2(n121), .ZN(n3197) );
  OAI22_X2 U907 ( .A1(n3882), .A2(n412), .B1(n415), .B2(n120), .ZN(n3198) );
  OAI22_X2 U908 ( .A1(n3881), .A2(n412), .B1(n415), .B2(n119), .ZN(n3199) );
  OAI22_X2 U909 ( .A1(n3880), .A2(n412), .B1(n416), .B2(n118), .ZN(n3200) );
  OAI22_X2 U910 ( .A1(n3879), .A2(n412), .B1(n416), .B2(n117), .ZN(n3201) );
  OAI22_X2 U911 ( .A1(n3878), .A2(n412), .B1(n416), .B2(n116), .ZN(n3202) );
  OAI22_X2 U912 ( .A1(n3877), .A2(n412), .B1(n416), .B2(n115), .ZN(n3203) );
  OAI22_X2 U913 ( .A1(n3876), .A2(n412), .B1(n416), .B2(n114), .ZN(n3204) );
  OAI22_X2 U914 ( .A1(n3875), .A2(n412), .B1(n545), .B2(n113), .ZN(n3205) );
  OAI22_X2 U915 ( .A1(n3874), .A2(n412), .B1(n545), .B2(n112), .ZN(n3206) );
  OAI22_X2 U916 ( .A1(n3873), .A2(n412), .B1(n545), .B2(n111), .ZN(n3207) );
  OAI22_X2 U917 ( .A1(n3872), .A2(n412), .B1(n545), .B2(n110), .ZN(n3208) );
  OAI22_X2 U918 ( .A1(n3871), .A2(n412), .B1(n545), .B2(n109), .ZN(n3209) );
  OAI22_X2 U919 ( .A1(n3870), .A2(n411), .B1(n546), .B2(n108), .ZN(n3210) );
  OAI22_X2 U920 ( .A1(n3869), .A2(n411), .B1(n546), .B2(n107), .ZN(n3211) );
  OAI22_X2 U921 ( .A1(n3868), .A2(n411), .B1(n546), .B2(n106), .ZN(n3212) );
  OAI22_X2 U922 ( .A1(n3867), .A2(n411), .B1(n546), .B2(n105), .ZN(n3213) );
  OAI22_X2 U923 ( .A1(n3866), .A2(n411), .B1(n546), .B2(n104), .ZN(n3214) );
  OAI22_X2 U924 ( .A1(n3865), .A2(n411), .B1(n547), .B2(n103), .ZN(n3215) );
  OAI22_X2 U925 ( .A1(n3864), .A2(n411), .B1(n547), .B2(n102), .ZN(n3216) );
  OAI22_X2 U926 ( .A1(n3863), .A2(n411), .B1(n547), .B2(n101), .ZN(n3217) );
  OAI22_X2 U927 ( .A1(n3862), .A2(n411), .B1(n547), .B2(n100), .ZN(n3218) );
  OAI22_X2 U928 ( .A1(n3861), .A2(n411), .B1(n547), .B2(n99), .ZN(n3219) );
  OAI22_X2 U929 ( .A1(n3860), .A2(n411), .B1(n548), .B2(n98), .ZN(n3220) );
  OAI22_X2 U930 ( .A1(n3859), .A2(n411), .B1(n548), .B2(n97), .ZN(n3221) );
  NAND2_X2 U931 ( .A1(n1521), .A2(n1140), .ZN(n1556) );
  NOR3_X2 U932 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n3850), .ZN(n1140) );
  OAI22_X2 U933 ( .A1(n3890), .A2(n402), .B1(n403), .B2(n96), .ZN(n3222) );
  OAI22_X2 U934 ( .A1(n3889), .A2(n402), .B1(n403), .B2(n95), .ZN(n3223) );
  OAI22_X2 U935 ( .A1(n3888), .A2(n402), .B1(n403), .B2(n94), .ZN(n3224) );
  OAI22_X2 U936 ( .A1(n3887), .A2(n402), .B1(n403), .B2(n93), .ZN(n3225) );
  OAI22_X2 U937 ( .A1(n3886), .A2(n402), .B1(n403), .B2(n92), .ZN(n3226) );
  OAI22_X2 U938 ( .A1(n3885), .A2(n402), .B1(n404), .B2(n91), .ZN(n3227) );
  OAI22_X2 U939 ( .A1(n3884), .A2(n402), .B1(n404), .B2(n90), .ZN(n3228) );
  OAI22_X2 U940 ( .A1(n3883), .A2(n402), .B1(n404), .B2(n89), .ZN(n3229) );
  OAI22_X2 U941 ( .A1(n3882), .A2(n401), .B1(n404), .B2(n88), .ZN(n3230) );
  OAI22_X2 U942 ( .A1(n3881), .A2(n401), .B1(n404), .B2(n87), .ZN(n3231) );
  OAI22_X2 U943 ( .A1(n3880), .A2(n401), .B1(n405), .B2(n86), .ZN(n3232) );
  OAI22_X2 U944 ( .A1(n3879), .A2(n401), .B1(n405), .B2(n85), .ZN(n3233) );
  OAI22_X2 U945 ( .A1(n3878), .A2(n401), .B1(n405), .B2(n84), .ZN(n3234) );
  OAI22_X2 U946 ( .A1(n3877), .A2(n401), .B1(n405), .B2(n83), .ZN(n3235) );
  OAI22_X2 U947 ( .A1(n3876), .A2(n401), .B1(n405), .B2(n82), .ZN(n3236) );
  OAI22_X2 U948 ( .A1(n3875), .A2(n401), .B1(n406), .B2(n81), .ZN(n3237) );
  OAI22_X2 U949 ( .A1(n3874), .A2(n401), .B1(n406), .B2(n80), .ZN(n3238) );
  OAI22_X2 U950 ( .A1(n3873), .A2(n401), .B1(n406), .B2(n79), .ZN(n3239) );
  OAI22_X2 U951 ( .A1(n3872), .A2(n401), .B1(n406), .B2(n78), .ZN(n3240) );
  OAI22_X2 U952 ( .A1(n3871), .A2(n401), .B1(n406), .B2(n77), .ZN(n3241) );
  OAI22_X2 U953 ( .A1(n3870), .A2(n400), .B1(n407), .B2(n76), .ZN(n3242) );
  OAI22_X2 U954 ( .A1(n3869), .A2(n400), .B1(n407), .B2(n75), .ZN(n3243) );
  OAI22_X2 U955 ( .A1(n3868), .A2(n400), .B1(n407), .B2(n74), .ZN(n3244) );
  OAI22_X2 U956 ( .A1(n3867), .A2(n400), .B1(n407), .B2(n73), .ZN(n3245) );
  OAI22_X2 U957 ( .A1(n3866), .A2(n400), .B1(n407), .B2(n72), .ZN(n3246) );
  OAI22_X2 U958 ( .A1(n3865), .A2(n400), .B1(n408), .B2(n71), .ZN(n3247) );
  OAI22_X2 U959 ( .A1(n3864), .A2(n400), .B1(n408), .B2(n70), .ZN(n3248) );
  OAI22_X2 U960 ( .A1(n3863), .A2(n400), .B1(n408), .B2(n69), .ZN(n3249) );
  OAI22_X2 U961 ( .A1(n3862), .A2(n400), .B1(n408), .B2(n68), .ZN(n3250) );
  OAI22_X2 U962 ( .A1(n3861), .A2(n400), .B1(n408), .B2(n67), .ZN(n3251) );
  OAI22_X2 U963 ( .A1(n3860), .A2(n400), .B1(n409), .B2(n66), .ZN(n3252) );
  OAI22_X2 U964 ( .A1(n3859), .A2(n400), .B1(n409), .B2(n65), .ZN(n3253) );
  NAND2_X2 U965 ( .A1(n1521), .A2(n1142), .ZN(n1557) );
  NOR3_X2 U966 ( .A1(n3852), .A2(ADD_WR[2]), .A3(n3851), .ZN(n1142) );
  OAI22_X2 U967 ( .A1(n3890), .A2(n391), .B1(n392), .B2(n64), .ZN(n3254) );
  OAI22_X2 U968 ( .A1(n3889), .A2(n391), .B1(n392), .B2(n63), .ZN(n3255) );
  OAI22_X2 U969 ( .A1(n3888), .A2(n391), .B1(n392), .B2(n62), .ZN(n3256) );
  OAI22_X2 U970 ( .A1(n3887), .A2(n391), .B1(n392), .B2(n61), .ZN(n3257) );
  OAI22_X2 U971 ( .A1(n3886), .A2(n391), .B1(n392), .B2(n60), .ZN(n3258) );
  OAI22_X2 U972 ( .A1(n3885), .A2(n391), .B1(n393), .B2(n59), .ZN(n3259) );
  OAI22_X2 U973 ( .A1(n3884), .A2(n391), .B1(n393), .B2(n58), .ZN(n3260) );
  OAI22_X2 U974 ( .A1(n3883), .A2(n391), .B1(n393), .B2(n57), .ZN(n3261) );
  OAI22_X2 U975 ( .A1(n3882), .A2(n390), .B1(n393), .B2(n56), .ZN(n3262) );
  OAI22_X2 U976 ( .A1(n3881), .A2(n390), .B1(n393), .B2(n55), .ZN(n3263) );
  OAI22_X2 U977 ( .A1(n3880), .A2(n390), .B1(n394), .B2(n54), .ZN(n3264) );
  OAI22_X2 U978 ( .A1(n3879), .A2(n390), .B1(n394), .B2(n53), .ZN(n3265) );
  OAI22_X2 U979 ( .A1(n3878), .A2(n390), .B1(n394), .B2(n52), .ZN(n3266) );
  OAI22_X2 U980 ( .A1(n3877), .A2(n390), .B1(n394), .B2(n51), .ZN(n3267) );
  OAI22_X2 U981 ( .A1(n3876), .A2(n390), .B1(n394), .B2(n50), .ZN(n3268) );
  OAI22_X2 U982 ( .A1(n3875), .A2(n390), .B1(n395), .B2(n49), .ZN(n3269) );
  OAI22_X2 U983 ( .A1(n3874), .A2(n390), .B1(n395), .B2(n48), .ZN(n3270) );
  OAI22_X2 U984 ( .A1(n3873), .A2(n390), .B1(n395), .B2(n47), .ZN(n3271) );
  OAI22_X2 U985 ( .A1(n3872), .A2(n390), .B1(n395), .B2(n46), .ZN(n3272) );
  OAI22_X2 U986 ( .A1(n3871), .A2(n390), .B1(n395), .B2(n45), .ZN(n3273) );
  OAI22_X2 U987 ( .A1(n3870), .A2(n389), .B1(n396), .B2(n44), .ZN(n3274) );
  OAI22_X2 U988 ( .A1(n3869), .A2(n389), .B1(n396), .B2(n43), .ZN(n3275) );
  OAI22_X2 U989 ( .A1(n3868), .A2(n389), .B1(n396), .B2(n42), .ZN(n3276) );
  OAI22_X2 U990 ( .A1(n3867), .A2(n389), .B1(n396), .B2(n41), .ZN(n3277) );
  OAI22_X2 U991 ( .A1(n3866), .A2(n389), .B1(n396), .B2(n40), .ZN(n3278) );
  OAI22_X2 U992 ( .A1(n3865), .A2(n389), .B1(n397), .B2(n39), .ZN(n3279) );
  OAI22_X2 U993 ( .A1(n3864), .A2(n389), .B1(n397), .B2(n38), .ZN(n3280) );
  OAI22_X2 U994 ( .A1(n3863), .A2(n389), .B1(n397), .B2(n37), .ZN(n3281) );
  OAI22_X2 U995 ( .A1(n3862), .A2(n389), .B1(n397), .B2(n36), .ZN(n3282) );
  OAI22_X2 U996 ( .A1(n3861), .A2(n389), .B1(n397), .B2(n35), .ZN(n3283) );
  OAI22_X2 U997 ( .A1(n3860), .A2(n389), .B1(n398), .B2(n34), .ZN(n3284) );
  OAI22_X2 U998 ( .A1(n3859), .A2(n389), .B1(n398), .B2(n33), .ZN(n3285) );
  NAND2_X2 U999 ( .A1(n1521), .A2(n1144), .ZN(n1558) );
  NOR3_X2 U1000 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n3851), .ZN(n1144) );
  AOI22_X2 U1001 ( .A1(DATAIN[0]), .A2(n381), .B1(n382), .B2(\registers[1][0] ), .ZN(n1559) );
  AOI22_X2 U1002 ( .A1(DATAIN[1]), .A2(n381), .B1(n382), .B2(\registers[1][1] ), .ZN(n1561) );
  AOI22_X2 U1003 ( .A1(DATAIN[2]), .A2(n381), .B1(n382), .B2(\registers[1][2] ), .ZN(n1562) );
  AOI22_X2 U1004 ( .A1(DATAIN[3]), .A2(n381), .B1(n382), .B2(\registers[1][3] ), .ZN(n1563) );
  AOI22_X2 U1005 ( .A1(DATAIN[4]), .A2(n381), .B1(n382), .B2(\registers[1][4] ), .ZN(n1564) );
  AOI22_X2 U1006 ( .A1(DATAIN[5]), .A2(n381), .B1(n383), .B2(\registers[1][5] ), .ZN(n1565) );
  AOI22_X2 U1007 ( .A1(DATAIN[6]), .A2(n381), .B1(n383), .B2(\registers[1][6] ), .ZN(n1566) );
  AOI22_X2 U1008 ( .A1(DATAIN[7]), .A2(n381), .B1(n383), .B2(\registers[1][7] ), .ZN(n1567) );
  AOI22_X2 U1009 ( .A1(DATAIN[8]), .A2(n380), .B1(n383), .B2(\registers[1][8] ), .ZN(n1568) );
  AOI22_X2 U1010 ( .A1(DATAIN[9]), .A2(n380), .B1(n383), .B2(\registers[1][9] ), .ZN(n1569) );
  AOI22_X2 U1011 ( .A1(DATAIN[10]), .A2(n380), .B1(n384), .B2(
        \registers[1][10] ), .ZN(n1570) );
  AOI22_X2 U1012 ( .A1(DATAIN[11]), .A2(n380), .B1(n384), .B2(
        \registers[1][11] ), .ZN(n1571) );
  AOI22_X2 U1013 ( .A1(DATAIN[12]), .A2(n380), .B1(n384), .B2(
        \registers[1][12] ), .ZN(n1572) );
  AOI22_X2 U1014 ( .A1(DATAIN[13]), .A2(n380), .B1(n384), .B2(
        \registers[1][13] ), .ZN(n1573) );
  AOI22_X2 U1015 ( .A1(DATAIN[14]), .A2(n380), .B1(n384), .B2(
        \registers[1][14] ), .ZN(n1574) );
  AOI22_X2 U1016 ( .A1(DATAIN[15]), .A2(n380), .B1(n385), .B2(
        \registers[1][15] ), .ZN(n1575) );
  AOI22_X2 U1017 ( .A1(DATAIN[16]), .A2(n380), .B1(n385), .B2(
        \registers[1][16] ), .ZN(n1576) );
  AOI22_X2 U1018 ( .A1(DATAIN[17]), .A2(n380), .B1(n385), .B2(
        \registers[1][17] ), .ZN(n1577) );
  AOI22_X2 U1019 ( .A1(DATAIN[18]), .A2(n380), .B1(n385), .B2(
        \registers[1][18] ), .ZN(n1578) );
  AOI22_X2 U1020 ( .A1(DATAIN[19]), .A2(n380), .B1(n385), .B2(
        \registers[1][19] ), .ZN(n1579) );
  AOI22_X2 U1021 ( .A1(DATAIN[20]), .A2(n379), .B1(n386), .B2(
        \registers[1][20] ), .ZN(n1580) );
  AOI22_X2 U1022 ( .A1(DATAIN[21]), .A2(n379), .B1(n386), .B2(
        \registers[1][21] ), .ZN(n1581) );
  AOI22_X2 U1023 ( .A1(DATAIN[22]), .A2(n379), .B1(n386), .B2(
        \registers[1][22] ), .ZN(n1582) );
  AOI22_X2 U1024 ( .A1(DATAIN[23]), .A2(n379), .B1(n386), .B2(
        \registers[1][23] ), .ZN(n1583) );
  AOI22_X2 U1025 ( .A1(DATAIN[24]), .A2(n379), .B1(n386), .B2(
        \registers[1][24] ), .ZN(n1584) );
  AOI22_X2 U1026 ( .A1(DATAIN[25]), .A2(n379), .B1(n387), .B2(
        \registers[1][25] ), .ZN(n1585) );
  AOI22_X2 U1027 ( .A1(DATAIN[26]), .A2(n379), .B1(n387), .B2(
        \registers[1][26] ), .ZN(n1586) );
  AOI22_X2 U1028 ( .A1(DATAIN[27]), .A2(n379), .B1(n387), .B2(
        \registers[1][27] ), .ZN(n1587) );
  AOI22_X2 U1029 ( .A1(DATAIN[28]), .A2(n379), .B1(n387), .B2(
        \registers[1][28] ), .ZN(n1588) );
  AOI22_X2 U1030 ( .A1(DATAIN[29]), .A2(n379), .B1(n387), .B2(
        \registers[1][29] ), .ZN(n1589) );
  AOI22_X2 U1031 ( .A1(DATAIN[30]), .A2(n379), .B1(n388), .B2(
        \registers[1][30] ), .ZN(n1590) );
  AOI22_X2 U1032 ( .A1(DATAIN[31]), .A2(n379), .B1(n388), .B2(
        \registers[1][31] ), .ZN(n1591) );
  NAND2_X2 U1033 ( .A1(n1521), .A2(n1178), .ZN(n1560) );
  NOR3_X2 U1034 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n3852), .ZN(n1178) );
  NOR3_X2 U1035 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n1212)
         );
  AND3_X2 U1036 ( .A1(n3849), .A2(n3592), .A3(n1213), .ZN(n1521) );
  AND2_X2 U1037 ( .A1(WR), .A2(ENABLE), .ZN(n1213) );
  AND2_X2 U1038 ( .A1(RD1), .A2(ENABLE), .ZN(N83) );
  NAND4_X2 U1039 ( .A1(n1592), .A2(n1593), .A3(n1594), .A4(n1595), .ZN(N352)
         );
  NOR4_X2 U1040 ( .A1(n1596), .A2(n1597), .A3(n1598), .A4(n1599), .ZN(n1595)
         );
  OAI221_X2 U1041 ( .B1(n513), .B2(n378), .C1(n481), .C2(n375), .A(n1602), 
        .ZN(n1599) );
  AOI22_X2 U1042 ( .A1(n372), .A2(\registers[19][31] ), .B1(n369), .B2(
        \registers[18][31] ), .ZN(n1602) );
  OAI221_X2 U1043 ( .B1(n641), .B2(n366), .C1(n609), .C2(n363), .A(n1607), 
        .ZN(n1598) );
  AOI22_X2 U1044 ( .A1(n360), .A2(\registers[23][31] ), .B1(n357), .B2(
        \registers[22][31] ), .ZN(n1607) );
  OAI221_X2 U1045 ( .B1(n833), .B2(n354), .C1(n801), .C2(n287), .A(n1612), 
        .ZN(n1597) );
  AOI22_X2 U1046 ( .A1(n284), .A2(\registers[25][31] ), .B1(n281), .B2(
        \registers[24][31] ), .ZN(n1612) );
  OAI221_X2 U1047 ( .B1(n961), .B2(n278), .C1(n929), .C2(n275), .A(n1617), 
        .ZN(n1596) );
  AOI22_X2 U1048 ( .A1(n272), .A2(\registers[29][31] ), .B1(n269), .B2(
        \registers[28][31] ), .ZN(n1617) );
  AOI211_X2 U1049 ( .C1(n266), .C2(\registers[1][31] ), .A(n1621), .B(n1622), 
        .ZN(n1594) );
  OAI22_X2 U1050 ( .A1(n33), .A2(n263), .B1(n65), .B2(n260), .ZN(n1622) );
  OAI221_X2 U1051 ( .B1(n129), .B2(n257), .C1(n97), .C2(n254), .A(n1627), .ZN(
        n1621) );
  AOI22_X2 U1052 ( .A1(n251), .A2(\registers[7][31] ), .B1(n248), .B2(
        \registers[6][31] ), .ZN(n1627) );
  AOI221_X2 U1053 ( .B1(n245), .B2(\registers[13][31] ), .C1(n242), .C2(
        \registers[12][31] ), .A(n1632), .ZN(n1593) );
  OAI22_X2 U1054 ( .A1(n417), .A2(n239), .B1(n449), .B2(n236), .ZN(n1632) );
  AOI221_X2 U1055 ( .B1(n233), .B2(\registers[9][31] ), .C1(n230), .C2(
        \registers[8][31] ), .A(n1637), .ZN(n1592) );
  OAI22_X2 U1056 ( .A1(n289), .A2(n227), .B1(n321), .B2(n224), .ZN(n1637) );
  NAND4_X2 U1057 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .ZN(N351)
         );
  NOR4_X2 U1058 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .ZN(n1643)
         );
  OAI221_X2 U1059 ( .B1(n514), .B2(n378), .C1(n482), .C2(n375), .A(n1648), 
        .ZN(n1647) );
  AOI22_X2 U1060 ( .A1(n372), .A2(\registers[19][30] ), .B1(n369), .B2(
        \registers[18][30] ), .ZN(n1648) );
  OAI221_X2 U1061 ( .B1(n642), .B2(n366), .C1(n610), .C2(n363), .A(n1649), 
        .ZN(n1646) );
  AOI22_X2 U1062 ( .A1(n360), .A2(\registers[23][30] ), .B1(n357), .B2(
        \registers[22][30] ), .ZN(n1649) );
  OAI221_X2 U1063 ( .B1(n834), .B2(n354), .C1(n802), .C2(n287), .A(n1650), 
        .ZN(n1645) );
  AOI22_X2 U1064 ( .A1(n284), .A2(\registers[25][30] ), .B1(n281), .B2(
        \registers[24][30] ), .ZN(n1650) );
  OAI221_X2 U1065 ( .B1(n962), .B2(n278), .C1(n930), .C2(n275), .A(n1651), 
        .ZN(n1644) );
  AOI22_X2 U1066 ( .A1(n272), .A2(\registers[29][30] ), .B1(n269), .B2(
        \registers[28][30] ), .ZN(n1651) );
  AOI211_X2 U1067 ( .C1(n266), .C2(\registers[1][30] ), .A(n1652), .B(n1653), 
        .ZN(n1642) );
  OAI22_X2 U1068 ( .A1(n34), .A2(n263), .B1(n66), .B2(n260), .ZN(n1653) );
  OAI221_X2 U1069 ( .B1(n130), .B2(n257), .C1(n98), .C2(n254), .A(n1654), .ZN(
        n1652) );
  AOI22_X2 U1070 ( .A1(n251), .A2(\registers[7][30] ), .B1(n248), .B2(
        \registers[6][30] ), .ZN(n1654) );
  AOI221_X2 U1071 ( .B1(n245), .B2(\registers[13][30] ), .C1(n242), .C2(
        \registers[12][30] ), .A(n1655), .ZN(n1641) );
  OAI22_X2 U1072 ( .A1(n418), .A2(n239), .B1(n450), .B2(n236), .ZN(n1655) );
  AOI221_X2 U1073 ( .B1(n233), .B2(\registers[9][30] ), .C1(n230), .C2(
        \registers[8][30] ), .A(n1656), .ZN(n1640) );
  OAI22_X2 U1074 ( .A1(n290), .A2(n227), .B1(n322), .B2(n224), .ZN(n1656) );
  NAND4_X2 U1075 ( .A1(n1657), .A2(n1658), .A3(n1659), .A4(n1660), .ZN(N350)
         );
  NOR4_X2 U1076 ( .A1(n1661), .A2(n1662), .A3(n1663), .A4(n1664), .ZN(n1660)
         );
  OAI221_X2 U1077 ( .B1(n515), .B2(n378), .C1(n483), .C2(n375), .A(n1665), 
        .ZN(n1664) );
  AOI22_X2 U1078 ( .A1(n372), .A2(\registers[19][29] ), .B1(n369), .B2(
        \registers[18][29] ), .ZN(n1665) );
  OAI221_X2 U1079 ( .B1(n643), .B2(n366), .C1(n611), .C2(n363), .A(n1666), 
        .ZN(n1663) );
  AOI22_X2 U1080 ( .A1(n360), .A2(\registers[23][29] ), .B1(n357), .B2(
        \registers[22][29] ), .ZN(n1666) );
  OAI221_X2 U1081 ( .B1(n835), .B2(n354), .C1(n803), .C2(n287), .A(n1667), 
        .ZN(n1662) );
  AOI22_X2 U1082 ( .A1(n284), .A2(\registers[25][29] ), .B1(n281), .B2(
        \registers[24][29] ), .ZN(n1667) );
  OAI221_X2 U1083 ( .B1(n963), .B2(n278), .C1(n931), .C2(n275), .A(n1668), 
        .ZN(n1661) );
  AOI22_X2 U1084 ( .A1(n272), .A2(\registers[29][29] ), .B1(n269), .B2(
        \registers[28][29] ), .ZN(n1668) );
  AOI211_X2 U1085 ( .C1(n266), .C2(\registers[1][29] ), .A(n1669), .B(n1670), 
        .ZN(n1659) );
  OAI22_X2 U1086 ( .A1(n35), .A2(n263), .B1(n67), .B2(n260), .ZN(n1670) );
  OAI221_X2 U1087 ( .B1(n131), .B2(n257), .C1(n99), .C2(n254), .A(n1671), .ZN(
        n1669) );
  AOI22_X2 U1088 ( .A1(n251), .A2(\registers[7][29] ), .B1(n248), .B2(
        \registers[6][29] ), .ZN(n1671) );
  AOI221_X2 U1089 ( .B1(n245), .B2(\registers[13][29] ), .C1(n242), .C2(
        \registers[12][29] ), .A(n1672), .ZN(n1658) );
  OAI22_X2 U1090 ( .A1(n419), .A2(n239), .B1(n451), .B2(n236), .ZN(n1672) );
  AOI221_X2 U1091 ( .B1(n233), .B2(\registers[9][29] ), .C1(n230), .C2(
        \registers[8][29] ), .A(n1673), .ZN(n1657) );
  OAI22_X2 U1092 ( .A1(n291), .A2(n227), .B1(n323), .B2(n224), .ZN(n1673) );
  NAND4_X2 U1093 ( .A1(n1674), .A2(n1675), .A3(n1676), .A4(n1677), .ZN(N349)
         );
  NOR4_X2 U1094 ( .A1(n1678), .A2(n1679), .A3(n1680), .A4(n1681), .ZN(n1677)
         );
  OAI221_X2 U1095 ( .B1(n516), .B2(n378), .C1(n484), .C2(n375), .A(n1682), 
        .ZN(n1681) );
  AOI22_X2 U1096 ( .A1(n372), .A2(\registers[19][28] ), .B1(n369), .B2(
        \registers[18][28] ), .ZN(n1682) );
  OAI221_X2 U1097 ( .B1(n644), .B2(n366), .C1(n612), .C2(n363), .A(n1683), 
        .ZN(n1680) );
  AOI22_X2 U1098 ( .A1(n360), .A2(\registers[23][28] ), .B1(n357), .B2(
        \registers[22][28] ), .ZN(n1683) );
  OAI221_X2 U1099 ( .B1(n836), .B2(n354), .C1(n804), .C2(n287), .A(n1684), 
        .ZN(n1679) );
  AOI22_X2 U1100 ( .A1(n284), .A2(\registers[25][28] ), .B1(n281), .B2(
        \registers[24][28] ), .ZN(n1684) );
  OAI221_X2 U1101 ( .B1(n964), .B2(n278), .C1(n932), .C2(n275), .A(n1685), 
        .ZN(n1678) );
  AOI22_X2 U1102 ( .A1(n272), .A2(\registers[29][28] ), .B1(n269), .B2(
        \registers[28][28] ), .ZN(n1685) );
  AOI211_X2 U1103 ( .C1(n266), .C2(\registers[1][28] ), .A(n1686), .B(n1687), 
        .ZN(n1676) );
  OAI22_X2 U1104 ( .A1(n36), .A2(n263), .B1(n68), .B2(n260), .ZN(n1687) );
  OAI221_X2 U1105 ( .B1(n132), .B2(n257), .C1(n100), .C2(n254), .A(n1688), 
        .ZN(n1686) );
  AOI22_X2 U1106 ( .A1(n251), .A2(\registers[7][28] ), .B1(n248), .B2(
        \registers[6][28] ), .ZN(n1688) );
  AOI221_X2 U1107 ( .B1(n245), .B2(\registers[13][28] ), .C1(n242), .C2(
        \registers[12][28] ), .A(n1689), .ZN(n1675) );
  OAI22_X2 U1108 ( .A1(n420), .A2(n239), .B1(n452), .B2(n236), .ZN(n1689) );
  AOI221_X2 U1109 ( .B1(n233), .B2(\registers[9][28] ), .C1(n230), .C2(
        \registers[8][28] ), .A(n1690), .ZN(n1674) );
  OAI22_X2 U1110 ( .A1(n292), .A2(n227), .B1(n324), .B2(n224), .ZN(n1690) );
  NAND4_X2 U1111 ( .A1(n1691), .A2(n1692), .A3(n1693), .A4(n1694), .ZN(N348)
         );
  NOR4_X2 U1112 ( .A1(n1695), .A2(n1696), .A3(n1697), .A4(n1698), .ZN(n1694)
         );
  OAI221_X2 U1113 ( .B1(n517), .B2(n378), .C1(n485), .C2(n375), .A(n1699), 
        .ZN(n1698) );
  AOI22_X2 U1114 ( .A1(n372), .A2(\registers[19][27] ), .B1(n369), .B2(
        \registers[18][27] ), .ZN(n1699) );
  OAI221_X2 U1115 ( .B1(n645), .B2(n366), .C1(n613), .C2(n363), .A(n1700), 
        .ZN(n1697) );
  AOI22_X2 U1116 ( .A1(n360), .A2(\registers[23][27] ), .B1(n357), .B2(
        \registers[22][27] ), .ZN(n1700) );
  OAI221_X2 U1117 ( .B1(n837), .B2(n354), .C1(n805), .C2(n287), .A(n1701), 
        .ZN(n1696) );
  AOI22_X2 U1118 ( .A1(n284), .A2(\registers[25][27] ), .B1(n281), .B2(
        \registers[24][27] ), .ZN(n1701) );
  OAI221_X2 U1119 ( .B1(n965), .B2(n278), .C1(n933), .C2(n275), .A(n1702), 
        .ZN(n1695) );
  AOI22_X2 U1120 ( .A1(n272), .A2(\registers[29][27] ), .B1(n269), .B2(
        \registers[28][27] ), .ZN(n1702) );
  AOI211_X2 U1121 ( .C1(n266), .C2(\registers[1][27] ), .A(n1703), .B(n1704), 
        .ZN(n1693) );
  OAI22_X2 U1122 ( .A1(n37), .A2(n263), .B1(n69), .B2(n260), .ZN(n1704) );
  OAI221_X2 U1123 ( .B1(n133), .B2(n257), .C1(n101), .C2(n254), .A(n1705), 
        .ZN(n1703) );
  AOI22_X2 U1124 ( .A1(n251), .A2(\registers[7][27] ), .B1(n248), .B2(
        \registers[6][27] ), .ZN(n1705) );
  AOI221_X2 U1125 ( .B1(n245), .B2(\registers[13][27] ), .C1(n242), .C2(
        \registers[12][27] ), .A(n1706), .ZN(n1692) );
  OAI22_X2 U1126 ( .A1(n421), .A2(n239), .B1(n453), .B2(n236), .ZN(n1706) );
  AOI221_X2 U1127 ( .B1(n233), .B2(\registers[9][27] ), .C1(n230), .C2(
        \registers[8][27] ), .A(n1707), .ZN(n1691) );
  OAI22_X2 U1128 ( .A1(n293), .A2(n227), .B1(n325), .B2(n224), .ZN(n1707) );
  NAND4_X2 U1129 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(N347)
         );
  NOR4_X2 U1130 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711)
         );
  OAI221_X2 U1131 ( .B1(n518), .B2(n378), .C1(n486), .C2(n375), .A(n1716), 
        .ZN(n1715) );
  AOI22_X2 U1132 ( .A1(n372), .A2(\registers[19][26] ), .B1(n369), .B2(
        \registers[18][26] ), .ZN(n1716) );
  OAI221_X2 U1133 ( .B1(n646), .B2(n366), .C1(n614), .C2(n363), .A(n1717), 
        .ZN(n1714) );
  AOI22_X2 U1134 ( .A1(n360), .A2(\registers[23][26] ), .B1(n357), .B2(
        \registers[22][26] ), .ZN(n1717) );
  OAI221_X2 U1135 ( .B1(n838), .B2(n354), .C1(n806), .C2(n287), .A(n1718), 
        .ZN(n1713) );
  AOI22_X2 U1136 ( .A1(n284), .A2(\registers[25][26] ), .B1(n281), .B2(
        \registers[24][26] ), .ZN(n1718) );
  OAI221_X2 U1137 ( .B1(n966), .B2(n278), .C1(n934), .C2(n275), .A(n1719), 
        .ZN(n1712) );
  AOI22_X2 U1138 ( .A1(n272), .A2(\registers[29][26] ), .B1(n269), .B2(
        \registers[28][26] ), .ZN(n1719) );
  AOI211_X2 U1139 ( .C1(n266), .C2(\registers[1][26] ), .A(n1720), .B(n1721), 
        .ZN(n1710) );
  OAI22_X2 U1140 ( .A1(n38), .A2(n263), .B1(n70), .B2(n260), .ZN(n1721) );
  OAI221_X2 U1141 ( .B1(n134), .B2(n257), .C1(n102), .C2(n254), .A(n1722), 
        .ZN(n1720) );
  AOI22_X2 U1142 ( .A1(n251), .A2(\registers[7][26] ), .B1(n248), .B2(
        \registers[6][26] ), .ZN(n1722) );
  AOI221_X2 U1143 ( .B1(n245), .B2(\registers[13][26] ), .C1(n242), .C2(
        \registers[12][26] ), .A(n1723), .ZN(n1709) );
  OAI22_X2 U1144 ( .A1(n422), .A2(n239), .B1(n454), .B2(n236), .ZN(n1723) );
  AOI221_X2 U1145 ( .B1(n233), .B2(\registers[9][26] ), .C1(n230), .C2(
        \registers[8][26] ), .A(n1724), .ZN(n1708) );
  OAI22_X2 U1146 ( .A1(n294), .A2(n227), .B1(n326), .B2(n224), .ZN(n1724) );
  NAND4_X2 U1147 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(N346)
         );
  NOR4_X2 U1148 ( .A1(n1729), .A2(n1730), .A3(n1731), .A4(n1732), .ZN(n1728)
         );
  OAI221_X2 U1149 ( .B1(n519), .B2(n378), .C1(n487), .C2(n375), .A(n1733), 
        .ZN(n1732) );
  AOI22_X2 U1150 ( .A1(n372), .A2(\registers[19][25] ), .B1(n369), .B2(
        \registers[18][25] ), .ZN(n1733) );
  OAI221_X2 U1151 ( .B1(n647), .B2(n366), .C1(n615), .C2(n363), .A(n1734), 
        .ZN(n1731) );
  AOI22_X2 U1152 ( .A1(n360), .A2(\registers[23][25] ), .B1(n357), .B2(
        \registers[22][25] ), .ZN(n1734) );
  OAI221_X2 U1153 ( .B1(n839), .B2(n354), .C1(n807), .C2(n287), .A(n1735), 
        .ZN(n1730) );
  AOI22_X2 U1154 ( .A1(n284), .A2(\registers[25][25] ), .B1(n281), .B2(
        \registers[24][25] ), .ZN(n1735) );
  OAI221_X2 U1155 ( .B1(n967), .B2(n278), .C1(n935), .C2(n275), .A(n1736), 
        .ZN(n1729) );
  AOI22_X2 U1156 ( .A1(n272), .A2(\registers[29][25] ), .B1(n269), .B2(
        \registers[28][25] ), .ZN(n1736) );
  AOI211_X2 U1157 ( .C1(n266), .C2(\registers[1][25] ), .A(n1737), .B(n1738), 
        .ZN(n1727) );
  OAI22_X2 U1158 ( .A1(n39), .A2(n263), .B1(n71), .B2(n260), .ZN(n1738) );
  OAI221_X2 U1159 ( .B1(n135), .B2(n257), .C1(n103), .C2(n254), .A(n1739), 
        .ZN(n1737) );
  AOI22_X2 U1160 ( .A1(n251), .A2(\registers[7][25] ), .B1(n248), .B2(
        \registers[6][25] ), .ZN(n1739) );
  AOI221_X2 U1161 ( .B1(n245), .B2(\registers[13][25] ), .C1(n242), .C2(
        \registers[12][25] ), .A(n1740), .ZN(n1726) );
  OAI22_X2 U1162 ( .A1(n423), .A2(n239), .B1(n455), .B2(n236), .ZN(n1740) );
  AOI221_X2 U1163 ( .B1(n233), .B2(\registers[9][25] ), .C1(n230), .C2(
        \registers[8][25] ), .A(n1741), .ZN(n1725) );
  OAI22_X2 U1164 ( .A1(n295), .A2(n227), .B1(n327), .B2(n224), .ZN(n1741) );
  NAND4_X2 U1165 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(N345)
         );
  NOR4_X2 U1166 ( .A1(n1746), .A2(n1747), .A3(n1748), .A4(n1749), .ZN(n1745)
         );
  OAI221_X2 U1167 ( .B1(n520), .B2(n378), .C1(n488), .C2(n375), .A(n1750), 
        .ZN(n1749) );
  AOI22_X2 U1168 ( .A1(n372), .A2(\registers[19][24] ), .B1(n369), .B2(
        \registers[18][24] ), .ZN(n1750) );
  OAI221_X2 U1169 ( .B1(n648), .B2(n366), .C1(n616), .C2(n363), .A(n1751), 
        .ZN(n1748) );
  AOI22_X2 U1170 ( .A1(n360), .A2(\registers[23][24] ), .B1(n357), .B2(
        \registers[22][24] ), .ZN(n1751) );
  OAI221_X2 U1171 ( .B1(n840), .B2(n354), .C1(n808), .C2(n287), .A(n1752), 
        .ZN(n1747) );
  AOI22_X2 U1172 ( .A1(n284), .A2(\registers[25][24] ), .B1(n281), .B2(
        \registers[24][24] ), .ZN(n1752) );
  OAI221_X2 U1173 ( .B1(n968), .B2(n278), .C1(n936), .C2(n275), .A(n1753), 
        .ZN(n1746) );
  AOI22_X2 U1174 ( .A1(n272), .A2(\registers[29][24] ), .B1(n269), .B2(
        \registers[28][24] ), .ZN(n1753) );
  AOI211_X2 U1175 ( .C1(n266), .C2(\registers[1][24] ), .A(n1754), .B(n1755), 
        .ZN(n1744) );
  OAI22_X2 U1176 ( .A1(n40), .A2(n263), .B1(n72), .B2(n260), .ZN(n1755) );
  OAI221_X2 U1177 ( .B1(n136), .B2(n257), .C1(n104), .C2(n254), .A(n1756), 
        .ZN(n1754) );
  AOI22_X2 U1178 ( .A1(n251), .A2(\registers[7][24] ), .B1(n248), .B2(
        \registers[6][24] ), .ZN(n1756) );
  AOI221_X2 U1179 ( .B1(n245), .B2(\registers[13][24] ), .C1(n242), .C2(
        \registers[12][24] ), .A(n1757), .ZN(n1743) );
  OAI22_X2 U1180 ( .A1(n424), .A2(n239), .B1(n456), .B2(n236), .ZN(n1757) );
  AOI221_X2 U1181 ( .B1(n233), .B2(\registers[9][24] ), .C1(n230), .C2(
        \registers[8][24] ), .A(n1758), .ZN(n1742) );
  OAI22_X2 U1182 ( .A1(n296), .A2(n227), .B1(n328), .B2(n224), .ZN(n1758) );
  NAND4_X2 U1183 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(N344)
         );
  NOR4_X2 U1184 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .ZN(n1762)
         );
  OAI221_X2 U1185 ( .B1(n521), .B2(n378), .C1(n489), .C2(n375), .A(n1767), 
        .ZN(n1766) );
  AOI22_X2 U1186 ( .A1(n372), .A2(\registers[19][23] ), .B1(n369), .B2(
        \registers[18][23] ), .ZN(n1767) );
  OAI221_X2 U1187 ( .B1(n649), .B2(n366), .C1(n617), .C2(n363), .A(n1768), 
        .ZN(n1765) );
  AOI22_X2 U1188 ( .A1(n360), .A2(\registers[23][23] ), .B1(n357), .B2(
        \registers[22][23] ), .ZN(n1768) );
  OAI221_X2 U1189 ( .B1(n841), .B2(n354), .C1(n809), .C2(n287), .A(n1769), 
        .ZN(n1764) );
  AOI22_X2 U1190 ( .A1(n284), .A2(\registers[25][23] ), .B1(n281), .B2(
        \registers[24][23] ), .ZN(n1769) );
  OAI221_X2 U1191 ( .B1(n969), .B2(n278), .C1(n937), .C2(n275), .A(n1770), 
        .ZN(n1763) );
  AOI22_X2 U1192 ( .A1(n272), .A2(\registers[29][23] ), .B1(n269), .B2(
        \registers[28][23] ), .ZN(n1770) );
  AOI211_X2 U1193 ( .C1(n266), .C2(\registers[1][23] ), .A(n1771), .B(n1772), 
        .ZN(n1761) );
  OAI22_X2 U1194 ( .A1(n41), .A2(n262), .B1(n73), .B2(n259), .ZN(n1772) );
  OAI221_X2 U1195 ( .B1(n137), .B2(n257), .C1(n105), .C2(n254), .A(n1773), 
        .ZN(n1771) );
  AOI22_X2 U1196 ( .A1(n251), .A2(\registers[7][23] ), .B1(n248), .B2(
        \registers[6][23] ), .ZN(n1773) );
  AOI221_X2 U1197 ( .B1(n245), .B2(\registers[13][23] ), .C1(n242), .C2(
        \registers[12][23] ), .A(n1774), .ZN(n1760) );
  OAI22_X2 U1198 ( .A1(n425), .A2(n238), .B1(n457), .B2(n235), .ZN(n1774) );
  AOI221_X2 U1199 ( .B1(n233), .B2(\registers[9][23] ), .C1(n230), .C2(
        \registers[8][23] ), .A(n1775), .ZN(n1759) );
  OAI22_X2 U1200 ( .A1(n297), .A2(n226), .B1(n329), .B2(n223), .ZN(n1775) );
  NAND4_X2 U1201 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(N343)
         );
  NOR4_X2 U1202 ( .A1(n1780), .A2(n1781), .A3(n1782), .A4(n1783), .ZN(n1779)
         );
  OAI221_X2 U1203 ( .B1(n522), .B2(n378), .C1(n490), .C2(n375), .A(n1784), 
        .ZN(n1783) );
  AOI22_X2 U1204 ( .A1(n372), .A2(\registers[19][22] ), .B1(n369), .B2(
        \registers[18][22] ), .ZN(n1784) );
  OAI221_X2 U1205 ( .B1(n650), .B2(n366), .C1(n618), .C2(n363), .A(n1785), 
        .ZN(n1782) );
  AOI22_X2 U1206 ( .A1(n360), .A2(\registers[23][22] ), .B1(n357), .B2(
        \registers[22][22] ), .ZN(n1785) );
  OAI221_X2 U1207 ( .B1(n842), .B2(n354), .C1(n810), .C2(n287), .A(n1786), 
        .ZN(n1781) );
  AOI22_X2 U1208 ( .A1(n284), .A2(\registers[25][22] ), .B1(n281), .B2(
        \registers[24][22] ), .ZN(n1786) );
  OAI221_X2 U1209 ( .B1(n970), .B2(n278), .C1(n938), .C2(n275), .A(n1787), 
        .ZN(n1780) );
  AOI22_X2 U1210 ( .A1(n272), .A2(\registers[29][22] ), .B1(n269), .B2(
        \registers[28][22] ), .ZN(n1787) );
  AOI211_X2 U1211 ( .C1(n266), .C2(\registers[1][22] ), .A(n1788), .B(n1789), 
        .ZN(n1778) );
  OAI22_X2 U1212 ( .A1(n42), .A2(n262), .B1(n74), .B2(n259), .ZN(n1789) );
  OAI221_X2 U1213 ( .B1(n138), .B2(n257), .C1(n106), .C2(n254), .A(n1790), 
        .ZN(n1788) );
  AOI22_X2 U1214 ( .A1(n251), .A2(\registers[7][22] ), .B1(n248), .B2(
        \registers[6][22] ), .ZN(n1790) );
  AOI221_X2 U1215 ( .B1(n245), .B2(\registers[13][22] ), .C1(n242), .C2(
        \registers[12][22] ), .A(n1791), .ZN(n1777) );
  OAI22_X2 U1216 ( .A1(n426), .A2(n238), .B1(n458), .B2(n235), .ZN(n1791) );
  AOI221_X2 U1217 ( .B1(n233), .B2(\registers[9][22] ), .C1(n230), .C2(
        \registers[8][22] ), .A(n1792), .ZN(n1776) );
  OAI22_X2 U1218 ( .A1(n298), .A2(n226), .B1(n330), .B2(n223), .ZN(n1792) );
  NAND4_X2 U1219 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .ZN(N342)
         );
  NOR4_X2 U1220 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1796)
         );
  OAI221_X2 U1221 ( .B1(n523), .B2(n377), .C1(n491), .C2(n374), .A(n1801), 
        .ZN(n1800) );
  AOI22_X2 U1222 ( .A1(n371), .A2(\registers[19][21] ), .B1(n368), .B2(
        \registers[18][21] ), .ZN(n1801) );
  OAI221_X2 U1223 ( .B1(n651), .B2(n365), .C1(n619), .C2(n362), .A(n1802), 
        .ZN(n1799) );
  AOI22_X2 U1224 ( .A1(n359), .A2(\registers[23][21] ), .B1(n356), .B2(
        \registers[22][21] ), .ZN(n1802) );
  OAI221_X2 U1225 ( .B1(n843), .B2(n353), .C1(n811), .C2(n286), .A(n1803), 
        .ZN(n1798) );
  AOI22_X2 U1226 ( .A1(n283), .A2(\registers[25][21] ), .B1(n280), .B2(
        \registers[24][21] ), .ZN(n1803) );
  OAI221_X2 U1227 ( .B1(n971), .B2(n277), .C1(n939), .C2(n274), .A(n1804), 
        .ZN(n1797) );
  AOI22_X2 U1228 ( .A1(n271), .A2(\registers[29][21] ), .B1(n268), .B2(
        \registers[28][21] ), .ZN(n1804) );
  AOI211_X2 U1229 ( .C1(n265), .C2(\registers[1][21] ), .A(n1805), .B(n1806), 
        .ZN(n1795) );
  OAI22_X2 U1230 ( .A1(n43), .A2(n262), .B1(n75), .B2(n259), .ZN(n1806) );
  OAI221_X2 U1231 ( .B1(n139), .B2(n256), .C1(n107), .C2(n253), .A(n1807), 
        .ZN(n1805) );
  AOI22_X2 U1232 ( .A1(n250), .A2(\registers[7][21] ), .B1(n247), .B2(
        \registers[6][21] ), .ZN(n1807) );
  AOI221_X2 U1233 ( .B1(n244), .B2(\registers[13][21] ), .C1(n241), .C2(
        \registers[12][21] ), .A(n1808), .ZN(n1794) );
  OAI22_X2 U1234 ( .A1(n427), .A2(n238), .B1(n459), .B2(n235), .ZN(n1808) );
  AOI221_X2 U1235 ( .B1(n232), .B2(\registers[9][21] ), .C1(n229), .C2(
        \registers[8][21] ), .A(n1809), .ZN(n1793) );
  OAI22_X2 U1236 ( .A1(n299), .A2(n226), .B1(n331), .B2(n223), .ZN(n1809) );
  NAND4_X2 U1237 ( .A1(n1810), .A2(n1811), .A3(n1812), .A4(n1813), .ZN(N341)
         );
  NOR4_X2 U1238 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .ZN(n1813)
         );
  OAI221_X2 U1239 ( .B1(n524), .B2(n377), .C1(n492), .C2(n374), .A(n1818), 
        .ZN(n1817) );
  AOI22_X2 U1240 ( .A1(n371), .A2(\registers[19][20] ), .B1(n368), .B2(
        \registers[18][20] ), .ZN(n1818) );
  OAI221_X2 U1241 ( .B1(n652), .B2(n365), .C1(n620), .C2(n362), .A(n1819), 
        .ZN(n1816) );
  AOI22_X2 U1242 ( .A1(n359), .A2(\registers[23][20] ), .B1(n356), .B2(
        \registers[22][20] ), .ZN(n1819) );
  OAI221_X2 U1243 ( .B1(n844), .B2(n353), .C1(n812), .C2(n286), .A(n1820), 
        .ZN(n1815) );
  AOI22_X2 U1244 ( .A1(n283), .A2(\registers[25][20] ), .B1(n280), .B2(
        \registers[24][20] ), .ZN(n1820) );
  OAI221_X2 U1245 ( .B1(n972), .B2(n277), .C1(n940), .C2(n274), .A(n1821), 
        .ZN(n1814) );
  AOI22_X2 U1246 ( .A1(n271), .A2(\registers[29][20] ), .B1(n268), .B2(
        \registers[28][20] ), .ZN(n1821) );
  AOI211_X2 U1247 ( .C1(n265), .C2(\registers[1][20] ), .A(n1822), .B(n1823), 
        .ZN(n1812) );
  OAI22_X2 U1248 ( .A1(n44), .A2(n262), .B1(n76), .B2(n259), .ZN(n1823) );
  OAI221_X2 U1249 ( .B1(n140), .B2(n256), .C1(n108), .C2(n253), .A(n1824), 
        .ZN(n1822) );
  AOI22_X2 U1250 ( .A1(n250), .A2(\registers[7][20] ), .B1(n247), .B2(
        \registers[6][20] ), .ZN(n1824) );
  AOI221_X2 U1251 ( .B1(n244), .B2(\registers[13][20] ), .C1(n241), .C2(
        \registers[12][20] ), .A(n1825), .ZN(n1811) );
  OAI22_X2 U1252 ( .A1(n428), .A2(n238), .B1(n460), .B2(n235), .ZN(n1825) );
  AOI221_X2 U1253 ( .B1(n232), .B2(\registers[9][20] ), .C1(n229), .C2(
        \registers[8][20] ), .A(n1826), .ZN(n1810) );
  OAI22_X2 U1254 ( .A1(n300), .A2(n226), .B1(n332), .B2(n223), .ZN(n1826) );
  NAND4_X2 U1255 ( .A1(n1827), .A2(n1828), .A3(n1829), .A4(n1830), .ZN(N340)
         );
  NOR4_X2 U1256 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(n1830)
         );
  OAI221_X2 U1257 ( .B1(n525), .B2(n377), .C1(n493), .C2(n374), .A(n1835), 
        .ZN(n1834) );
  AOI22_X2 U1258 ( .A1(n371), .A2(\registers[19][19] ), .B1(n368), .B2(
        \registers[18][19] ), .ZN(n1835) );
  OAI221_X2 U1259 ( .B1(n653), .B2(n365), .C1(n621), .C2(n362), .A(n1836), 
        .ZN(n1833) );
  AOI22_X2 U1260 ( .A1(n359), .A2(\registers[23][19] ), .B1(n356), .B2(
        \registers[22][19] ), .ZN(n1836) );
  OAI221_X2 U1261 ( .B1(n845), .B2(n353), .C1(n813), .C2(n286), .A(n1837), 
        .ZN(n1832) );
  AOI22_X2 U1262 ( .A1(n283), .A2(\registers[25][19] ), .B1(n280), .B2(
        \registers[24][19] ), .ZN(n1837) );
  OAI221_X2 U1263 ( .B1(n973), .B2(n277), .C1(n941), .C2(n274), .A(n1838), 
        .ZN(n1831) );
  AOI22_X2 U1264 ( .A1(n271), .A2(\registers[29][19] ), .B1(n268), .B2(
        \registers[28][19] ), .ZN(n1838) );
  AOI211_X2 U1265 ( .C1(n265), .C2(\registers[1][19] ), .A(n1839), .B(n1840), 
        .ZN(n1829) );
  OAI22_X2 U1266 ( .A1(n45), .A2(n262), .B1(n77), .B2(n259), .ZN(n1840) );
  OAI221_X2 U1267 ( .B1(n141), .B2(n256), .C1(n109), .C2(n253), .A(n1841), 
        .ZN(n1839) );
  AOI22_X2 U1268 ( .A1(n250), .A2(\registers[7][19] ), .B1(n247), .B2(
        \registers[6][19] ), .ZN(n1841) );
  AOI221_X2 U1269 ( .B1(n244), .B2(\registers[13][19] ), .C1(n241), .C2(
        \registers[12][19] ), .A(n1842), .ZN(n1828) );
  OAI22_X2 U1270 ( .A1(n429), .A2(n238), .B1(n461), .B2(n235), .ZN(n1842) );
  AOI221_X2 U1271 ( .B1(n232), .B2(\registers[9][19] ), .C1(n229), .C2(
        \registers[8][19] ), .A(n1843), .ZN(n1827) );
  OAI22_X2 U1272 ( .A1(n301), .A2(n226), .B1(n333), .B2(n223), .ZN(n1843) );
  NAND4_X2 U1273 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .ZN(N339)
         );
  NOR4_X2 U1274 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1847)
         );
  OAI221_X2 U1275 ( .B1(n526), .B2(n377), .C1(n494), .C2(n374), .A(n1852), 
        .ZN(n1851) );
  AOI22_X2 U1276 ( .A1(n371), .A2(\registers[19][18] ), .B1(n368), .B2(
        \registers[18][18] ), .ZN(n1852) );
  OAI221_X2 U1277 ( .B1(n654), .B2(n365), .C1(n622), .C2(n362), .A(n1853), 
        .ZN(n1850) );
  AOI22_X2 U1278 ( .A1(n359), .A2(\registers[23][18] ), .B1(n356), .B2(
        \registers[22][18] ), .ZN(n1853) );
  OAI221_X2 U1279 ( .B1(n846), .B2(n353), .C1(n814), .C2(n286), .A(n1854), 
        .ZN(n1849) );
  AOI22_X2 U1280 ( .A1(n283), .A2(\registers[25][18] ), .B1(n280), .B2(
        \registers[24][18] ), .ZN(n1854) );
  OAI221_X2 U1281 ( .B1(n974), .B2(n277), .C1(n942), .C2(n274), .A(n1855), 
        .ZN(n1848) );
  AOI22_X2 U1282 ( .A1(n271), .A2(\registers[29][18] ), .B1(n268), .B2(
        \registers[28][18] ), .ZN(n1855) );
  AOI211_X2 U1283 ( .C1(n265), .C2(\registers[1][18] ), .A(n1856), .B(n1857), 
        .ZN(n1846) );
  OAI22_X2 U1284 ( .A1(n46), .A2(n262), .B1(n78), .B2(n259), .ZN(n1857) );
  OAI221_X2 U1285 ( .B1(n142), .B2(n256), .C1(n110), .C2(n253), .A(n1858), 
        .ZN(n1856) );
  AOI22_X2 U1286 ( .A1(n250), .A2(\registers[7][18] ), .B1(n247), .B2(
        \registers[6][18] ), .ZN(n1858) );
  AOI221_X2 U1287 ( .B1(n244), .B2(\registers[13][18] ), .C1(n241), .C2(
        \registers[12][18] ), .A(n1859), .ZN(n1845) );
  OAI22_X2 U1288 ( .A1(n430), .A2(n238), .B1(n462), .B2(n235), .ZN(n1859) );
  AOI221_X2 U1289 ( .B1(n232), .B2(\registers[9][18] ), .C1(n229), .C2(
        \registers[8][18] ), .A(n1860), .ZN(n1844) );
  OAI22_X2 U1290 ( .A1(n302), .A2(n226), .B1(n334), .B2(n223), .ZN(n1860) );
  NAND4_X2 U1291 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .ZN(N338)
         );
  NOR4_X2 U1292 ( .A1(n1865), .A2(n1866), .A3(n1867), .A4(n1868), .ZN(n1864)
         );
  OAI221_X2 U1293 ( .B1(n527), .B2(n377), .C1(n495), .C2(n374), .A(n1869), 
        .ZN(n1868) );
  AOI22_X2 U1294 ( .A1(n371), .A2(\registers[19][17] ), .B1(n368), .B2(
        \registers[18][17] ), .ZN(n1869) );
  OAI221_X2 U1295 ( .B1(n655), .B2(n365), .C1(n623), .C2(n362), .A(n1870), 
        .ZN(n1867) );
  AOI22_X2 U1296 ( .A1(n359), .A2(\registers[23][17] ), .B1(n356), .B2(
        \registers[22][17] ), .ZN(n1870) );
  OAI221_X2 U1297 ( .B1(n847), .B2(n353), .C1(n815), .C2(n286), .A(n1871), 
        .ZN(n1866) );
  AOI22_X2 U1298 ( .A1(n283), .A2(\registers[25][17] ), .B1(n280), .B2(
        \registers[24][17] ), .ZN(n1871) );
  OAI221_X2 U1299 ( .B1(n975), .B2(n277), .C1(n943), .C2(n274), .A(n1872), 
        .ZN(n1865) );
  AOI22_X2 U1300 ( .A1(n271), .A2(\registers[29][17] ), .B1(n268), .B2(
        \registers[28][17] ), .ZN(n1872) );
  AOI211_X2 U1301 ( .C1(n265), .C2(\registers[1][17] ), .A(n1873), .B(n1874), 
        .ZN(n1863) );
  OAI22_X2 U1302 ( .A1(n47), .A2(n262), .B1(n79), .B2(n259), .ZN(n1874) );
  OAI221_X2 U1303 ( .B1(n143), .B2(n256), .C1(n111), .C2(n253), .A(n1875), 
        .ZN(n1873) );
  AOI22_X2 U1304 ( .A1(n250), .A2(\registers[7][17] ), .B1(n247), .B2(
        \registers[6][17] ), .ZN(n1875) );
  AOI221_X2 U1305 ( .B1(n244), .B2(\registers[13][17] ), .C1(n241), .C2(
        \registers[12][17] ), .A(n1876), .ZN(n1862) );
  OAI22_X2 U1306 ( .A1(n431), .A2(n238), .B1(n463), .B2(n235), .ZN(n1876) );
  AOI221_X2 U1307 ( .B1(n232), .B2(\registers[9][17] ), .C1(n229), .C2(
        \registers[8][17] ), .A(n1877), .ZN(n1861) );
  OAI22_X2 U1308 ( .A1(n303), .A2(n226), .B1(n335), .B2(n223), .ZN(n1877) );
  NAND4_X2 U1309 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .ZN(N337)
         );
  NOR4_X2 U1310 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .ZN(n1881)
         );
  OAI221_X2 U1311 ( .B1(n528), .B2(n377), .C1(n496), .C2(n374), .A(n1886), 
        .ZN(n1885) );
  AOI22_X2 U1312 ( .A1(n371), .A2(\registers[19][16] ), .B1(n368), .B2(
        \registers[18][16] ), .ZN(n1886) );
  OAI221_X2 U1313 ( .B1(n656), .B2(n365), .C1(n624), .C2(n362), .A(n1887), 
        .ZN(n1884) );
  AOI22_X2 U1314 ( .A1(n359), .A2(\registers[23][16] ), .B1(n356), .B2(
        \registers[22][16] ), .ZN(n1887) );
  OAI221_X2 U1315 ( .B1(n848), .B2(n353), .C1(n816), .C2(n286), .A(n1888), 
        .ZN(n1883) );
  AOI22_X2 U1316 ( .A1(n283), .A2(\registers[25][16] ), .B1(n280), .B2(
        \registers[24][16] ), .ZN(n1888) );
  OAI221_X2 U1317 ( .B1(n976), .B2(n277), .C1(n944), .C2(n274), .A(n1889), 
        .ZN(n1882) );
  AOI22_X2 U1318 ( .A1(n271), .A2(\registers[29][16] ), .B1(n268), .B2(
        \registers[28][16] ), .ZN(n1889) );
  AOI211_X2 U1319 ( .C1(n265), .C2(\registers[1][16] ), .A(n1890), .B(n1891), 
        .ZN(n1880) );
  OAI22_X2 U1320 ( .A1(n48), .A2(n262), .B1(n80), .B2(n259), .ZN(n1891) );
  OAI221_X2 U1321 ( .B1(n144), .B2(n256), .C1(n112), .C2(n253), .A(n1892), 
        .ZN(n1890) );
  AOI22_X2 U1322 ( .A1(n250), .A2(\registers[7][16] ), .B1(n247), .B2(
        \registers[6][16] ), .ZN(n1892) );
  AOI221_X2 U1323 ( .B1(n244), .B2(\registers[13][16] ), .C1(n241), .C2(
        \registers[12][16] ), .A(n1893), .ZN(n1879) );
  OAI22_X2 U1324 ( .A1(n432), .A2(n238), .B1(n464), .B2(n235), .ZN(n1893) );
  AOI221_X2 U1325 ( .B1(n232), .B2(\registers[9][16] ), .C1(n229), .C2(
        \registers[8][16] ), .A(n1894), .ZN(n1878) );
  OAI22_X2 U1326 ( .A1(n304), .A2(n226), .B1(n336), .B2(n223), .ZN(n1894) );
  NAND4_X2 U1327 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(N336)
         );
  NOR4_X2 U1328 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898)
         );
  OAI221_X2 U1329 ( .B1(n529), .B2(n377), .C1(n497), .C2(n374), .A(n1903), 
        .ZN(n1902) );
  AOI22_X2 U1330 ( .A1(n371), .A2(\registers[19][15] ), .B1(n368), .B2(
        \registers[18][15] ), .ZN(n1903) );
  OAI221_X2 U1331 ( .B1(n657), .B2(n365), .C1(n625), .C2(n362), .A(n1904), 
        .ZN(n1901) );
  AOI22_X2 U1332 ( .A1(n359), .A2(\registers[23][15] ), .B1(n356), .B2(
        \registers[22][15] ), .ZN(n1904) );
  OAI221_X2 U1333 ( .B1(n849), .B2(n353), .C1(n817), .C2(n286), .A(n1905), 
        .ZN(n1900) );
  AOI22_X2 U1334 ( .A1(n283), .A2(\registers[25][15] ), .B1(n280), .B2(
        \registers[24][15] ), .ZN(n1905) );
  OAI221_X2 U1335 ( .B1(n977), .B2(n277), .C1(n945), .C2(n274), .A(n1906), 
        .ZN(n1899) );
  AOI22_X2 U1336 ( .A1(n271), .A2(\registers[29][15] ), .B1(n268), .B2(
        \registers[28][15] ), .ZN(n1906) );
  AOI211_X2 U1337 ( .C1(n265), .C2(\registers[1][15] ), .A(n1907), .B(n1908), 
        .ZN(n1897) );
  OAI22_X2 U1338 ( .A1(n49), .A2(n262), .B1(n81), .B2(n259), .ZN(n1908) );
  OAI221_X2 U1339 ( .B1(n145), .B2(n256), .C1(n113), .C2(n253), .A(n1909), 
        .ZN(n1907) );
  AOI22_X2 U1340 ( .A1(n250), .A2(\registers[7][15] ), .B1(n247), .B2(
        \registers[6][15] ), .ZN(n1909) );
  AOI221_X2 U1341 ( .B1(n244), .B2(\registers[13][15] ), .C1(n241), .C2(
        \registers[12][15] ), .A(n1910), .ZN(n1896) );
  OAI22_X2 U1342 ( .A1(n433), .A2(n238), .B1(n465), .B2(n235), .ZN(n1910) );
  AOI221_X2 U1343 ( .B1(n232), .B2(\registers[9][15] ), .C1(n229), .C2(
        \registers[8][15] ), .A(n1911), .ZN(n1895) );
  OAI22_X2 U1344 ( .A1(n305), .A2(n226), .B1(n337), .B2(n223), .ZN(n1911) );
  NAND4_X2 U1345 ( .A1(n1912), .A2(n1913), .A3(n1914), .A4(n1915), .ZN(N335)
         );
  NOR4_X2 U1346 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(n1915)
         );
  OAI221_X2 U1347 ( .B1(n530), .B2(n377), .C1(n498), .C2(n374), .A(n1920), 
        .ZN(n1919) );
  AOI22_X2 U1348 ( .A1(n371), .A2(\registers[19][14] ), .B1(n368), .B2(
        \registers[18][14] ), .ZN(n1920) );
  OAI221_X2 U1349 ( .B1(n658), .B2(n365), .C1(n626), .C2(n362), .A(n1921), 
        .ZN(n1918) );
  AOI22_X2 U1350 ( .A1(n359), .A2(\registers[23][14] ), .B1(n356), .B2(
        \registers[22][14] ), .ZN(n1921) );
  OAI221_X2 U1351 ( .B1(n850), .B2(n353), .C1(n818), .C2(n286), .A(n1922), 
        .ZN(n1917) );
  AOI22_X2 U1352 ( .A1(n283), .A2(\registers[25][14] ), .B1(n280), .B2(
        \registers[24][14] ), .ZN(n1922) );
  OAI221_X2 U1353 ( .B1(n978), .B2(n277), .C1(n946), .C2(n274), .A(n1923), 
        .ZN(n1916) );
  AOI22_X2 U1354 ( .A1(n271), .A2(\registers[29][14] ), .B1(n268), .B2(
        \registers[28][14] ), .ZN(n1923) );
  AOI211_X2 U1355 ( .C1(n265), .C2(\registers[1][14] ), .A(n1924), .B(n1925), 
        .ZN(n1914) );
  OAI22_X2 U1356 ( .A1(n50), .A2(n262), .B1(n82), .B2(n259), .ZN(n1925) );
  OAI221_X2 U1357 ( .B1(n146), .B2(n256), .C1(n114), .C2(n253), .A(n1926), 
        .ZN(n1924) );
  AOI22_X2 U1358 ( .A1(n250), .A2(\registers[7][14] ), .B1(n247), .B2(
        \registers[6][14] ), .ZN(n1926) );
  AOI221_X2 U1359 ( .B1(n244), .B2(\registers[13][14] ), .C1(n241), .C2(
        \registers[12][14] ), .A(n1927), .ZN(n1913) );
  OAI22_X2 U1360 ( .A1(n434), .A2(n238), .B1(n466), .B2(n235), .ZN(n1927) );
  AOI221_X2 U1361 ( .B1(n232), .B2(\registers[9][14] ), .C1(n229), .C2(
        \registers[8][14] ), .A(n1928), .ZN(n1912) );
  OAI22_X2 U1362 ( .A1(n306), .A2(n226), .B1(n338), .B2(n223), .ZN(n1928) );
  NAND4_X2 U1363 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(N334)
         );
  NOR4_X2 U1364 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(n1932)
         );
  OAI221_X2 U1365 ( .B1(n531), .B2(n377), .C1(n499), .C2(n374), .A(n1937), 
        .ZN(n1936) );
  AOI22_X2 U1366 ( .A1(n371), .A2(\registers[19][13] ), .B1(n368), .B2(
        \registers[18][13] ), .ZN(n1937) );
  OAI221_X2 U1367 ( .B1(n659), .B2(n365), .C1(n627), .C2(n362), .A(n1938), 
        .ZN(n1935) );
  AOI22_X2 U1368 ( .A1(n359), .A2(\registers[23][13] ), .B1(n356), .B2(
        \registers[22][13] ), .ZN(n1938) );
  OAI221_X2 U1369 ( .B1(n851), .B2(n353), .C1(n819), .C2(n286), .A(n1939), 
        .ZN(n1934) );
  AOI22_X2 U1370 ( .A1(n283), .A2(\registers[25][13] ), .B1(n280), .B2(
        \registers[24][13] ), .ZN(n1939) );
  OAI221_X2 U1371 ( .B1(n979), .B2(n277), .C1(n947), .C2(n274), .A(n1940), 
        .ZN(n1933) );
  AOI22_X2 U1372 ( .A1(n271), .A2(\registers[29][13] ), .B1(n268), .B2(
        \registers[28][13] ), .ZN(n1940) );
  AOI211_X2 U1373 ( .C1(n265), .C2(\registers[1][13] ), .A(n1941), .B(n1942), 
        .ZN(n1931) );
  OAI22_X2 U1374 ( .A1(n51), .A2(n262), .B1(n83), .B2(n259), .ZN(n1942) );
  OAI221_X2 U1375 ( .B1(n147), .B2(n256), .C1(n115), .C2(n253), .A(n1943), 
        .ZN(n1941) );
  AOI22_X2 U1376 ( .A1(n250), .A2(\registers[7][13] ), .B1(n247), .B2(
        \registers[6][13] ), .ZN(n1943) );
  AOI221_X2 U1377 ( .B1(n244), .B2(\registers[13][13] ), .C1(n241), .C2(
        \registers[12][13] ), .A(n1944), .ZN(n1930) );
  OAI22_X2 U1378 ( .A1(n435), .A2(n238), .B1(n467), .B2(n235), .ZN(n1944) );
  AOI221_X2 U1379 ( .B1(n232), .B2(\registers[9][13] ), .C1(n229), .C2(
        \registers[8][13] ), .A(n1945), .ZN(n1929) );
  OAI22_X2 U1380 ( .A1(n307), .A2(n226), .B1(n339), .B2(n223), .ZN(n1945) );
  NAND4_X2 U1381 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(N333)
         );
  NOR4_X2 U1382 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1949)
         );
  OAI221_X2 U1383 ( .B1(n532), .B2(n377), .C1(n500), .C2(n374), .A(n1954), 
        .ZN(n1953) );
  AOI22_X2 U1384 ( .A1(n371), .A2(\registers[19][12] ), .B1(n368), .B2(
        \registers[18][12] ), .ZN(n1954) );
  OAI221_X2 U1385 ( .B1(n660), .B2(n365), .C1(n628), .C2(n362), .A(n1955), 
        .ZN(n1952) );
  AOI22_X2 U1386 ( .A1(n359), .A2(\registers[23][12] ), .B1(n356), .B2(
        \registers[22][12] ), .ZN(n1955) );
  OAI221_X2 U1387 ( .B1(n852), .B2(n353), .C1(n820), .C2(n286), .A(n1956), 
        .ZN(n1951) );
  AOI22_X2 U1388 ( .A1(n283), .A2(\registers[25][12] ), .B1(n280), .B2(
        \registers[24][12] ), .ZN(n1956) );
  OAI221_X2 U1389 ( .B1(n980), .B2(n277), .C1(n948), .C2(n274), .A(n1957), 
        .ZN(n1950) );
  AOI22_X2 U1390 ( .A1(n271), .A2(\registers[29][12] ), .B1(n268), .B2(
        \registers[28][12] ), .ZN(n1957) );
  AOI211_X2 U1391 ( .C1(n265), .C2(\registers[1][12] ), .A(n1958), .B(n1959), 
        .ZN(n1948) );
  OAI22_X2 U1392 ( .A1(n52), .A2(n262), .B1(n84), .B2(n259), .ZN(n1959) );
  OAI221_X2 U1393 ( .B1(n148), .B2(n256), .C1(n116), .C2(n253), .A(n1960), 
        .ZN(n1958) );
  AOI22_X2 U1394 ( .A1(n250), .A2(\registers[7][12] ), .B1(n247), .B2(
        \registers[6][12] ), .ZN(n1960) );
  AOI221_X2 U1395 ( .B1(n244), .B2(\registers[13][12] ), .C1(n241), .C2(
        \registers[12][12] ), .A(n1961), .ZN(n1947) );
  OAI22_X2 U1396 ( .A1(n436), .A2(n238), .B1(n468), .B2(n235), .ZN(n1961) );
  AOI221_X2 U1397 ( .B1(n232), .B2(\registers[9][12] ), .C1(n229), .C2(
        \registers[8][12] ), .A(n1962), .ZN(n1946) );
  OAI22_X2 U1398 ( .A1(n308), .A2(n226), .B1(n340), .B2(n223), .ZN(n1962) );
  NAND4_X2 U1399 ( .A1(n1963), .A2(n1964), .A3(n1965), .A4(n1966), .ZN(N332)
         );
  NOR4_X2 U1400 ( .A1(n1967), .A2(n1968), .A3(n1969), .A4(n1970), .ZN(n1966)
         );
  OAI221_X2 U1401 ( .B1(n533), .B2(n377), .C1(n501), .C2(n374), .A(n1971), 
        .ZN(n1970) );
  AOI22_X2 U1402 ( .A1(n371), .A2(\registers[19][11] ), .B1(n368), .B2(
        \registers[18][11] ), .ZN(n1971) );
  OAI221_X2 U1403 ( .B1(n661), .B2(n365), .C1(n629), .C2(n362), .A(n1972), 
        .ZN(n1969) );
  AOI22_X2 U1404 ( .A1(n359), .A2(\registers[23][11] ), .B1(n356), .B2(
        \registers[22][11] ), .ZN(n1972) );
  OAI221_X2 U1405 ( .B1(n853), .B2(n353), .C1(n821), .C2(n286), .A(n1973), 
        .ZN(n1968) );
  AOI22_X2 U1406 ( .A1(n283), .A2(\registers[25][11] ), .B1(n280), .B2(
        \registers[24][11] ), .ZN(n1973) );
  OAI221_X2 U1407 ( .B1(n981), .B2(n277), .C1(n949), .C2(n274), .A(n1974), 
        .ZN(n1967) );
  AOI22_X2 U1408 ( .A1(n271), .A2(\registers[29][11] ), .B1(n268), .B2(
        \registers[28][11] ), .ZN(n1974) );
  AOI211_X2 U1409 ( .C1(n265), .C2(\registers[1][11] ), .A(n1975), .B(n1976), 
        .ZN(n1965) );
  OAI22_X2 U1410 ( .A1(n53), .A2(n261), .B1(n85), .B2(n258), .ZN(n1976) );
  OAI221_X2 U1411 ( .B1(n149), .B2(n256), .C1(n117), .C2(n253), .A(n1977), 
        .ZN(n1975) );
  AOI22_X2 U1412 ( .A1(n250), .A2(\registers[7][11] ), .B1(n247), .B2(
        \registers[6][11] ), .ZN(n1977) );
  AOI221_X2 U1413 ( .B1(n244), .B2(\registers[13][11] ), .C1(n241), .C2(
        \registers[12][11] ), .A(n1978), .ZN(n1964) );
  OAI22_X2 U1414 ( .A1(n437), .A2(n237), .B1(n469), .B2(n234), .ZN(n1978) );
  AOI221_X2 U1415 ( .B1(n232), .B2(\registers[9][11] ), .C1(n229), .C2(
        \registers[8][11] ), .A(n1979), .ZN(n1963) );
  OAI22_X2 U1416 ( .A1(n309), .A2(n225), .B1(n341), .B2(n222), .ZN(n1979) );
  NAND4_X2 U1417 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .ZN(N331)
         );
  NOR4_X2 U1418 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(n1983)
         );
  OAI221_X2 U1419 ( .B1(n534), .B2(n376), .C1(n502), .C2(n373), .A(n1988), 
        .ZN(n1987) );
  AOI22_X2 U1420 ( .A1(n370), .A2(\registers[19][10] ), .B1(n367), .B2(
        \registers[18][10] ), .ZN(n1988) );
  OAI221_X2 U1421 ( .B1(n662), .B2(n364), .C1(n630), .C2(n361), .A(n1989), 
        .ZN(n1986) );
  AOI22_X2 U1422 ( .A1(n358), .A2(\registers[23][10] ), .B1(n355), .B2(
        \registers[22][10] ), .ZN(n1989) );
  OAI221_X2 U1423 ( .B1(n854), .B2(n288), .C1(n822), .C2(n285), .A(n1990), 
        .ZN(n1985) );
  AOI22_X2 U1424 ( .A1(n282), .A2(\registers[25][10] ), .B1(n279), .B2(
        \registers[24][10] ), .ZN(n1990) );
  OAI221_X2 U1425 ( .B1(n982), .B2(n276), .C1(n950), .C2(n273), .A(n1991), 
        .ZN(n1984) );
  AOI22_X2 U1426 ( .A1(n270), .A2(\registers[29][10] ), .B1(n267), .B2(
        \registers[28][10] ), .ZN(n1991) );
  AOI211_X2 U1427 ( .C1(n264), .C2(\registers[1][10] ), .A(n1992), .B(n1993), 
        .ZN(n1982) );
  OAI22_X2 U1428 ( .A1(n54), .A2(n261), .B1(n86), .B2(n258), .ZN(n1993) );
  OAI221_X2 U1429 ( .B1(n150), .B2(n255), .C1(n118), .C2(n252), .A(n1994), 
        .ZN(n1992) );
  AOI22_X2 U1430 ( .A1(n249), .A2(\registers[7][10] ), .B1(n246), .B2(
        \registers[6][10] ), .ZN(n1994) );
  AOI221_X2 U1431 ( .B1(n243), .B2(\registers[13][10] ), .C1(n240), .C2(
        \registers[12][10] ), .A(n1995), .ZN(n1981) );
  OAI22_X2 U1432 ( .A1(n438), .A2(n237), .B1(n470), .B2(n234), .ZN(n1995) );
  AOI221_X2 U1433 ( .B1(n231), .B2(\registers[9][10] ), .C1(n228), .C2(
        \registers[8][10] ), .A(n1996), .ZN(n1980) );
  OAI22_X2 U1434 ( .A1(n310), .A2(n225), .B1(n342), .B2(n222), .ZN(n1996) );
  NAND4_X2 U1435 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(N330)
         );
  NOR4_X2 U1436 ( .A1(n2001), .A2(n2002), .A3(n2003), .A4(n2004), .ZN(n2000)
         );
  OAI221_X2 U1437 ( .B1(n535), .B2(n376), .C1(n503), .C2(n373), .A(n2005), 
        .ZN(n2004) );
  AOI22_X2 U1438 ( .A1(n370), .A2(\registers[19][9] ), .B1(n367), .B2(
        \registers[18][9] ), .ZN(n2005) );
  OAI221_X2 U1439 ( .B1(n663), .B2(n364), .C1(n631), .C2(n361), .A(n2006), 
        .ZN(n2003) );
  AOI22_X2 U1440 ( .A1(n358), .A2(\registers[23][9] ), .B1(n355), .B2(
        \registers[22][9] ), .ZN(n2006) );
  OAI221_X2 U1441 ( .B1(n855), .B2(n288), .C1(n823), .C2(n285), .A(n2007), 
        .ZN(n2002) );
  AOI22_X2 U1442 ( .A1(n282), .A2(\registers[25][9] ), .B1(n279), .B2(
        \registers[24][9] ), .ZN(n2007) );
  OAI221_X2 U1443 ( .B1(n983), .B2(n276), .C1(n951), .C2(n273), .A(n2008), 
        .ZN(n2001) );
  AOI22_X2 U1444 ( .A1(n270), .A2(\registers[29][9] ), .B1(n267), .B2(
        \registers[28][9] ), .ZN(n2008) );
  AOI211_X2 U1445 ( .C1(n264), .C2(\registers[1][9] ), .A(n2009), .B(n2010), 
        .ZN(n1999) );
  OAI22_X2 U1446 ( .A1(n55), .A2(n261), .B1(n87), .B2(n258), .ZN(n2010) );
  OAI221_X2 U1447 ( .B1(n151), .B2(n255), .C1(n119), .C2(n252), .A(n2011), 
        .ZN(n2009) );
  AOI22_X2 U1448 ( .A1(n249), .A2(\registers[7][9] ), .B1(n246), .B2(
        \registers[6][9] ), .ZN(n2011) );
  AOI221_X2 U1449 ( .B1(n243), .B2(\registers[13][9] ), .C1(n240), .C2(
        \registers[12][9] ), .A(n2012), .ZN(n1998) );
  OAI22_X2 U1450 ( .A1(n439), .A2(n237), .B1(n471), .B2(n234), .ZN(n2012) );
  AOI221_X2 U1451 ( .B1(n231), .B2(\registers[9][9] ), .C1(n228), .C2(
        \registers[8][9] ), .A(n2013), .ZN(n1997) );
  OAI22_X2 U1452 ( .A1(n311), .A2(n225), .B1(n343), .B2(n222), .ZN(n2013) );
  NAND4_X2 U1453 ( .A1(n2014), .A2(n2015), .A3(n2016), .A4(n2017), .ZN(N329)
         );
  NOR4_X2 U1454 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2017)
         );
  OAI221_X2 U1455 ( .B1(n536), .B2(n376), .C1(n504), .C2(n373), .A(n2022), 
        .ZN(n2021) );
  AOI22_X2 U1456 ( .A1(n370), .A2(\registers[19][8] ), .B1(n367), .B2(
        \registers[18][8] ), .ZN(n2022) );
  OAI221_X2 U1457 ( .B1(n664), .B2(n364), .C1(n632), .C2(n361), .A(n2023), 
        .ZN(n2020) );
  AOI22_X2 U1458 ( .A1(n358), .A2(\registers[23][8] ), .B1(n355), .B2(
        \registers[22][8] ), .ZN(n2023) );
  OAI221_X2 U1459 ( .B1(n856), .B2(n288), .C1(n824), .C2(n285), .A(n2024), 
        .ZN(n2019) );
  AOI22_X2 U1460 ( .A1(n282), .A2(\registers[25][8] ), .B1(n279), .B2(
        \registers[24][8] ), .ZN(n2024) );
  OAI221_X2 U1461 ( .B1(n984), .B2(n276), .C1(n952), .C2(n273), .A(n2025), 
        .ZN(n2018) );
  AOI22_X2 U1462 ( .A1(n270), .A2(\registers[29][8] ), .B1(n267), .B2(
        \registers[28][8] ), .ZN(n2025) );
  AOI211_X2 U1463 ( .C1(n264), .C2(\registers[1][8] ), .A(n2026), .B(n2027), 
        .ZN(n2016) );
  OAI22_X2 U1464 ( .A1(n56), .A2(n261), .B1(n88), .B2(n258), .ZN(n2027) );
  OAI221_X2 U1465 ( .B1(n152), .B2(n255), .C1(n120), .C2(n252), .A(n2028), 
        .ZN(n2026) );
  AOI22_X2 U1466 ( .A1(n249), .A2(\registers[7][8] ), .B1(n246), .B2(
        \registers[6][8] ), .ZN(n2028) );
  AOI221_X2 U1467 ( .B1(n243), .B2(\registers[13][8] ), .C1(n240), .C2(
        \registers[12][8] ), .A(n2029), .ZN(n2015) );
  OAI22_X2 U1468 ( .A1(n440), .A2(n237), .B1(n472), .B2(n234), .ZN(n2029) );
  AOI221_X2 U1469 ( .B1(n231), .B2(\registers[9][8] ), .C1(n228), .C2(
        \registers[8][8] ), .A(n2030), .ZN(n2014) );
  OAI22_X2 U1470 ( .A1(n312), .A2(n225), .B1(n344), .B2(n222), .ZN(n2030) );
  NAND4_X2 U1471 ( .A1(n2031), .A2(n2032), .A3(n2033), .A4(n2034), .ZN(N328)
         );
  NOR4_X2 U1472 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .ZN(n2034)
         );
  OAI221_X2 U1473 ( .B1(n537), .B2(n376), .C1(n505), .C2(n373), .A(n2039), 
        .ZN(n2038) );
  AOI22_X2 U1474 ( .A1(n370), .A2(\registers[19][7] ), .B1(n367), .B2(
        \registers[18][7] ), .ZN(n2039) );
  OAI221_X2 U1475 ( .B1(n665), .B2(n364), .C1(n633), .C2(n361), .A(n2040), 
        .ZN(n2037) );
  AOI22_X2 U1476 ( .A1(n358), .A2(\registers[23][7] ), .B1(n355), .B2(
        \registers[22][7] ), .ZN(n2040) );
  OAI221_X2 U1477 ( .B1(n857), .B2(n288), .C1(n825), .C2(n285), .A(n2041), 
        .ZN(n2036) );
  AOI22_X2 U1478 ( .A1(n282), .A2(\registers[25][7] ), .B1(n279), .B2(
        \registers[24][7] ), .ZN(n2041) );
  OAI221_X2 U1479 ( .B1(n985), .B2(n276), .C1(n953), .C2(n273), .A(n2042), 
        .ZN(n2035) );
  AOI22_X2 U1480 ( .A1(n270), .A2(\registers[29][7] ), .B1(n267), .B2(
        \registers[28][7] ), .ZN(n2042) );
  AOI211_X2 U1481 ( .C1(n264), .C2(\registers[1][7] ), .A(n2043), .B(n2044), 
        .ZN(n2033) );
  OAI22_X2 U1482 ( .A1(n57), .A2(n261), .B1(n89), .B2(n258), .ZN(n2044) );
  OAI221_X2 U1483 ( .B1(n153), .B2(n255), .C1(n121), .C2(n252), .A(n2045), 
        .ZN(n2043) );
  AOI22_X2 U1484 ( .A1(n249), .A2(\registers[7][7] ), .B1(n246), .B2(
        \registers[6][7] ), .ZN(n2045) );
  AOI221_X2 U1485 ( .B1(n243), .B2(\registers[13][7] ), .C1(n240), .C2(
        \registers[12][7] ), .A(n2046), .ZN(n2032) );
  OAI22_X2 U1486 ( .A1(n441), .A2(n237), .B1(n473), .B2(n234), .ZN(n2046) );
  AOI221_X2 U1487 ( .B1(n231), .B2(\registers[9][7] ), .C1(n228), .C2(
        \registers[8][7] ), .A(n2047), .ZN(n2031) );
  OAI22_X2 U1488 ( .A1(n313), .A2(n225), .B1(n345), .B2(n222), .ZN(n2047) );
  NAND4_X2 U1489 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(N327)
         );
  NOR4_X2 U1490 ( .A1(n2052), .A2(n2053), .A3(n2054), .A4(n2055), .ZN(n2051)
         );
  OAI221_X2 U1491 ( .B1(n538), .B2(n376), .C1(n506), .C2(n373), .A(n2056), 
        .ZN(n2055) );
  AOI22_X2 U1492 ( .A1(n370), .A2(\registers[19][6] ), .B1(n367), .B2(
        \registers[18][6] ), .ZN(n2056) );
  OAI221_X2 U1493 ( .B1(n666), .B2(n364), .C1(n634), .C2(n361), .A(n2057), 
        .ZN(n2054) );
  AOI22_X2 U1494 ( .A1(n358), .A2(\registers[23][6] ), .B1(n355), .B2(
        \registers[22][6] ), .ZN(n2057) );
  OAI221_X2 U1495 ( .B1(n858), .B2(n288), .C1(n826), .C2(n285), .A(n2058), 
        .ZN(n2053) );
  AOI22_X2 U1496 ( .A1(n282), .A2(\registers[25][6] ), .B1(n279), .B2(
        \registers[24][6] ), .ZN(n2058) );
  OAI221_X2 U1497 ( .B1(n986), .B2(n276), .C1(n954), .C2(n273), .A(n2059), 
        .ZN(n2052) );
  AOI22_X2 U1498 ( .A1(n270), .A2(\registers[29][6] ), .B1(n267), .B2(
        \registers[28][6] ), .ZN(n2059) );
  AOI211_X2 U1499 ( .C1(n264), .C2(\registers[1][6] ), .A(n2060), .B(n2061), 
        .ZN(n2050) );
  OAI22_X2 U1500 ( .A1(n58), .A2(n261), .B1(n90), .B2(n258), .ZN(n2061) );
  OAI221_X2 U1501 ( .B1(n154), .B2(n255), .C1(n122), .C2(n252), .A(n2062), 
        .ZN(n2060) );
  AOI22_X2 U1502 ( .A1(n249), .A2(\registers[7][6] ), .B1(n246), .B2(
        \registers[6][6] ), .ZN(n2062) );
  AOI221_X2 U1503 ( .B1(n243), .B2(\registers[13][6] ), .C1(n240), .C2(
        \registers[12][6] ), .A(n2063), .ZN(n2049) );
  OAI22_X2 U1504 ( .A1(n442), .A2(n237), .B1(n474), .B2(n234), .ZN(n2063) );
  AOI221_X2 U1505 ( .B1(n231), .B2(\registers[9][6] ), .C1(n228), .C2(
        \registers[8][6] ), .A(n2064), .ZN(n2048) );
  OAI22_X2 U1506 ( .A1(n314), .A2(n225), .B1(n346), .B2(n222), .ZN(n2064) );
  NAND4_X2 U1507 ( .A1(n2065), .A2(n2066), .A3(n2067), .A4(n2068), .ZN(N326)
         );
  NOR4_X2 U1508 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2068)
         );
  OAI221_X2 U1509 ( .B1(n539), .B2(n376), .C1(n507), .C2(n373), .A(n2073), 
        .ZN(n2072) );
  AOI22_X2 U1510 ( .A1(n370), .A2(\registers[19][5] ), .B1(n367), .B2(
        \registers[18][5] ), .ZN(n2073) );
  OAI221_X2 U1511 ( .B1(n667), .B2(n364), .C1(n635), .C2(n361), .A(n2074), 
        .ZN(n2071) );
  AOI22_X2 U1512 ( .A1(n358), .A2(\registers[23][5] ), .B1(n355), .B2(
        \registers[22][5] ), .ZN(n2074) );
  OAI221_X2 U1513 ( .B1(n859), .B2(n288), .C1(n827), .C2(n285), .A(n2075), 
        .ZN(n2070) );
  AOI22_X2 U1514 ( .A1(n282), .A2(\registers[25][5] ), .B1(n279), .B2(
        \registers[24][5] ), .ZN(n2075) );
  OAI221_X2 U1515 ( .B1(n987), .B2(n276), .C1(n955), .C2(n273), .A(n2076), 
        .ZN(n2069) );
  AOI22_X2 U1516 ( .A1(n270), .A2(\registers[29][5] ), .B1(n267), .B2(
        \registers[28][5] ), .ZN(n2076) );
  AOI211_X2 U1517 ( .C1(n264), .C2(\registers[1][5] ), .A(n2077), .B(n2078), 
        .ZN(n2067) );
  OAI22_X2 U1518 ( .A1(n59), .A2(n261), .B1(n91), .B2(n258), .ZN(n2078) );
  OAI221_X2 U1519 ( .B1(n155), .B2(n255), .C1(n123), .C2(n252), .A(n2079), 
        .ZN(n2077) );
  AOI22_X2 U1520 ( .A1(n249), .A2(\registers[7][5] ), .B1(n246), .B2(
        \registers[6][5] ), .ZN(n2079) );
  AOI221_X2 U1521 ( .B1(n243), .B2(\registers[13][5] ), .C1(n240), .C2(
        \registers[12][5] ), .A(n2080), .ZN(n2066) );
  OAI22_X2 U1522 ( .A1(n443), .A2(n237), .B1(n475), .B2(n234), .ZN(n2080) );
  AOI221_X2 U1523 ( .B1(n231), .B2(\registers[9][5] ), .C1(n228), .C2(
        \registers[8][5] ), .A(n2081), .ZN(n2065) );
  OAI22_X2 U1524 ( .A1(n315), .A2(n225), .B1(n347), .B2(n222), .ZN(n2081) );
  NAND4_X2 U1525 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(N325)
         );
  NOR4_X2 U1526 ( .A1(n2086), .A2(n2087), .A3(n2088), .A4(n2089), .ZN(n2085)
         );
  OAI221_X2 U1527 ( .B1(n540), .B2(n376), .C1(n508), .C2(n373), .A(n2090), 
        .ZN(n2089) );
  AOI22_X2 U1528 ( .A1(n370), .A2(\registers[19][4] ), .B1(n367), .B2(
        \registers[18][4] ), .ZN(n2090) );
  OAI221_X2 U1529 ( .B1(n668), .B2(n364), .C1(n636), .C2(n361), .A(n2091), 
        .ZN(n2088) );
  AOI22_X2 U1530 ( .A1(n358), .A2(\registers[23][4] ), .B1(n355), .B2(
        \registers[22][4] ), .ZN(n2091) );
  OAI221_X2 U1531 ( .B1(n860), .B2(n288), .C1(n828), .C2(n285), .A(n2092), 
        .ZN(n2087) );
  AOI22_X2 U1532 ( .A1(n282), .A2(\registers[25][4] ), .B1(n279), .B2(
        \registers[24][4] ), .ZN(n2092) );
  OAI221_X2 U1533 ( .B1(n988), .B2(n276), .C1(n956), .C2(n273), .A(n2093), 
        .ZN(n2086) );
  AOI22_X2 U1534 ( .A1(n270), .A2(\registers[29][4] ), .B1(n267), .B2(
        \registers[28][4] ), .ZN(n2093) );
  AOI211_X2 U1535 ( .C1(n264), .C2(\registers[1][4] ), .A(n2094), .B(n2095), 
        .ZN(n2084) );
  OAI22_X2 U1536 ( .A1(n60), .A2(n261), .B1(n92), .B2(n258), .ZN(n2095) );
  OAI221_X2 U1537 ( .B1(n156), .B2(n255), .C1(n124), .C2(n252), .A(n2096), 
        .ZN(n2094) );
  AOI22_X2 U1538 ( .A1(n249), .A2(\registers[7][4] ), .B1(n246), .B2(
        \registers[6][4] ), .ZN(n2096) );
  AOI221_X2 U1539 ( .B1(n243), .B2(\registers[13][4] ), .C1(n240), .C2(
        \registers[12][4] ), .A(n2097), .ZN(n2083) );
  OAI22_X2 U1540 ( .A1(n444), .A2(n237), .B1(n476), .B2(n234), .ZN(n2097) );
  AOI221_X2 U1541 ( .B1(n231), .B2(\registers[9][4] ), .C1(n228), .C2(
        \registers[8][4] ), .A(n2098), .ZN(n2082) );
  OAI22_X2 U1542 ( .A1(n316), .A2(n225), .B1(n348), .B2(n222), .ZN(n2098) );
  NAND4_X2 U1543 ( .A1(n2099), .A2(n2100), .A3(n2101), .A4(n2102), .ZN(N324)
         );
  NOR4_X2 U1544 ( .A1(n2103), .A2(n2104), .A3(n2105), .A4(n2106), .ZN(n2102)
         );
  OAI221_X2 U1545 ( .B1(n541), .B2(n376), .C1(n509), .C2(n373), .A(n2107), 
        .ZN(n2106) );
  AOI22_X2 U1546 ( .A1(n370), .A2(\registers[19][3] ), .B1(n367), .B2(
        \registers[18][3] ), .ZN(n2107) );
  OAI221_X2 U1547 ( .B1(n669), .B2(n364), .C1(n637), .C2(n361), .A(n2108), 
        .ZN(n2105) );
  AOI22_X2 U1548 ( .A1(n358), .A2(\registers[23][3] ), .B1(n355), .B2(
        \registers[22][3] ), .ZN(n2108) );
  OAI221_X2 U1549 ( .B1(n861), .B2(n288), .C1(n829), .C2(n285), .A(n2109), 
        .ZN(n2104) );
  AOI22_X2 U1550 ( .A1(n282), .A2(\registers[25][3] ), .B1(n279), .B2(
        \registers[24][3] ), .ZN(n2109) );
  OAI221_X2 U1551 ( .B1(n989), .B2(n276), .C1(n957), .C2(n273), .A(n2110), 
        .ZN(n2103) );
  AOI22_X2 U1552 ( .A1(n270), .A2(\registers[29][3] ), .B1(n267), .B2(
        \registers[28][3] ), .ZN(n2110) );
  AOI211_X2 U1553 ( .C1(n264), .C2(\registers[1][3] ), .A(n2111), .B(n2112), 
        .ZN(n2101) );
  OAI22_X2 U1554 ( .A1(n61), .A2(n261), .B1(n93), .B2(n258), .ZN(n2112) );
  OAI221_X2 U1555 ( .B1(n157), .B2(n255), .C1(n125), .C2(n252), .A(n2113), 
        .ZN(n2111) );
  AOI22_X2 U1556 ( .A1(n249), .A2(\registers[7][3] ), .B1(n246), .B2(
        \registers[6][3] ), .ZN(n2113) );
  AOI221_X2 U1557 ( .B1(n243), .B2(\registers[13][3] ), .C1(n240), .C2(
        \registers[12][3] ), .A(n2114), .ZN(n2100) );
  OAI22_X2 U1558 ( .A1(n445), .A2(n237), .B1(n477), .B2(n234), .ZN(n2114) );
  AOI221_X2 U1559 ( .B1(n231), .B2(\registers[9][3] ), .C1(n228), .C2(
        \registers[8][3] ), .A(n2115), .ZN(n2099) );
  OAI22_X2 U1560 ( .A1(n317), .A2(n225), .B1(n349), .B2(n222), .ZN(n2115) );
  NAND4_X2 U1561 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(N323)
         );
  NOR4_X2 U1562 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2119)
         );
  OAI221_X2 U1563 ( .B1(n542), .B2(n376), .C1(n510), .C2(n373), .A(n2124), 
        .ZN(n2123) );
  AOI22_X2 U1564 ( .A1(n370), .A2(\registers[19][2] ), .B1(n367), .B2(
        \registers[18][2] ), .ZN(n2124) );
  OAI221_X2 U1565 ( .B1(n670), .B2(n364), .C1(n638), .C2(n361), .A(n2125), 
        .ZN(n2122) );
  AOI22_X2 U1566 ( .A1(n358), .A2(\registers[23][2] ), .B1(n355), .B2(
        \registers[22][2] ), .ZN(n2125) );
  OAI221_X2 U1567 ( .B1(n862), .B2(n288), .C1(n830), .C2(n285), .A(n2126), 
        .ZN(n2121) );
  AOI22_X2 U1568 ( .A1(n282), .A2(\registers[25][2] ), .B1(n279), .B2(
        \registers[24][2] ), .ZN(n2126) );
  OAI221_X2 U1569 ( .B1(n990), .B2(n276), .C1(n958), .C2(n273), .A(n2127), 
        .ZN(n2120) );
  AOI22_X2 U1570 ( .A1(n270), .A2(\registers[29][2] ), .B1(n267), .B2(
        \registers[28][2] ), .ZN(n2127) );
  AOI211_X2 U1571 ( .C1(n264), .C2(\registers[1][2] ), .A(n2128), .B(n2129), 
        .ZN(n2118) );
  OAI22_X2 U1572 ( .A1(n62), .A2(n261), .B1(n94), .B2(n258), .ZN(n2129) );
  OAI221_X2 U1573 ( .B1(n158), .B2(n255), .C1(n126), .C2(n252), .A(n2130), 
        .ZN(n2128) );
  AOI22_X2 U1574 ( .A1(n249), .A2(\registers[7][2] ), .B1(n246), .B2(
        \registers[6][2] ), .ZN(n2130) );
  AOI221_X2 U1575 ( .B1(n243), .B2(\registers[13][2] ), .C1(n240), .C2(
        \registers[12][2] ), .A(n2131), .ZN(n2117) );
  OAI22_X2 U1576 ( .A1(n446), .A2(n237), .B1(n478), .B2(n234), .ZN(n2131) );
  AOI221_X2 U1577 ( .B1(n231), .B2(\registers[9][2] ), .C1(n228), .C2(
        \registers[8][2] ), .A(n2132), .ZN(n2116) );
  OAI22_X2 U1578 ( .A1(n318), .A2(n225), .B1(n350), .B2(n222), .ZN(n2132) );
  NAND4_X2 U1579 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(N322)
         );
  NOR4_X2 U1580 ( .A1(n2137), .A2(n2138), .A3(n2139), .A4(n2140), .ZN(n2136)
         );
  OAI221_X2 U1581 ( .B1(n543), .B2(n376), .C1(n511), .C2(n373), .A(n2141), 
        .ZN(n2140) );
  AOI22_X2 U1582 ( .A1(n370), .A2(\registers[19][1] ), .B1(n367), .B2(
        \registers[18][1] ), .ZN(n2141) );
  OAI221_X2 U1583 ( .B1(n671), .B2(n364), .C1(n639), .C2(n361), .A(n2142), 
        .ZN(n2139) );
  AOI22_X2 U1584 ( .A1(n358), .A2(\registers[23][1] ), .B1(n355), .B2(
        \registers[22][1] ), .ZN(n2142) );
  OAI221_X2 U1585 ( .B1(n863), .B2(n288), .C1(n831), .C2(n285), .A(n2143), 
        .ZN(n2138) );
  AOI22_X2 U1586 ( .A1(n282), .A2(\registers[25][1] ), .B1(n279), .B2(
        \registers[24][1] ), .ZN(n2143) );
  OAI221_X2 U1587 ( .B1(n991), .B2(n276), .C1(n959), .C2(n273), .A(n2144), 
        .ZN(n2137) );
  AOI22_X2 U1588 ( .A1(n270), .A2(\registers[29][1] ), .B1(n267), .B2(
        \registers[28][1] ), .ZN(n2144) );
  AOI211_X2 U1589 ( .C1(n264), .C2(\registers[1][1] ), .A(n2145), .B(n2146), 
        .ZN(n2135) );
  OAI22_X2 U1590 ( .A1(n63), .A2(n261), .B1(n95), .B2(n258), .ZN(n2146) );
  OAI221_X2 U1591 ( .B1(n159), .B2(n255), .C1(n127), .C2(n252), .A(n2147), 
        .ZN(n2145) );
  AOI22_X2 U1592 ( .A1(n249), .A2(\registers[7][1] ), .B1(n246), .B2(
        \registers[6][1] ), .ZN(n2147) );
  AOI221_X2 U1593 ( .B1(n243), .B2(\registers[13][1] ), .C1(n240), .C2(
        \registers[12][1] ), .A(n2148), .ZN(n2134) );
  OAI22_X2 U1594 ( .A1(n447), .A2(n237), .B1(n479), .B2(n234), .ZN(n2148) );
  AOI221_X2 U1595 ( .B1(n231), .B2(\registers[9][1] ), .C1(n228), .C2(
        \registers[8][1] ), .A(n2149), .ZN(n2133) );
  OAI22_X2 U1596 ( .A1(n319), .A2(n225), .B1(n351), .B2(n222), .ZN(n2149) );
  NAND4_X2 U1597 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .ZN(N321)
         );
  NOR4_X2 U1598 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2153)
         );
  OAI221_X2 U1599 ( .B1(n544), .B2(n376), .C1(n512), .C2(n373), .A(n2158), 
        .ZN(n2157) );
  AOI22_X2 U1600 ( .A1(n370), .A2(\registers[19][0] ), .B1(n367), .B2(
        \registers[18][0] ), .ZN(n2158) );
  AND2_X2 U1601 ( .A1(n2159), .A2(n2160), .ZN(n1604) );
  AND2_X2 U1602 ( .A1(n2161), .A2(n2160), .ZN(n1603) );
  NAND2_X2 U1603 ( .A1(n2159), .A2(n2162), .ZN(n1601) );
  NAND2_X2 U1604 ( .A1(n2161), .A2(n2162), .ZN(n1600) );
  OAI221_X2 U1605 ( .B1(n672), .B2(n364), .C1(n640), .C2(n361), .A(n2163), 
        .ZN(n2156) );
  AOI22_X2 U1606 ( .A1(n358), .A2(\registers[23][0] ), .B1(n355), .B2(
        \registers[22][0] ), .ZN(n2163) );
  AND2_X2 U1607 ( .A1(n2159), .A2(n2164), .ZN(n1609) );
  AND2_X2 U1608 ( .A1(n2161), .A2(n2164), .ZN(n1608) );
  NAND2_X2 U1609 ( .A1(n2159), .A2(n2165), .ZN(n1606) );
  AND2_X2 U1610 ( .A1(n2166), .A2(n3858), .ZN(n2159) );
  NAND2_X2 U1611 ( .A1(n2161), .A2(n2165), .ZN(n1605) );
  AND2_X2 U1612 ( .A1(n2166), .A2(ADD_RD2[0]), .ZN(n2161) );
  AND2_X2 U1613 ( .A1(ADD_RD2[4]), .A2(n3856), .ZN(n2166) );
  OAI221_X2 U1614 ( .B1(n864), .B2(n288), .C1(n832), .C2(n285), .A(n2167), 
        .ZN(n2155) );
  AOI22_X2 U1615 ( .A1(n282), .A2(\registers[25][0] ), .B1(n279), .B2(
        \registers[24][0] ), .ZN(n2167) );
  AND2_X2 U1616 ( .A1(n2162), .A2(n2168), .ZN(n1614) );
  AND2_X2 U1617 ( .A1(n2162), .A2(n2169), .ZN(n1613) );
  NAND2_X2 U1618 ( .A1(n2160), .A2(n2168), .ZN(n1611) );
  NAND2_X2 U1619 ( .A1(n2160), .A2(n2169), .ZN(n1610) );
  OAI221_X2 U1620 ( .B1(n992), .B2(n276), .C1(n960), .C2(n273), .A(n2170), 
        .ZN(n2154) );
  AOI22_X2 U1621 ( .A1(n270), .A2(\registers[29][0] ), .B1(n267), .B2(
        \registers[28][0] ), .ZN(n2170) );
  AND2_X2 U1622 ( .A1(n2165), .A2(n2168), .ZN(n1619) );
  AND2_X2 U1623 ( .A1(n2165), .A2(n2169), .ZN(n1618) );
  NAND2_X2 U1624 ( .A1(n2168), .A2(n2164), .ZN(n1616) );
  AND2_X2 U1625 ( .A1(n2171), .A2(n3858), .ZN(n2168) );
  NAND2_X2 U1626 ( .A1(n2164), .A2(n2169), .ZN(n1615) );
  AND2_X2 U1627 ( .A1(ADD_RD2[0]), .A2(n2171), .ZN(n2169) );
  AND2_X2 U1628 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n2171) );
  AOI211_X2 U1629 ( .C1(n264), .C2(\registers[1][0] ), .A(n2172), .B(n2173), 
        .ZN(n2152) );
  OAI22_X2 U1630 ( .A1(n64), .A2(n261), .B1(n96), .B2(n258), .ZN(n2173) );
  NAND2_X2 U1631 ( .A1(n2174), .A2(n2160), .ZN(n1624) );
  NAND2_X2 U1632 ( .A1(n2175), .A2(n2160), .ZN(n1623) );
  OAI221_X2 U1633 ( .B1(n160), .B2(n255), .C1(n128), .C2(n252), .A(n2176), 
        .ZN(n2172) );
  AOI22_X2 U1634 ( .A1(n249), .A2(\registers[7][0] ), .B1(n246), .B2(
        \registers[6][0] ), .ZN(n2176) );
  AND2_X2 U1635 ( .A1(n2175), .A2(n2164), .ZN(n1629) );
  AND2_X2 U1636 ( .A1(n2174), .A2(n2164), .ZN(n1628) );
  NAND2_X2 U1637 ( .A1(n2175), .A2(n2165), .ZN(n1626) );
  AND2_X2 U1638 ( .A1(n2177), .A2(n3858), .ZN(n2175) );
  NAND2_X2 U1639 ( .A1(n2174), .A2(n2165), .ZN(n1625) );
  AND2_X2 U1640 ( .A1(n2174), .A2(n2162), .ZN(n1620) );
  AND2_X2 U1641 ( .A1(n2177), .A2(ADD_RD2[0]), .ZN(n2174) );
  NOR2_X2 U1642 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n2177) );
  AOI221_X2 U1643 ( .B1(n243), .B2(\registers[13][0] ), .C1(n240), .C2(
        \registers[12][0] ), .A(n2178), .ZN(n2151) );
  OAI22_X2 U1644 ( .A1(n448), .A2(n237), .B1(n480), .B2(n234), .ZN(n2178) );
  NAND2_X2 U1645 ( .A1(n2179), .A2(n2164), .ZN(n1634) );
  NAND2_X2 U1646 ( .A1(n2180), .A2(n2164), .ZN(n1633) );
  AND2_X2 U1647 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n2164) );
  AND2_X2 U1648 ( .A1(n2180), .A2(n2165), .ZN(n1631) );
  AND2_X2 U1649 ( .A1(n2179), .A2(n2165), .ZN(n1630) );
  AND2_X2 U1650 ( .A1(ADD_RD2[2]), .A2(n3857), .ZN(n2165) );
  AOI221_X2 U1651 ( .B1(n231), .B2(\registers[9][0] ), .C1(n228), .C2(
        \registers[8][0] ), .A(n2181), .ZN(n2150) );
  OAI22_X2 U1652 ( .A1(n320), .A2(n225), .B1(n352), .B2(n222), .ZN(n2181) );
  NAND2_X2 U1653 ( .A1(n2179), .A2(n2160), .ZN(n1639) );
  NAND2_X2 U1654 ( .A1(n2180), .A2(n2160), .ZN(n1638) );
  NOR2_X2 U1655 ( .A1(n3857), .A2(ADD_RD2[2]), .ZN(n2160) );
  AND2_X2 U1656 ( .A1(n2180), .A2(n2162), .ZN(n1636) );
  AND2_X2 U1657 ( .A1(n2182), .A2(n3858), .ZN(n2180) );
  AND2_X2 U1658 ( .A1(n2179), .A2(n2162), .ZN(n1635) );
  NOR2_X2 U1659 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n2162) );
  AND2_X2 U1660 ( .A1(n2182), .A2(ADD_RD2[0]), .ZN(n2179) );
  NOR2_X2 U1661 ( .A1(n3856), .A2(ADD_RD2[4]), .ZN(n2182) );
  AND2_X2 U1662 ( .A1(RD2), .A2(ENABLE), .ZN(N218) );
  NAND4_X2 U1663 ( .A1(n2183), .A2(n2184), .A3(n2185), .A4(n2186), .ZN(N217)
         );
  NOR4_X2 U1664 ( .A1(n2187), .A2(n2188), .A3(n2189), .A4(n2190), .ZN(n2186)
         );
  OAI221_X2 U1665 ( .B1(n513), .B2(n221), .C1(n481), .C2(n218), .A(n2193), 
        .ZN(n2190) );
  AOI22_X2 U1666 ( .A1(n215), .A2(\registers[19][31] ), .B1(n212), .B2(
        \registers[18][31] ), .ZN(n2193) );
  OAI221_X2 U1667 ( .B1(n641), .B2(n209), .C1(n609), .C2(n206), .A(n2198), 
        .ZN(n2189) );
  AOI22_X2 U1668 ( .A1(n203), .A2(\registers[23][31] ), .B1(n200), .B2(
        \registers[22][31] ), .ZN(n2198) );
  OAI221_X2 U1669 ( .B1(n833), .B2(n197), .C1(n801), .C2(n194), .A(n2203), 
        .ZN(n2188) );
  AOI22_X2 U1670 ( .A1(n191), .A2(\registers[25][31] ), .B1(n188), .B2(
        \registers[24][31] ), .ZN(n2203) );
  OAI221_X2 U1671 ( .B1(n961), .B2(n185), .C1(n929), .C2(n182), .A(n2208), 
        .ZN(n2187) );
  AOI22_X2 U1672 ( .A1(n179), .A2(\registers[29][31] ), .B1(n176), .B2(
        \registers[28][31] ), .ZN(n2208) );
  AOI211_X2 U1673 ( .C1(n173), .C2(\registers[1][31] ), .A(n2212), .B(n2213), 
        .ZN(n2185) );
  OAI22_X2 U1674 ( .A1(n33), .A2(n170), .B1(n65), .B2(n167), .ZN(n2213) );
  OAI221_X2 U1675 ( .B1(n129), .B2(n164), .C1(n97), .C2(n161), .A(n2218), .ZN(
        n2212) );
  AOI22_X2 U1676 ( .A1(n30), .A2(\registers[7][31] ), .B1(n27), .B2(
        \registers[6][31] ), .ZN(n2218) );
  AOI221_X2 U1677 ( .B1(n24), .B2(\registers[13][31] ), .C1(n21), .C2(
        \registers[12][31] ), .A(n2223), .ZN(n2184) );
  OAI22_X2 U1678 ( .A1(n417), .A2(n18), .B1(n449), .B2(n15), .ZN(n2223) );
  AOI221_X2 U1679 ( .B1(n12), .B2(\registers[9][31] ), .C1(n9), .C2(
        \registers[8][31] ), .A(n2228), .ZN(n2183) );
  OAI22_X2 U1680 ( .A1(n289), .A2(n6), .B1(n321), .B2(n3), .ZN(n2228) );
  NAND4_X2 U1681 ( .A1(n2231), .A2(n2232), .A3(n2233), .A4(n2234), .ZN(N216)
         );
  NOR4_X2 U1682 ( .A1(n2235), .A2(n2236), .A3(n2237), .A4(n2238), .ZN(n2234)
         );
  OAI221_X2 U1683 ( .B1(n514), .B2(n221), .C1(n482), .C2(n218), .A(n2239), 
        .ZN(n2238) );
  AOI22_X2 U1684 ( .A1(n215), .A2(\registers[19][30] ), .B1(n212), .B2(
        \registers[18][30] ), .ZN(n2239) );
  OAI221_X2 U1685 ( .B1(n642), .B2(n209), .C1(n610), .C2(n206), .A(n2240), 
        .ZN(n2237) );
  AOI22_X2 U1686 ( .A1(n203), .A2(\registers[23][30] ), .B1(n200), .B2(
        \registers[22][30] ), .ZN(n2240) );
  OAI221_X2 U1687 ( .B1(n834), .B2(n197), .C1(n802), .C2(n194), .A(n2241), 
        .ZN(n2236) );
  AOI22_X2 U1688 ( .A1(n191), .A2(\registers[25][30] ), .B1(n188), .B2(
        \registers[24][30] ), .ZN(n2241) );
  OAI221_X2 U1689 ( .B1(n962), .B2(n185), .C1(n930), .C2(n182), .A(n2242), 
        .ZN(n2235) );
  AOI22_X2 U1690 ( .A1(n179), .A2(\registers[29][30] ), .B1(n176), .B2(
        \registers[28][30] ), .ZN(n2242) );
  AOI211_X2 U1691 ( .C1(n173), .C2(\registers[1][30] ), .A(n2243), .B(n2244), 
        .ZN(n2233) );
  OAI22_X2 U1692 ( .A1(n34), .A2(n170), .B1(n66), .B2(n167), .ZN(n2244) );
  OAI221_X2 U1693 ( .B1(n130), .B2(n164), .C1(n98), .C2(n161), .A(n2245), .ZN(
        n2243) );
  AOI22_X2 U1694 ( .A1(n30), .A2(\registers[7][30] ), .B1(n27), .B2(
        \registers[6][30] ), .ZN(n2245) );
  AOI221_X2 U1695 ( .B1(n24), .B2(\registers[13][30] ), .C1(n21), .C2(
        \registers[12][30] ), .A(n2246), .ZN(n2232) );
  OAI22_X2 U1696 ( .A1(n418), .A2(n18), .B1(n450), .B2(n15), .ZN(n2246) );
  AOI221_X2 U1697 ( .B1(n12), .B2(\registers[9][30] ), .C1(n9), .C2(
        \registers[8][30] ), .A(n2247), .ZN(n2231) );
  OAI22_X2 U1698 ( .A1(n290), .A2(n6), .B1(n322), .B2(n3), .ZN(n2247) );
  NAND4_X2 U1699 ( .A1(n2248), .A2(n2249), .A3(n2250), .A4(n2251), .ZN(N215)
         );
  NOR4_X2 U1700 ( .A1(n2252), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2251)
         );
  OAI221_X2 U1701 ( .B1(n515), .B2(n221), .C1(n483), .C2(n218), .A(n2256), 
        .ZN(n2255) );
  AOI22_X2 U1702 ( .A1(n215), .A2(\registers[19][29] ), .B1(n212), .B2(
        \registers[18][29] ), .ZN(n2256) );
  OAI221_X2 U1703 ( .B1(n643), .B2(n209), .C1(n611), .C2(n206), .A(n2257), 
        .ZN(n2254) );
  AOI22_X2 U1704 ( .A1(n203), .A2(\registers[23][29] ), .B1(n200), .B2(
        \registers[22][29] ), .ZN(n2257) );
  OAI221_X2 U1705 ( .B1(n835), .B2(n197), .C1(n803), .C2(n194), .A(n2258), 
        .ZN(n2253) );
  AOI22_X2 U1706 ( .A1(n191), .A2(\registers[25][29] ), .B1(n188), .B2(
        \registers[24][29] ), .ZN(n2258) );
  OAI221_X2 U1707 ( .B1(n963), .B2(n185), .C1(n931), .C2(n182), .A(n2259), 
        .ZN(n2252) );
  AOI22_X2 U1708 ( .A1(n179), .A2(\registers[29][29] ), .B1(n176), .B2(
        \registers[28][29] ), .ZN(n2259) );
  AOI211_X2 U1709 ( .C1(n173), .C2(\registers[1][29] ), .A(n2260), .B(n2261), 
        .ZN(n2250) );
  OAI22_X2 U1710 ( .A1(n35), .A2(n170), .B1(n67), .B2(n167), .ZN(n2261) );
  OAI221_X2 U1711 ( .B1(n131), .B2(n164), .C1(n99), .C2(n161), .A(n2262), .ZN(
        n2260) );
  AOI22_X2 U1712 ( .A1(n30), .A2(\registers[7][29] ), .B1(n27), .B2(
        \registers[6][29] ), .ZN(n2262) );
  AOI221_X2 U1713 ( .B1(n24), .B2(\registers[13][29] ), .C1(n21), .C2(
        \registers[12][29] ), .A(n2263), .ZN(n2249) );
  OAI22_X2 U1714 ( .A1(n419), .A2(n18), .B1(n451), .B2(n15), .ZN(n2263) );
  AOI221_X2 U1715 ( .B1(n12), .B2(\registers[9][29] ), .C1(n9), .C2(
        \registers[8][29] ), .A(n2264), .ZN(n2248) );
  OAI22_X2 U1716 ( .A1(n291), .A2(n6), .B1(n323), .B2(n3), .ZN(n2264) );
  NAND4_X2 U1717 ( .A1(n2265), .A2(n2266), .A3(n2267), .A4(n2268), .ZN(N214)
         );
  NOR4_X2 U1718 ( .A1(n2269), .A2(n2270), .A3(n2271), .A4(n2272), .ZN(n2268)
         );
  OAI221_X2 U1719 ( .B1(n516), .B2(n221), .C1(n484), .C2(n218), .A(n2273), 
        .ZN(n2272) );
  AOI22_X2 U1720 ( .A1(n215), .A2(\registers[19][28] ), .B1(n212), .B2(
        \registers[18][28] ), .ZN(n2273) );
  OAI221_X2 U1721 ( .B1(n644), .B2(n209), .C1(n612), .C2(n206), .A(n2274), 
        .ZN(n2271) );
  AOI22_X2 U1722 ( .A1(n203), .A2(\registers[23][28] ), .B1(n200), .B2(
        \registers[22][28] ), .ZN(n2274) );
  OAI221_X2 U1723 ( .B1(n836), .B2(n197), .C1(n804), .C2(n194), .A(n2275), 
        .ZN(n2270) );
  AOI22_X2 U1724 ( .A1(n191), .A2(\registers[25][28] ), .B1(n188), .B2(
        \registers[24][28] ), .ZN(n2275) );
  OAI221_X2 U1725 ( .B1(n964), .B2(n185), .C1(n932), .C2(n182), .A(n2276), 
        .ZN(n2269) );
  AOI22_X2 U1726 ( .A1(n179), .A2(\registers[29][28] ), .B1(n176), .B2(
        \registers[28][28] ), .ZN(n2276) );
  AOI211_X2 U1727 ( .C1(n173), .C2(\registers[1][28] ), .A(n2277), .B(n2278), 
        .ZN(n2267) );
  OAI22_X2 U1728 ( .A1(n36), .A2(n170), .B1(n68), .B2(n167), .ZN(n2278) );
  OAI221_X2 U1729 ( .B1(n132), .B2(n164), .C1(n100), .C2(n161), .A(n2279), 
        .ZN(n2277) );
  AOI22_X2 U1730 ( .A1(n30), .A2(\registers[7][28] ), .B1(n27), .B2(
        \registers[6][28] ), .ZN(n2279) );
  AOI221_X2 U1731 ( .B1(n24), .B2(\registers[13][28] ), .C1(n21), .C2(
        \registers[12][28] ), .A(n2280), .ZN(n2266) );
  OAI22_X2 U1732 ( .A1(n420), .A2(n18), .B1(n452), .B2(n15), .ZN(n2280) );
  AOI221_X2 U1733 ( .B1(n12), .B2(\registers[9][28] ), .C1(n9), .C2(
        \registers[8][28] ), .A(n2281), .ZN(n2265) );
  OAI22_X2 U1734 ( .A1(n292), .A2(n6), .B1(n324), .B2(n3), .ZN(n2281) );
  NAND4_X2 U1735 ( .A1(n2282), .A2(n2283), .A3(n2284), .A4(n2285), .ZN(N213)
         );
  NOR4_X2 U1736 ( .A1(n2286), .A2(n2287), .A3(n2288), .A4(n2289), .ZN(n2285)
         );
  OAI221_X2 U1737 ( .B1(n517), .B2(n221), .C1(n485), .C2(n218), .A(n2290), 
        .ZN(n2289) );
  AOI22_X2 U1738 ( .A1(n215), .A2(\registers[19][27] ), .B1(n212), .B2(
        \registers[18][27] ), .ZN(n2290) );
  OAI221_X2 U1739 ( .B1(n645), .B2(n209), .C1(n613), .C2(n206), .A(n2291), 
        .ZN(n2288) );
  AOI22_X2 U1740 ( .A1(n203), .A2(\registers[23][27] ), .B1(n200), .B2(
        \registers[22][27] ), .ZN(n2291) );
  OAI221_X2 U1741 ( .B1(n837), .B2(n197), .C1(n805), .C2(n194), .A(n2292), 
        .ZN(n2287) );
  AOI22_X2 U1742 ( .A1(n191), .A2(\registers[25][27] ), .B1(n188), .B2(
        \registers[24][27] ), .ZN(n2292) );
  OAI221_X2 U1743 ( .B1(n965), .B2(n185), .C1(n933), .C2(n182), .A(n2293), 
        .ZN(n2286) );
  AOI22_X2 U1744 ( .A1(n179), .A2(\registers[29][27] ), .B1(n176), .B2(
        \registers[28][27] ), .ZN(n2293) );
  AOI211_X2 U1745 ( .C1(n173), .C2(\registers[1][27] ), .A(n2294), .B(n2295), 
        .ZN(n2284) );
  OAI22_X2 U1746 ( .A1(n37), .A2(n170), .B1(n69), .B2(n167), .ZN(n2295) );
  OAI221_X2 U1747 ( .B1(n133), .B2(n164), .C1(n101), .C2(n161), .A(n2296), 
        .ZN(n2294) );
  AOI22_X2 U1748 ( .A1(n30), .A2(\registers[7][27] ), .B1(n27), .B2(
        \registers[6][27] ), .ZN(n2296) );
  AOI221_X2 U1749 ( .B1(n24), .B2(\registers[13][27] ), .C1(n21), .C2(
        \registers[12][27] ), .A(n2297), .ZN(n2283) );
  OAI22_X2 U1750 ( .A1(n421), .A2(n18), .B1(n453), .B2(n15), .ZN(n2297) );
  AOI221_X2 U1751 ( .B1(n12), .B2(\registers[9][27] ), .C1(n9), .C2(
        \registers[8][27] ), .A(n2298), .ZN(n2282) );
  OAI22_X2 U1752 ( .A1(n293), .A2(n6), .B1(n325), .B2(n3), .ZN(n2298) );
  NAND4_X2 U1753 ( .A1(n2299), .A2(n2300), .A3(n2301), .A4(n2302), .ZN(N212)
         );
  NOR4_X2 U1754 ( .A1(n2303), .A2(n2304), .A3(n2305), .A4(n2306), .ZN(n2302)
         );
  OAI221_X2 U1755 ( .B1(n518), .B2(n221), .C1(n486), .C2(n218), .A(n2307), 
        .ZN(n2306) );
  AOI22_X2 U1756 ( .A1(n215), .A2(\registers[19][26] ), .B1(n212), .B2(
        \registers[18][26] ), .ZN(n2307) );
  OAI221_X2 U1757 ( .B1(n646), .B2(n209), .C1(n614), .C2(n206), .A(n2308), 
        .ZN(n2305) );
  AOI22_X2 U1758 ( .A1(n203), .A2(\registers[23][26] ), .B1(n200), .B2(
        \registers[22][26] ), .ZN(n2308) );
  OAI221_X2 U1759 ( .B1(n838), .B2(n197), .C1(n806), .C2(n194), .A(n2309), 
        .ZN(n2304) );
  AOI22_X2 U1760 ( .A1(n191), .A2(\registers[25][26] ), .B1(n188), .B2(
        \registers[24][26] ), .ZN(n2309) );
  OAI221_X2 U1761 ( .B1(n966), .B2(n185), .C1(n934), .C2(n182), .A(n2310), 
        .ZN(n2303) );
  AOI22_X2 U1762 ( .A1(n179), .A2(\registers[29][26] ), .B1(n176), .B2(
        \registers[28][26] ), .ZN(n2310) );
  AOI211_X2 U1763 ( .C1(n173), .C2(\registers[1][26] ), .A(n2311), .B(n2312), 
        .ZN(n2301) );
  OAI22_X2 U1764 ( .A1(n38), .A2(n170), .B1(n70), .B2(n167), .ZN(n2312) );
  OAI221_X2 U1765 ( .B1(n134), .B2(n164), .C1(n102), .C2(n161), .A(n2313), 
        .ZN(n2311) );
  AOI22_X2 U1766 ( .A1(n30), .A2(\registers[7][26] ), .B1(n27), .B2(
        \registers[6][26] ), .ZN(n2313) );
  AOI221_X2 U1767 ( .B1(n24), .B2(\registers[13][26] ), .C1(n21), .C2(
        \registers[12][26] ), .A(n2314), .ZN(n2300) );
  OAI22_X2 U1768 ( .A1(n422), .A2(n18), .B1(n454), .B2(n15), .ZN(n2314) );
  AOI221_X2 U1769 ( .B1(n12), .B2(\registers[9][26] ), .C1(n9), .C2(
        \registers[8][26] ), .A(n2315), .ZN(n2299) );
  OAI22_X2 U1770 ( .A1(n294), .A2(n6), .B1(n326), .B2(n3), .ZN(n2315) );
  NAND4_X2 U1771 ( .A1(n2316), .A2(n2317), .A3(n2318), .A4(n2319), .ZN(N211)
         );
  NOR4_X2 U1772 ( .A1(n2320), .A2(n2321), .A3(n2322), .A4(n2323), .ZN(n2319)
         );
  OAI221_X2 U1773 ( .B1(n519), .B2(n221), .C1(n487), .C2(n218), .A(n2324), 
        .ZN(n2323) );
  AOI22_X2 U1774 ( .A1(n215), .A2(\registers[19][25] ), .B1(n212), .B2(
        \registers[18][25] ), .ZN(n2324) );
  OAI221_X2 U1775 ( .B1(n647), .B2(n209), .C1(n615), .C2(n206), .A(n2325), 
        .ZN(n2322) );
  AOI22_X2 U1776 ( .A1(n203), .A2(\registers[23][25] ), .B1(n200), .B2(
        \registers[22][25] ), .ZN(n2325) );
  OAI221_X2 U1777 ( .B1(n839), .B2(n197), .C1(n807), .C2(n194), .A(n2326), 
        .ZN(n2321) );
  AOI22_X2 U1778 ( .A1(n191), .A2(\registers[25][25] ), .B1(n188), .B2(
        \registers[24][25] ), .ZN(n2326) );
  OAI221_X2 U1779 ( .B1(n967), .B2(n185), .C1(n935), .C2(n182), .A(n2327), 
        .ZN(n2320) );
  AOI22_X2 U1780 ( .A1(n179), .A2(\registers[29][25] ), .B1(n176), .B2(
        \registers[28][25] ), .ZN(n2327) );
  AOI211_X2 U1781 ( .C1(n173), .C2(\registers[1][25] ), .A(n2328), .B(n2329), 
        .ZN(n2318) );
  OAI22_X2 U1782 ( .A1(n39), .A2(n170), .B1(n71), .B2(n167), .ZN(n2329) );
  OAI221_X2 U1783 ( .B1(n135), .B2(n164), .C1(n103), .C2(n161), .A(n2330), 
        .ZN(n2328) );
  AOI22_X2 U1784 ( .A1(n30), .A2(\registers[7][25] ), .B1(n27), .B2(
        \registers[6][25] ), .ZN(n2330) );
  AOI221_X2 U1785 ( .B1(n24), .B2(\registers[13][25] ), .C1(n21), .C2(
        \registers[12][25] ), .A(n2331), .ZN(n2317) );
  OAI22_X2 U1786 ( .A1(n423), .A2(n18), .B1(n455), .B2(n15), .ZN(n2331) );
  AOI221_X2 U1787 ( .B1(n12), .B2(\registers[9][25] ), .C1(n9), .C2(
        \registers[8][25] ), .A(n2332), .ZN(n2316) );
  OAI22_X2 U1788 ( .A1(n295), .A2(n6), .B1(n327), .B2(n3), .ZN(n2332) );
  NAND4_X2 U1789 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(N210)
         );
  NOR4_X2 U1790 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n2336)
         );
  OAI221_X2 U1791 ( .B1(n520), .B2(n221), .C1(n488), .C2(n218), .A(n2341), 
        .ZN(n2340) );
  AOI22_X2 U1792 ( .A1(n215), .A2(\registers[19][24] ), .B1(n212), .B2(
        \registers[18][24] ), .ZN(n2341) );
  OAI221_X2 U1793 ( .B1(n648), .B2(n209), .C1(n616), .C2(n206), .A(n2342), 
        .ZN(n2339) );
  AOI22_X2 U1794 ( .A1(n203), .A2(\registers[23][24] ), .B1(n200), .B2(
        \registers[22][24] ), .ZN(n2342) );
  OAI221_X2 U1795 ( .B1(n840), .B2(n197), .C1(n808), .C2(n194), .A(n2343), 
        .ZN(n2338) );
  AOI22_X2 U1796 ( .A1(n191), .A2(\registers[25][24] ), .B1(n188), .B2(
        \registers[24][24] ), .ZN(n2343) );
  OAI221_X2 U1797 ( .B1(n968), .B2(n185), .C1(n936), .C2(n182), .A(n2344), 
        .ZN(n2337) );
  AOI22_X2 U1798 ( .A1(n179), .A2(\registers[29][24] ), .B1(n176), .B2(
        \registers[28][24] ), .ZN(n2344) );
  AOI211_X2 U1799 ( .C1(n173), .C2(\registers[1][24] ), .A(n2345), .B(n2346), 
        .ZN(n2335) );
  OAI22_X2 U1800 ( .A1(n40), .A2(n170), .B1(n72), .B2(n167), .ZN(n2346) );
  OAI221_X2 U1801 ( .B1(n136), .B2(n164), .C1(n104), .C2(n161), .A(n2347), 
        .ZN(n2345) );
  AOI22_X2 U1802 ( .A1(n30), .A2(\registers[7][24] ), .B1(n27), .B2(
        \registers[6][24] ), .ZN(n2347) );
  AOI221_X2 U1803 ( .B1(n24), .B2(\registers[13][24] ), .C1(n21), .C2(
        \registers[12][24] ), .A(n2348), .ZN(n2334) );
  OAI22_X2 U1804 ( .A1(n424), .A2(n18), .B1(n456), .B2(n15), .ZN(n2348) );
  AOI221_X2 U1805 ( .B1(n12), .B2(\registers[9][24] ), .C1(n9), .C2(
        \registers[8][24] ), .A(n2349), .ZN(n2333) );
  OAI22_X2 U1806 ( .A1(n296), .A2(n6), .B1(n328), .B2(n3), .ZN(n2349) );
  NAND4_X2 U1807 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(N209)
         );
  NOR4_X2 U1808 ( .A1(n2354), .A2(n2355), .A3(n2356), .A4(n2357), .ZN(n2353)
         );
  OAI221_X2 U1809 ( .B1(n521), .B2(n221), .C1(n489), .C2(n218), .A(n2358), 
        .ZN(n2357) );
  AOI22_X2 U1810 ( .A1(n215), .A2(\registers[19][23] ), .B1(n212), .B2(
        \registers[18][23] ), .ZN(n2358) );
  OAI221_X2 U1811 ( .B1(n649), .B2(n209), .C1(n617), .C2(n206), .A(n2359), 
        .ZN(n2356) );
  AOI22_X2 U1812 ( .A1(n203), .A2(\registers[23][23] ), .B1(n200), .B2(
        \registers[22][23] ), .ZN(n2359) );
  OAI221_X2 U1813 ( .B1(n841), .B2(n197), .C1(n809), .C2(n194), .A(n2360), 
        .ZN(n2355) );
  AOI22_X2 U1814 ( .A1(n191), .A2(\registers[25][23] ), .B1(n188), .B2(
        \registers[24][23] ), .ZN(n2360) );
  OAI221_X2 U1815 ( .B1(n969), .B2(n185), .C1(n937), .C2(n182), .A(n2361), 
        .ZN(n2354) );
  AOI22_X2 U1816 ( .A1(n179), .A2(\registers[29][23] ), .B1(n176), .B2(
        \registers[28][23] ), .ZN(n2361) );
  AOI211_X2 U1817 ( .C1(n173), .C2(\registers[1][23] ), .A(n2362), .B(n2363), 
        .ZN(n2352) );
  OAI22_X2 U1818 ( .A1(n41), .A2(n169), .B1(n73), .B2(n166), .ZN(n2363) );
  OAI221_X2 U1819 ( .B1(n137), .B2(n164), .C1(n105), .C2(n161), .A(n2364), 
        .ZN(n2362) );
  AOI22_X2 U1820 ( .A1(n30), .A2(\registers[7][23] ), .B1(n27), .B2(
        \registers[6][23] ), .ZN(n2364) );
  AOI221_X2 U1821 ( .B1(n24), .B2(\registers[13][23] ), .C1(n21), .C2(
        \registers[12][23] ), .A(n2365), .ZN(n2351) );
  OAI22_X2 U1822 ( .A1(n425), .A2(n17), .B1(n457), .B2(n14), .ZN(n2365) );
  AOI221_X2 U1823 ( .B1(n12), .B2(\registers[9][23] ), .C1(n9), .C2(
        \registers[8][23] ), .A(n2366), .ZN(n2350) );
  OAI22_X2 U1824 ( .A1(n297), .A2(n5), .B1(n329), .B2(n2), .ZN(n2366) );
  NAND4_X2 U1825 ( .A1(n2367), .A2(n2368), .A3(n2369), .A4(n2370), .ZN(N208)
         );
  NOR4_X2 U1826 ( .A1(n2371), .A2(n2372), .A3(n2373), .A4(n2374), .ZN(n2370)
         );
  OAI221_X2 U1827 ( .B1(n522), .B2(n221), .C1(n490), .C2(n218), .A(n2375), 
        .ZN(n2374) );
  AOI22_X2 U1828 ( .A1(n215), .A2(\registers[19][22] ), .B1(n212), .B2(
        \registers[18][22] ), .ZN(n2375) );
  OAI221_X2 U1829 ( .B1(n650), .B2(n209), .C1(n618), .C2(n206), .A(n2376), 
        .ZN(n2373) );
  AOI22_X2 U1830 ( .A1(n203), .A2(\registers[23][22] ), .B1(n200), .B2(
        \registers[22][22] ), .ZN(n2376) );
  OAI221_X2 U1831 ( .B1(n842), .B2(n197), .C1(n810), .C2(n194), .A(n2377), 
        .ZN(n2372) );
  AOI22_X2 U1832 ( .A1(n191), .A2(\registers[25][22] ), .B1(n188), .B2(
        \registers[24][22] ), .ZN(n2377) );
  OAI221_X2 U1833 ( .B1(n970), .B2(n185), .C1(n938), .C2(n182), .A(n2378), 
        .ZN(n2371) );
  AOI22_X2 U1834 ( .A1(n179), .A2(\registers[29][22] ), .B1(n176), .B2(
        \registers[28][22] ), .ZN(n2378) );
  AOI211_X2 U1835 ( .C1(n173), .C2(\registers[1][22] ), .A(n2379), .B(n2380), 
        .ZN(n2369) );
  OAI22_X2 U1836 ( .A1(n42), .A2(n169), .B1(n74), .B2(n166), .ZN(n2380) );
  OAI221_X2 U1837 ( .B1(n138), .B2(n164), .C1(n106), .C2(n161), .A(n2381), 
        .ZN(n2379) );
  AOI22_X2 U1838 ( .A1(n30), .A2(\registers[7][22] ), .B1(n27), .B2(
        \registers[6][22] ), .ZN(n2381) );
  AOI221_X2 U1839 ( .B1(n24), .B2(\registers[13][22] ), .C1(n21), .C2(
        \registers[12][22] ), .A(n2382), .ZN(n2368) );
  OAI22_X2 U1840 ( .A1(n426), .A2(n17), .B1(n458), .B2(n14), .ZN(n2382) );
  AOI221_X2 U1841 ( .B1(n12), .B2(\registers[9][22] ), .C1(n9), .C2(
        \registers[8][22] ), .A(n2383), .ZN(n2367) );
  OAI22_X2 U1842 ( .A1(n298), .A2(n5), .B1(n330), .B2(n2), .ZN(n2383) );
  NAND4_X2 U1843 ( .A1(n2384), .A2(n2385), .A3(n2386), .A4(n2387), .ZN(N207)
         );
  NOR4_X2 U1844 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2387)
         );
  OAI221_X2 U1845 ( .B1(n523), .B2(n220), .C1(n491), .C2(n217), .A(n2392), 
        .ZN(n2391) );
  AOI22_X2 U1846 ( .A1(n214), .A2(\registers[19][21] ), .B1(n211), .B2(
        \registers[18][21] ), .ZN(n2392) );
  OAI221_X2 U1847 ( .B1(n651), .B2(n208), .C1(n619), .C2(n205), .A(n2393), 
        .ZN(n2390) );
  AOI22_X2 U1848 ( .A1(n202), .A2(\registers[23][21] ), .B1(n199), .B2(
        \registers[22][21] ), .ZN(n2393) );
  OAI221_X2 U1849 ( .B1(n843), .B2(n196), .C1(n811), .C2(n193), .A(n2394), 
        .ZN(n2389) );
  AOI22_X2 U1850 ( .A1(n190), .A2(\registers[25][21] ), .B1(n187), .B2(
        \registers[24][21] ), .ZN(n2394) );
  OAI221_X2 U1851 ( .B1(n971), .B2(n184), .C1(n939), .C2(n181), .A(n2395), 
        .ZN(n2388) );
  AOI22_X2 U1852 ( .A1(n178), .A2(\registers[29][21] ), .B1(n175), .B2(
        \registers[28][21] ), .ZN(n2395) );
  AOI211_X2 U1853 ( .C1(n172), .C2(\registers[1][21] ), .A(n2396), .B(n2397), 
        .ZN(n2386) );
  OAI22_X2 U1854 ( .A1(n43), .A2(n169), .B1(n75), .B2(n166), .ZN(n2397) );
  OAI221_X2 U1855 ( .B1(n139), .B2(n163), .C1(n107), .C2(n32), .A(n2398), .ZN(
        n2396) );
  AOI22_X2 U1856 ( .A1(n29), .A2(\registers[7][21] ), .B1(n26), .B2(
        \registers[6][21] ), .ZN(n2398) );
  AOI221_X2 U1857 ( .B1(n23), .B2(\registers[13][21] ), .C1(n20), .C2(
        \registers[12][21] ), .A(n2399), .ZN(n2385) );
  OAI22_X2 U1858 ( .A1(n427), .A2(n17), .B1(n459), .B2(n14), .ZN(n2399) );
  AOI221_X2 U1859 ( .B1(n11), .B2(\registers[9][21] ), .C1(n8), .C2(
        \registers[8][21] ), .A(n2400), .ZN(n2384) );
  OAI22_X2 U1860 ( .A1(n299), .A2(n5), .B1(n331), .B2(n2), .ZN(n2400) );
  NAND4_X2 U1861 ( .A1(n2401), .A2(n2402), .A3(n2403), .A4(n2404), .ZN(N206)
         );
  NOR4_X2 U1862 ( .A1(n2405), .A2(n2406), .A3(n2407), .A4(n2408), .ZN(n2404)
         );
  OAI221_X2 U1863 ( .B1(n524), .B2(n220), .C1(n492), .C2(n217), .A(n2409), 
        .ZN(n2408) );
  AOI22_X2 U1864 ( .A1(n214), .A2(\registers[19][20] ), .B1(n211), .B2(
        \registers[18][20] ), .ZN(n2409) );
  OAI221_X2 U1865 ( .B1(n652), .B2(n208), .C1(n620), .C2(n205), .A(n2410), 
        .ZN(n2407) );
  AOI22_X2 U1866 ( .A1(n202), .A2(\registers[23][20] ), .B1(n199), .B2(
        \registers[22][20] ), .ZN(n2410) );
  OAI221_X2 U1867 ( .B1(n844), .B2(n196), .C1(n812), .C2(n193), .A(n2411), 
        .ZN(n2406) );
  AOI22_X2 U1868 ( .A1(n190), .A2(\registers[25][20] ), .B1(n187), .B2(
        \registers[24][20] ), .ZN(n2411) );
  OAI221_X2 U1869 ( .B1(n972), .B2(n184), .C1(n940), .C2(n181), .A(n2412), 
        .ZN(n2405) );
  AOI22_X2 U1870 ( .A1(n178), .A2(\registers[29][20] ), .B1(n175), .B2(
        \registers[28][20] ), .ZN(n2412) );
  AOI211_X2 U1871 ( .C1(n172), .C2(\registers[1][20] ), .A(n2413), .B(n2414), 
        .ZN(n2403) );
  OAI22_X2 U1872 ( .A1(n44), .A2(n169), .B1(n76), .B2(n166), .ZN(n2414) );
  OAI221_X2 U1873 ( .B1(n140), .B2(n163), .C1(n108), .C2(n32), .A(n2415), .ZN(
        n2413) );
  AOI22_X2 U1874 ( .A1(n29), .A2(\registers[7][20] ), .B1(n26), .B2(
        \registers[6][20] ), .ZN(n2415) );
  AOI221_X2 U1875 ( .B1(n23), .B2(\registers[13][20] ), .C1(n20), .C2(
        \registers[12][20] ), .A(n2416), .ZN(n2402) );
  OAI22_X2 U1876 ( .A1(n428), .A2(n17), .B1(n460), .B2(n14), .ZN(n2416) );
  AOI221_X2 U1877 ( .B1(n11), .B2(\registers[9][20] ), .C1(n8), .C2(
        \registers[8][20] ), .A(n2417), .ZN(n2401) );
  OAI22_X2 U1878 ( .A1(n300), .A2(n5), .B1(n332), .B2(n2), .ZN(n2417) );
  NAND4_X2 U1879 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(N205)
         );
  NOR4_X2 U1880 ( .A1(n2422), .A2(n2423), .A3(n2424), .A4(n2425), .ZN(n2421)
         );
  OAI221_X2 U1881 ( .B1(n525), .B2(n220), .C1(n493), .C2(n217), .A(n2426), 
        .ZN(n2425) );
  AOI22_X2 U1882 ( .A1(n214), .A2(\registers[19][19] ), .B1(n211), .B2(
        \registers[18][19] ), .ZN(n2426) );
  OAI221_X2 U1883 ( .B1(n653), .B2(n208), .C1(n621), .C2(n205), .A(n2427), 
        .ZN(n2424) );
  AOI22_X2 U1884 ( .A1(n202), .A2(\registers[23][19] ), .B1(n199), .B2(
        \registers[22][19] ), .ZN(n2427) );
  OAI221_X2 U1885 ( .B1(n845), .B2(n196), .C1(n813), .C2(n193), .A(n2428), 
        .ZN(n2423) );
  AOI22_X2 U1886 ( .A1(n190), .A2(\registers[25][19] ), .B1(n187), .B2(
        \registers[24][19] ), .ZN(n2428) );
  OAI221_X2 U1887 ( .B1(n973), .B2(n184), .C1(n941), .C2(n181), .A(n2429), 
        .ZN(n2422) );
  AOI22_X2 U1888 ( .A1(n178), .A2(\registers[29][19] ), .B1(n175), .B2(
        \registers[28][19] ), .ZN(n2429) );
  AOI211_X2 U1889 ( .C1(n172), .C2(\registers[1][19] ), .A(n2430), .B(n2431), 
        .ZN(n2420) );
  OAI22_X2 U1890 ( .A1(n45), .A2(n169), .B1(n77), .B2(n166), .ZN(n2431) );
  OAI221_X2 U1891 ( .B1(n141), .B2(n163), .C1(n109), .C2(n32), .A(n2432), .ZN(
        n2430) );
  AOI22_X2 U1892 ( .A1(n29), .A2(\registers[7][19] ), .B1(n26), .B2(
        \registers[6][19] ), .ZN(n2432) );
  AOI221_X2 U1893 ( .B1(n23), .B2(\registers[13][19] ), .C1(n20), .C2(
        \registers[12][19] ), .A(n2433), .ZN(n2419) );
  OAI22_X2 U1894 ( .A1(n429), .A2(n17), .B1(n461), .B2(n14), .ZN(n2433) );
  AOI221_X2 U1895 ( .B1(n11), .B2(\registers[9][19] ), .C1(n8), .C2(
        \registers[8][19] ), .A(n2434), .ZN(n2418) );
  OAI22_X2 U1896 ( .A1(n301), .A2(n5), .B1(n333), .B2(n2), .ZN(n2434) );
  NAND4_X2 U1897 ( .A1(n2435), .A2(n2436), .A3(n2437), .A4(n2438), .ZN(N204)
         );
  NOR4_X2 U1898 ( .A1(n2439), .A2(n2440), .A3(n2441), .A4(n2442), .ZN(n2438)
         );
  OAI221_X2 U1899 ( .B1(n526), .B2(n220), .C1(n494), .C2(n217), .A(n2443), 
        .ZN(n2442) );
  AOI22_X2 U1900 ( .A1(n214), .A2(\registers[19][18] ), .B1(n211), .B2(
        \registers[18][18] ), .ZN(n2443) );
  OAI221_X2 U1901 ( .B1(n654), .B2(n208), .C1(n622), .C2(n205), .A(n2444), 
        .ZN(n2441) );
  AOI22_X2 U1902 ( .A1(n202), .A2(\registers[23][18] ), .B1(n199), .B2(
        \registers[22][18] ), .ZN(n2444) );
  OAI221_X2 U1903 ( .B1(n846), .B2(n196), .C1(n814), .C2(n193), .A(n2445), 
        .ZN(n2440) );
  AOI22_X2 U1904 ( .A1(n190), .A2(\registers[25][18] ), .B1(n187), .B2(
        \registers[24][18] ), .ZN(n2445) );
  OAI221_X2 U1905 ( .B1(n974), .B2(n184), .C1(n942), .C2(n181), .A(n2446), 
        .ZN(n2439) );
  AOI22_X2 U1906 ( .A1(n178), .A2(\registers[29][18] ), .B1(n175), .B2(
        \registers[28][18] ), .ZN(n2446) );
  AOI211_X2 U1907 ( .C1(n172), .C2(\registers[1][18] ), .A(n2447), .B(n2448), 
        .ZN(n2437) );
  OAI22_X2 U1908 ( .A1(n46), .A2(n169), .B1(n78), .B2(n166), .ZN(n2448) );
  OAI221_X2 U1909 ( .B1(n142), .B2(n163), .C1(n110), .C2(n32), .A(n2449), .ZN(
        n2447) );
  AOI22_X2 U1910 ( .A1(n29), .A2(\registers[7][18] ), .B1(n26), .B2(
        \registers[6][18] ), .ZN(n2449) );
  AOI221_X2 U1911 ( .B1(n23), .B2(\registers[13][18] ), .C1(n20), .C2(
        \registers[12][18] ), .A(n2450), .ZN(n2436) );
  OAI22_X2 U1912 ( .A1(n430), .A2(n17), .B1(n462), .B2(n14), .ZN(n2450) );
  AOI221_X2 U1913 ( .B1(n11), .B2(\registers[9][18] ), .C1(n8), .C2(
        \registers[8][18] ), .A(n2451), .ZN(n2435) );
  OAI22_X2 U1914 ( .A1(n302), .A2(n5), .B1(n334), .B2(n2), .ZN(n2451) );
  NAND4_X2 U1915 ( .A1(n2452), .A2(n2453), .A3(n2454), .A4(n2455), .ZN(N203)
         );
  NOR4_X2 U1916 ( .A1(n2456), .A2(n2457), .A3(n2458), .A4(n2459), .ZN(n2455)
         );
  OAI221_X2 U1917 ( .B1(n527), .B2(n220), .C1(n495), .C2(n217), .A(n2460), 
        .ZN(n2459) );
  AOI22_X2 U1918 ( .A1(n214), .A2(\registers[19][17] ), .B1(n211), .B2(
        \registers[18][17] ), .ZN(n2460) );
  OAI221_X2 U1919 ( .B1(n655), .B2(n208), .C1(n623), .C2(n205), .A(n2461), 
        .ZN(n2458) );
  AOI22_X2 U1920 ( .A1(n202), .A2(\registers[23][17] ), .B1(n199), .B2(
        \registers[22][17] ), .ZN(n2461) );
  OAI221_X2 U1921 ( .B1(n847), .B2(n196), .C1(n815), .C2(n193), .A(n2462), 
        .ZN(n2457) );
  AOI22_X2 U1922 ( .A1(n190), .A2(\registers[25][17] ), .B1(n187), .B2(
        \registers[24][17] ), .ZN(n2462) );
  OAI221_X2 U1923 ( .B1(n975), .B2(n184), .C1(n943), .C2(n181), .A(n2463), 
        .ZN(n2456) );
  AOI22_X2 U1924 ( .A1(n178), .A2(\registers[29][17] ), .B1(n175), .B2(
        \registers[28][17] ), .ZN(n2463) );
  AOI211_X2 U1925 ( .C1(n172), .C2(\registers[1][17] ), .A(n2464), .B(n2465), 
        .ZN(n2454) );
  OAI22_X2 U1926 ( .A1(n47), .A2(n169), .B1(n79), .B2(n166), .ZN(n2465) );
  OAI221_X2 U1927 ( .B1(n143), .B2(n163), .C1(n111), .C2(n32), .A(n2466), .ZN(
        n2464) );
  AOI22_X2 U1928 ( .A1(n29), .A2(\registers[7][17] ), .B1(n26), .B2(
        \registers[6][17] ), .ZN(n2466) );
  AOI221_X2 U1929 ( .B1(n23), .B2(\registers[13][17] ), .C1(n20), .C2(
        \registers[12][17] ), .A(n2467), .ZN(n2453) );
  OAI22_X2 U1930 ( .A1(n431), .A2(n17), .B1(n463), .B2(n14), .ZN(n2467) );
  AOI221_X2 U1931 ( .B1(n11), .B2(\registers[9][17] ), .C1(n8), .C2(
        \registers[8][17] ), .A(n2468), .ZN(n2452) );
  OAI22_X2 U1932 ( .A1(n303), .A2(n5), .B1(n335), .B2(n2), .ZN(n2468) );
  NAND4_X2 U1933 ( .A1(n2469), .A2(n2470), .A3(n2471), .A4(n2472), .ZN(N202)
         );
  NOR4_X2 U1934 ( .A1(n2473), .A2(n2474), .A3(n2475), .A4(n2476), .ZN(n2472)
         );
  OAI221_X2 U1935 ( .B1(n528), .B2(n220), .C1(n496), .C2(n217), .A(n2477), 
        .ZN(n2476) );
  AOI22_X2 U1936 ( .A1(n214), .A2(\registers[19][16] ), .B1(n211), .B2(
        \registers[18][16] ), .ZN(n2477) );
  OAI221_X2 U1937 ( .B1(n656), .B2(n208), .C1(n624), .C2(n205), .A(n2478), 
        .ZN(n2475) );
  AOI22_X2 U1938 ( .A1(n202), .A2(\registers[23][16] ), .B1(n199), .B2(
        \registers[22][16] ), .ZN(n2478) );
  OAI221_X2 U1939 ( .B1(n848), .B2(n196), .C1(n816), .C2(n193), .A(n2479), 
        .ZN(n2474) );
  AOI22_X2 U1940 ( .A1(n190), .A2(\registers[25][16] ), .B1(n187), .B2(
        \registers[24][16] ), .ZN(n2479) );
  OAI221_X2 U1941 ( .B1(n976), .B2(n184), .C1(n944), .C2(n181), .A(n2480), 
        .ZN(n2473) );
  AOI22_X2 U1942 ( .A1(n178), .A2(\registers[29][16] ), .B1(n175), .B2(
        \registers[28][16] ), .ZN(n2480) );
  AOI211_X2 U1943 ( .C1(n172), .C2(\registers[1][16] ), .A(n2481), .B(n2482), 
        .ZN(n2471) );
  OAI22_X2 U1944 ( .A1(n48), .A2(n169), .B1(n80), .B2(n166), .ZN(n2482) );
  OAI221_X2 U1945 ( .B1(n144), .B2(n163), .C1(n112), .C2(n32), .A(n2483), .ZN(
        n2481) );
  AOI22_X2 U1946 ( .A1(n29), .A2(\registers[7][16] ), .B1(n26), .B2(
        \registers[6][16] ), .ZN(n2483) );
  AOI221_X2 U1947 ( .B1(n23), .B2(\registers[13][16] ), .C1(n20), .C2(
        \registers[12][16] ), .A(n2484), .ZN(n2470) );
  OAI22_X2 U1948 ( .A1(n432), .A2(n17), .B1(n464), .B2(n14), .ZN(n2484) );
  AOI221_X2 U1949 ( .B1(n11), .B2(\registers[9][16] ), .C1(n8), .C2(
        \registers[8][16] ), .A(n2485), .ZN(n2469) );
  OAI22_X2 U1950 ( .A1(n304), .A2(n5), .B1(n336), .B2(n2), .ZN(n2485) );
  NAND4_X2 U1951 ( .A1(n2486), .A2(n2487), .A3(n2488), .A4(n2489), .ZN(N201)
         );
  NOR4_X2 U1952 ( .A1(n2490), .A2(n2491), .A3(n2492), .A4(n2493), .ZN(n2489)
         );
  OAI221_X2 U1953 ( .B1(n529), .B2(n220), .C1(n497), .C2(n217), .A(n2494), 
        .ZN(n2493) );
  AOI22_X2 U1954 ( .A1(n214), .A2(\registers[19][15] ), .B1(n211), .B2(
        \registers[18][15] ), .ZN(n2494) );
  OAI221_X2 U1955 ( .B1(n657), .B2(n208), .C1(n625), .C2(n205), .A(n2495), 
        .ZN(n2492) );
  AOI22_X2 U1956 ( .A1(n202), .A2(\registers[23][15] ), .B1(n199), .B2(
        \registers[22][15] ), .ZN(n2495) );
  OAI221_X2 U1957 ( .B1(n849), .B2(n196), .C1(n817), .C2(n193), .A(n2496), 
        .ZN(n2491) );
  AOI22_X2 U1958 ( .A1(n190), .A2(\registers[25][15] ), .B1(n187), .B2(
        \registers[24][15] ), .ZN(n2496) );
  OAI221_X2 U1959 ( .B1(n977), .B2(n184), .C1(n945), .C2(n181), .A(n2497), 
        .ZN(n2490) );
  AOI22_X2 U1960 ( .A1(n178), .A2(\registers[29][15] ), .B1(n175), .B2(
        \registers[28][15] ), .ZN(n2497) );
  AOI211_X2 U1961 ( .C1(n172), .C2(\registers[1][15] ), .A(n2498), .B(n2499), 
        .ZN(n2488) );
  OAI22_X2 U1962 ( .A1(n49), .A2(n169), .B1(n81), .B2(n166), .ZN(n2499) );
  OAI221_X2 U1963 ( .B1(n145), .B2(n163), .C1(n113), .C2(n32), .A(n2500), .ZN(
        n2498) );
  AOI22_X2 U1964 ( .A1(n29), .A2(\registers[7][15] ), .B1(n26), .B2(
        \registers[6][15] ), .ZN(n2500) );
  AOI221_X2 U1965 ( .B1(n23), .B2(\registers[13][15] ), .C1(n20), .C2(
        \registers[12][15] ), .A(n2501), .ZN(n2487) );
  OAI22_X2 U1966 ( .A1(n433), .A2(n17), .B1(n465), .B2(n14), .ZN(n2501) );
  AOI221_X2 U1967 ( .B1(n11), .B2(\registers[9][15] ), .C1(n8), .C2(
        \registers[8][15] ), .A(n2502), .ZN(n2486) );
  OAI22_X2 U1968 ( .A1(n305), .A2(n5), .B1(n337), .B2(n2), .ZN(n2502) );
  NAND4_X2 U1969 ( .A1(n2503), .A2(n2504), .A3(n2505), .A4(n2506), .ZN(N200)
         );
  NOR4_X2 U1970 ( .A1(n2507), .A2(n2508), .A3(n2509), .A4(n2510), .ZN(n2506)
         );
  OAI221_X2 U1971 ( .B1(n530), .B2(n220), .C1(n498), .C2(n217), .A(n2511), 
        .ZN(n2510) );
  AOI22_X2 U1972 ( .A1(n214), .A2(\registers[19][14] ), .B1(n211), .B2(
        \registers[18][14] ), .ZN(n2511) );
  OAI221_X2 U1973 ( .B1(n658), .B2(n208), .C1(n626), .C2(n205), .A(n2512), 
        .ZN(n2509) );
  AOI22_X2 U1974 ( .A1(n202), .A2(\registers[23][14] ), .B1(n199), .B2(
        \registers[22][14] ), .ZN(n2512) );
  OAI221_X2 U1975 ( .B1(n850), .B2(n196), .C1(n818), .C2(n193), .A(n2513), 
        .ZN(n2508) );
  AOI22_X2 U1976 ( .A1(n190), .A2(\registers[25][14] ), .B1(n187), .B2(
        \registers[24][14] ), .ZN(n2513) );
  OAI221_X2 U1977 ( .B1(n978), .B2(n184), .C1(n946), .C2(n181), .A(n2514), 
        .ZN(n2507) );
  AOI22_X2 U1978 ( .A1(n178), .A2(\registers[29][14] ), .B1(n175), .B2(
        \registers[28][14] ), .ZN(n2514) );
  AOI211_X2 U1979 ( .C1(n172), .C2(\registers[1][14] ), .A(n2515), .B(n2516), 
        .ZN(n2505) );
  OAI22_X2 U1980 ( .A1(n50), .A2(n169), .B1(n82), .B2(n166), .ZN(n2516) );
  OAI221_X2 U1981 ( .B1(n146), .B2(n163), .C1(n114), .C2(n32), .A(n2517), .ZN(
        n2515) );
  AOI22_X2 U1982 ( .A1(n29), .A2(\registers[7][14] ), .B1(n26), .B2(
        \registers[6][14] ), .ZN(n2517) );
  AOI221_X2 U1983 ( .B1(n23), .B2(\registers[13][14] ), .C1(n20), .C2(
        \registers[12][14] ), .A(n2518), .ZN(n2504) );
  OAI22_X2 U1984 ( .A1(n434), .A2(n17), .B1(n466), .B2(n14), .ZN(n2518) );
  AOI221_X2 U1985 ( .B1(n11), .B2(\registers[9][14] ), .C1(n8), .C2(
        \registers[8][14] ), .A(n2519), .ZN(n2503) );
  OAI22_X2 U1986 ( .A1(n306), .A2(n5), .B1(n338), .B2(n2), .ZN(n2519) );
  NAND4_X2 U1987 ( .A1(n2520), .A2(n2521), .A3(n2522), .A4(n2523), .ZN(N199)
         );
  NOR4_X2 U1988 ( .A1(n2524), .A2(n2525), .A3(n2526), .A4(n2527), .ZN(n2523)
         );
  OAI221_X2 U1989 ( .B1(n531), .B2(n220), .C1(n499), .C2(n217), .A(n2528), 
        .ZN(n2527) );
  AOI22_X2 U1990 ( .A1(n214), .A2(\registers[19][13] ), .B1(n211), .B2(
        \registers[18][13] ), .ZN(n2528) );
  OAI221_X2 U1991 ( .B1(n659), .B2(n208), .C1(n627), .C2(n205), .A(n2529), 
        .ZN(n2526) );
  AOI22_X2 U1992 ( .A1(n202), .A2(\registers[23][13] ), .B1(n199), .B2(
        \registers[22][13] ), .ZN(n2529) );
  OAI221_X2 U1993 ( .B1(n851), .B2(n196), .C1(n819), .C2(n193), .A(n2530), 
        .ZN(n2525) );
  AOI22_X2 U1994 ( .A1(n190), .A2(\registers[25][13] ), .B1(n187), .B2(
        \registers[24][13] ), .ZN(n2530) );
  OAI221_X2 U1995 ( .B1(n979), .B2(n184), .C1(n947), .C2(n181), .A(n2531), 
        .ZN(n2524) );
  AOI22_X2 U1996 ( .A1(n178), .A2(\registers[29][13] ), .B1(n175), .B2(
        \registers[28][13] ), .ZN(n2531) );
  AOI211_X2 U1997 ( .C1(n172), .C2(\registers[1][13] ), .A(n2532), .B(n2533), 
        .ZN(n2522) );
  OAI22_X2 U1998 ( .A1(n51), .A2(n169), .B1(n83), .B2(n166), .ZN(n2533) );
  OAI221_X2 U1999 ( .B1(n147), .B2(n163), .C1(n115), .C2(n32), .A(n2534), .ZN(
        n2532) );
  AOI22_X2 U2000 ( .A1(n29), .A2(\registers[7][13] ), .B1(n26), .B2(
        \registers[6][13] ), .ZN(n2534) );
  AOI221_X2 U2001 ( .B1(n23), .B2(\registers[13][13] ), .C1(n20), .C2(
        \registers[12][13] ), .A(n2535), .ZN(n2521) );
  OAI22_X2 U2002 ( .A1(n435), .A2(n17), .B1(n467), .B2(n14), .ZN(n2535) );
  AOI221_X2 U2003 ( .B1(n11), .B2(\registers[9][13] ), .C1(n8), .C2(
        \registers[8][13] ), .A(n2536), .ZN(n2520) );
  OAI22_X2 U2004 ( .A1(n307), .A2(n5), .B1(n339), .B2(n2), .ZN(n2536) );
  NAND4_X2 U2005 ( .A1(n2537), .A2(n2538), .A3(n2539), .A4(n2540), .ZN(N198)
         );
  NOR4_X2 U2006 ( .A1(n2541), .A2(n2542), .A3(n2543), .A4(n2544), .ZN(n2540)
         );
  OAI221_X2 U2007 ( .B1(n532), .B2(n220), .C1(n500), .C2(n217), .A(n2545), 
        .ZN(n2544) );
  AOI22_X2 U2008 ( .A1(n214), .A2(\registers[19][12] ), .B1(n211), .B2(
        \registers[18][12] ), .ZN(n2545) );
  OAI221_X2 U2009 ( .B1(n660), .B2(n208), .C1(n628), .C2(n205), .A(n2546), 
        .ZN(n2543) );
  AOI22_X2 U2010 ( .A1(n202), .A2(\registers[23][12] ), .B1(n199), .B2(
        \registers[22][12] ), .ZN(n2546) );
  OAI221_X2 U2011 ( .B1(n852), .B2(n196), .C1(n820), .C2(n193), .A(n2547), 
        .ZN(n2542) );
  AOI22_X2 U2012 ( .A1(n190), .A2(\registers[25][12] ), .B1(n187), .B2(
        \registers[24][12] ), .ZN(n2547) );
  OAI221_X2 U2013 ( .B1(n980), .B2(n184), .C1(n948), .C2(n181), .A(n2548), 
        .ZN(n2541) );
  AOI22_X2 U2014 ( .A1(n178), .A2(\registers[29][12] ), .B1(n175), .B2(
        \registers[28][12] ), .ZN(n2548) );
  AOI211_X2 U2015 ( .C1(n172), .C2(\registers[1][12] ), .A(n2549), .B(n2550), 
        .ZN(n2539) );
  OAI22_X2 U2016 ( .A1(n52), .A2(n169), .B1(n84), .B2(n166), .ZN(n2550) );
  OAI221_X2 U2017 ( .B1(n148), .B2(n163), .C1(n116), .C2(n32), .A(n2551), .ZN(
        n2549) );
  AOI22_X2 U2018 ( .A1(n29), .A2(\registers[7][12] ), .B1(n26), .B2(
        \registers[6][12] ), .ZN(n2551) );
  AOI221_X2 U2019 ( .B1(n23), .B2(\registers[13][12] ), .C1(n20), .C2(
        \registers[12][12] ), .A(n2552), .ZN(n2538) );
  OAI22_X2 U2020 ( .A1(n436), .A2(n17), .B1(n468), .B2(n14), .ZN(n2552) );
  AOI221_X2 U2021 ( .B1(n11), .B2(\registers[9][12] ), .C1(n8), .C2(
        \registers[8][12] ), .A(n2553), .ZN(n2537) );
  OAI22_X2 U2022 ( .A1(n308), .A2(n5), .B1(n340), .B2(n2), .ZN(n2553) );
  NAND4_X2 U2023 ( .A1(n2554), .A2(n2555), .A3(n2556), .A4(n2557), .ZN(N197)
         );
  NOR4_X2 U2024 ( .A1(n2558), .A2(n2559), .A3(n2560), .A4(n2561), .ZN(n2557)
         );
  OAI221_X2 U2025 ( .B1(n533), .B2(n220), .C1(n501), .C2(n217), .A(n2562), 
        .ZN(n2561) );
  AOI22_X2 U2026 ( .A1(n214), .A2(\registers[19][11] ), .B1(n211), .B2(
        \registers[18][11] ), .ZN(n2562) );
  OAI221_X2 U2027 ( .B1(n661), .B2(n208), .C1(n629), .C2(n205), .A(n2563), 
        .ZN(n2560) );
  AOI22_X2 U2028 ( .A1(n202), .A2(\registers[23][11] ), .B1(n199), .B2(
        \registers[22][11] ), .ZN(n2563) );
  OAI221_X2 U2029 ( .B1(n853), .B2(n196), .C1(n821), .C2(n193), .A(n2564), 
        .ZN(n2559) );
  AOI22_X2 U2030 ( .A1(n190), .A2(\registers[25][11] ), .B1(n187), .B2(
        \registers[24][11] ), .ZN(n2564) );
  OAI221_X2 U2031 ( .B1(n981), .B2(n184), .C1(n949), .C2(n181), .A(n2565), 
        .ZN(n2558) );
  AOI22_X2 U2032 ( .A1(n178), .A2(\registers[29][11] ), .B1(n175), .B2(
        \registers[28][11] ), .ZN(n2565) );
  AOI211_X2 U2033 ( .C1(n172), .C2(\registers[1][11] ), .A(n2566), .B(n2567), 
        .ZN(n2556) );
  OAI22_X2 U2034 ( .A1(n53), .A2(n168), .B1(n85), .B2(n165), .ZN(n2567) );
  OAI221_X2 U2035 ( .B1(n149), .B2(n163), .C1(n117), .C2(n32), .A(n2568), .ZN(
        n2566) );
  AOI22_X2 U2036 ( .A1(n29), .A2(\registers[7][11] ), .B1(n26), .B2(
        \registers[6][11] ), .ZN(n2568) );
  AOI221_X2 U2037 ( .B1(n23), .B2(\registers[13][11] ), .C1(n20), .C2(
        \registers[12][11] ), .A(n2569), .ZN(n2555) );
  OAI22_X2 U2038 ( .A1(n437), .A2(n16), .B1(n469), .B2(n13), .ZN(n2569) );
  AOI221_X2 U2039 ( .B1(n11), .B2(\registers[9][11] ), .C1(n8), .C2(
        \registers[8][11] ), .A(n2570), .ZN(n2554) );
  OAI22_X2 U2040 ( .A1(n309), .A2(n4), .B1(n341), .B2(n1), .ZN(n2570) );
  NAND4_X2 U2041 ( .A1(n2571), .A2(n2572), .A3(n2573), .A4(n2574), .ZN(N196)
         );
  NOR4_X2 U2042 ( .A1(n2575), .A2(n2576), .A3(n2577), .A4(n2578), .ZN(n2574)
         );
  OAI221_X2 U2043 ( .B1(n534), .B2(n219), .C1(n502), .C2(n216), .A(n2579), 
        .ZN(n2578) );
  AOI22_X2 U2044 ( .A1(n213), .A2(\registers[19][10] ), .B1(n210), .B2(
        \registers[18][10] ), .ZN(n2579) );
  OAI221_X2 U2045 ( .B1(n662), .B2(n207), .C1(n630), .C2(n204), .A(n2580), 
        .ZN(n2577) );
  AOI22_X2 U2046 ( .A1(n201), .A2(\registers[23][10] ), .B1(n198), .B2(
        \registers[22][10] ), .ZN(n2580) );
  OAI221_X2 U2047 ( .B1(n854), .B2(n195), .C1(n822), .C2(n192), .A(n2581), 
        .ZN(n2576) );
  AOI22_X2 U2048 ( .A1(n189), .A2(\registers[25][10] ), .B1(n186), .B2(
        \registers[24][10] ), .ZN(n2581) );
  OAI221_X2 U2049 ( .B1(n982), .B2(n183), .C1(n950), .C2(n180), .A(n2582), 
        .ZN(n2575) );
  AOI22_X2 U2050 ( .A1(n177), .A2(\registers[29][10] ), .B1(n174), .B2(
        \registers[28][10] ), .ZN(n2582) );
  AOI211_X2 U2051 ( .C1(n171), .C2(\registers[1][10] ), .A(n2583), .B(n2584), 
        .ZN(n2573) );
  OAI22_X2 U2052 ( .A1(n54), .A2(n168), .B1(n86), .B2(n165), .ZN(n2584) );
  OAI221_X2 U2053 ( .B1(n150), .B2(n162), .C1(n118), .C2(n31), .A(n2585), .ZN(
        n2583) );
  AOI22_X2 U2054 ( .A1(n28), .A2(\registers[7][10] ), .B1(n25), .B2(
        \registers[6][10] ), .ZN(n2585) );
  AOI221_X2 U2055 ( .B1(n22), .B2(\registers[13][10] ), .C1(n19), .C2(
        \registers[12][10] ), .A(n2586), .ZN(n2572) );
  OAI22_X2 U2056 ( .A1(n438), .A2(n16), .B1(n470), .B2(n13), .ZN(n2586) );
  AOI221_X2 U2057 ( .B1(n10), .B2(\registers[9][10] ), .C1(n7), .C2(
        \registers[8][10] ), .A(n2587), .ZN(n2571) );
  OAI22_X2 U2058 ( .A1(n310), .A2(n4), .B1(n342), .B2(n1), .ZN(n2587) );
  NAND4_X2 U2059 ( .A1(n2588), .A2(n2589), .A3(n2590), .A4(n2591), .ZN(N195)
         );
  NOR4_X2 U2060 ( .A1(n2592), .A2(n2593), .A3(n2594), .A4(n2595), .ZN(n2591)
         );
  OAI221_X2 U2061 ( .B1(n535), .B2(n219), .C1(n503), .C2(n216), .A(n2596), 
        .ZN(n2595) );
  AOI22_X2 U2062 ( .A1(n213), .A2(\registers[19][9] ), .B1(n210), .B2(
        \registers[18][9] ), .ZN(n2596) );
  OAI221_X2 U2063 ( .B1(n663), .B2(n207), .C1(n631), .C2(n204), .A(n2597), 
        .ZN(n2594) );
  AOI22_X2 U2064 ( .A1(n201), .A2(\registers[23][9] ), .B1(n198), .B2(
        \registers[22][9] ), .ZN(n2597) );
  OAI221_X2 U2065 ( .B1(n855), .B2(n195), .C1(n823), .C2(n192), .A(n2598), 
        .ZN(n2593) );
  AOI22_X2 U2066 ( .A1(n189), .A2(\registers[25][9] ), .B1(n186), .B2(
        \registers[24][9] ), .ZN(n2598) );
  OAI221_X2 U2067 ( .B1(n983), .B2(n183), .C1(n951), .C2(n180), .A(n2599), 
        .ZN(n2592) );
  AOI22_X2 U2068 ( .A1(n177), .A2(\registers[29][9] ), .B1(n174), .B2(
        \registers[28][9] ), .ZN(n2599) );
  AOI211_X2 U2069 ( .C1(n171), .C2(\registers[1][9] ), .A(n2600), .B(n2601), 
        .ZN(n2590) );
  OAI22_X2 U2070 ( .A1(n55), .A2(n168), .B1(n87), .B2(n165), .ZN(n2601) );
  OAI221_X2 U2071 ( .B1(n151), .B2(n162), .C1(n119), .C2(n31), .A(n2602), .ZN(
        n2600) );
  AOI22_X2 U2072 ( .A1(n28), .A2(\registers[7][9] ), .B1(n25), .B2(
        \registers[6][9] ), .ZN(n2602) );
  AOI221_X2 U2073 ( .B1(n22), .B2(\registers[13][9] ), .C1(n19), .C2(
        \registers[12][9] ), .A(n2603), .ZN(n2589) );
  OAI22_X2 U2074 ( .A1(n439), .A2(n16), .B1(n471), .B2(n13), .ZN(n2603) );
  AOI221_X2 U2075 ( .B1(n10), .B2(\registers[9][9] ), .C1(n7), .C2(
        \registers[8][9] ), .A(n2604), .ZN(n2588) );
  OAI22_X2 U2076 ( .A1(n311), .A2(n4), .B1(n343), .B2(n1), .ZN(n2604) );
  NAND4_X2 U2077 ( .A1(n2605), .A2(n2606), .A3(n2607), .A4(n2608), .ZN(N194)
         );
  NOR4_X2 U2078 ( .A1(n2609), .A2(n2610), .A3(n2611), .A4(n2612), .ZN(n2608)
         );
  OAI221_X2 U2079 ( .B1(n536), .B2(n219), .C1(n504), .C2(n216), .A(n2613), 
        .ZN(n2612) );
  AOI22_X2 U2080 ( .A1(n213), .A2(\registers[19][8] ), .B1(n210), .B2(
        \registers[18][8] ), .ZN(n2613) );
  OAI221_X2 U2081 ( .B1(n664), .B2(n207), .C1(n632), .C2(n204), .A(n2614), 
        .ZN(n2611) );
  AOI22_X2 U2082 ( .A1(n201), .A2(\registers[23][8] ), .B1(n198), .B2(
        \registers[22][8] ), .ZN(n2614) );
  OAI221_X2 U2083 ( .B1(n856), .B2(n195), .C1(n824), .C2(n192), .A(n2615), 
        .ZN(n2610) );
  AOI22_X2 U2084 ( .A1(n189), .A2(\registers[25][8] ), .B1(n186), .B2(
        \registers[24][8] ), .ZN(n2615) );
  OAI221_X2 U2085 ( .B1(n984), .B2(n183), .C1(n952), .C2(n180), .A(n2616), 
        .ZN(n2609) );
  AOI22_X2 U2086 ( .A1(n177), .A2(\registers[29][8] ), .B1(n174), .B2(
        \registers[28][8] ), .ZN(n2616) );
  AOI211_X2 U2087 ( .C1(n171), .C2(\registers[1][8] ), .A(n2617), .B(n2618), 
        .ZN(n2607) );
  OAI22_X2 U2088 ( .A1(n56), .A2(n168), .B1(n88), .B2(n165), .ZN(n2618) );
  OAI221_X2 U2089 ( .B1(n152), .B2(n162), .C1(n120), .C2(n31), .A(n2619), .ZN(
        n2617) );
  AOI22_X2 U2090 ( .A1(n28), .A2(\registers[7][8] ), .B1(n25), .B2(
        \registers[6][8] ), .ZN(n2619) );
  AOI221_X2 U2091 ( .B1(n22), .B2(\registers[13][8] ), .C1(n19), .C2(
        \registers[12][8] ), .A(n2620), .ZN(n2606) );
  OAI22_X2 U2092 ( .A1(n440), .A2(n16), .B1(n472), .B2(n13), .ZN(n2620) );
  AOI221_X2 U2093 ( .B1(n10), .B2(\registers[9][8] ), .C1(n7), .C2(
        \registers[8][8] ), .A(n2621), .ZN(n2605) );
  OAI22_X2 U2094 ( .A1(n312), .A2(n4), .B1(n344), .B2(n1), .ZN(n2621) );
  NAND4_X2 U2095 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(N193)
         );
  NOR4_X2 U2096 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(n2625)
         );
  OAI221_X2 U2097 ( .B1(n537), .B2(n219), .C1(n505), .C2(n216), .A(n2630), 
        .ZN(n2629) );
  AOI22_X2 U2098 ( .A1(n213), .A2(\registers[19][7] ), .B1(n210), .B2(
        \registers[18][7] ), .ZN(n2630) );
  OAI221_X2 U2099 ( .B1(n665), .B2(n207), .C1(n633), .C2(n204), .A(n2631), 
        .ZN(n2628) );
  AOI22_X2 U2100 ( .A1(n201), .A2(\registers[23][7] ), .B1(n198), .B2(
        \registers[22][7] ), .ZN(n2631) );
  OAI221_X2 U2101 ( .B1(n857), .B2(n195), .C1(n825), .C2(n192), .A(n2632), 
        .ZN(n2627) );
  AOI22_X2 U2102 ( .A1(n189), .A2(\registers[25][7] ), .B1(n186), .B2(
        \registers[24][7] ), .ZN(n2632) );
  OAI221_X2 U2103 ( .B1(n985), .B2(n183), .C1(n953), .C2(n180), .A(n2633), 
        .ZN(n2626) );
  AOI22_X2 U2104 ( .A1(n177), .A2(\registers[29][7] ), .B1(n174), .B2(
        \registers[28][7] ), .ZN(n2633) );
  AOI211_X2 U2105 ( .C1(n171), .C2(\registers[1][7] ), .A(n2634), .B(n2635), 
        .ZN(n2624) );
  OAI22_X2 U2106 ( .A1(n57), .A2(n168), .B1(n89), .B2(n165), .ZN(n2635) );
  OAI221_X2 U2107 ( .B1(n153), .B2(n162), .C1(n121), .C2(n31), .A(n2636), .ZN(
        n2634) );
  AOI22_X2 U2108 ( .A1(n28), .A2(\registers[7][7] ), .B1(n25), .B2(
        \registers[6][7] ), .ZN(n2636) );
  AOI221_X2 U2109 ( .B1(n22), .B2(\registers[13][7] ), .C1(n19), .C2(
        \registers[12][7] ), .A(n2637), .ZN(n2623) );
  OAI22_X2 U2110 ( .A1(n441), .A2(n16), .B1(n473), .B2(n13), .ZN(n2637) );
  AOI221_X2 U2111 ( .B1(n10), .B2(\registers[9][7] ), .C1(n7), .C2(
        \registers[8][7] ), .A(n2638), .ZN(n2622) );
  OAI22_X2 U2112 ( .A1(n313), .A2(n4), .B1(n345), .B2(n1), .ZN(n2638) );
  NAND4_X2 U2113 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2642), .ZN(N192)
         );
  NOR4_X2 U2114 ( .A1(n2643), .A2(n2644), .A3(n2645), .A4(n2646), .ZN(n2642)
         );
  OAI221_X2 U2115 ( .B1(n538), .B2(n219), .C1(n506), .C2(n216), .A(n2647), 
        .ZN(n2646) );
  AOI22_X2 U2116 ( .A1(n213), .A2(\registers[19][6] ), .B1(n210), .B2(
        \registers[18][6] ), .ZN(n2647) );
  OAI221_X2 U2117 ( .B1(n666), .B2(n207), .C1(n634), .C2(n204), .A(n2648), 
        .ZN(n2645) );
  AOI22_X2 U2118 ( .A1(n201), .A2(\registers[23][6] ), .B1(n198), .B2(
        \registers[22][6] ), .ZN(n2648) );
  OAI221_X2 U2119 ( .B1(n858), .B2(n195), .C1(n826), .C2(n192), .A(n2649), 
        .ZN(n2644) );
  AOI22_X2 U2120 ( .A1(n189), .A2(\registers[25][6] ), .B1(n186), .B2(
        \registers[24][6] ), .ZN(n2649) );
  OAI221_X2 U2121 ( .B1(n986), .B2(n183), .C1(n954), .C2(n180), .A(n2650), 
        .ZN(n2643) );
  AOI22_X2 U2122 ( .A1(n177), .A2(\registers[29][6] ), .B1(n174), .B2(
        \registers[28][6] ), .ZN(n2650) );
  AOI211_X2 U2123 ( .C1(n171), .C2(\registers[1][6] ), .A(n2651), .B(n2652), 
        .ZN(n2641) );
  OAI22_X2 U2124 ( .A1(n58), .A2(n168), .B1(n90), .B2(n165), .ZN(n2652) );
  OAI221_X2 U2125 ( .B1(n154), .B2(n162), .C1(n122), .C2(n31), .A(n2653), .ZN(
        n2651) );
  AOI22_X2 U2126 ( .A1(n28), .A2(\registers[7][6] ), .B1(n25), .B2(
        \registers[6][6] ), .ZN(n2653) );
  AOI221_X2 U2127 ( .B1(n22), .B2(\registers[13][6] ), .C1(n19), .C2(
        \registers[12][6] ), .A(n2654), .ZN(n2640) );
  OAI22_X2 U2128 ( .A1(n442), .A2(n16), .B1(n474), .B2(n13), .ZN(n2654) );
  AOI221_X2 U2129 ( .B1(n10), .B2(\registers[9][6] ), .C1(n7), .C2(
        \registers[8][6] ), .A(n2655), .ZN(n2639) );
  OAI22_X2 U2130 ( .A1(n314), .A2(n4), .B1(n346), .B2(n1), .ZN(n2655) );
  NAND4_X2 U2131 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(N191)
         );
  NOR4_X2 U2132 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(n2659)
         );
  OAI221_X2 U2133 ( .B1(n539), .B2(n219), .C1(n507), .C2(n216), .A(n2664), 
        .ZN(n2663) );
  AOI22_X2 U2134 ( .A1(n213), .A2(\registers[19][5] ), .B1(n210), .B2(
        \registers[18][5] ), .ZN(n2664) );
  OAI221_X2 U2135 ( .B1(n667), .B2(n207), .C1(n635), .C2(n204), .A(n2665), 
        .ZN(n2662) );
  AOI22_X2 U2136 ( .A1(n201), .A2(\registers[23][5] ), .B1(n198), .B2(
        \registers[22][5] ), .ZN(n2665) );
  OAI221_X2 U2137 ( .B1(n859), .B2(n195), .C1(n827), .C2(n192), .A(n2666), 
        .ZN(n2661) );
  AOI22_X2 U2138 ( .A1(n189), .A2(\registers[25][5] ), .B1(n186), .B2(
        \registers[24][5] ), .ZN(n2666) );
  OAI221_X2 U2139 ( .B1(n987), .B2(n183), .C1(n955), .C2(n180), .A(n2667), 
        .ZN(n2660) );
  AOI22_X2 U2140 ( .A1(n177), .A2(\registers[29][5] ), .B1(n174), .B2(
        \registers[28][5] ), .ZN(n2667) );
  AOI211_X2 U2141 ( .C1(n171), .C2(\registers[1][5] ), .A(n2668), .B(n2669), 
        .ZN(n2658) );
  OAI22_X2 U2142 ( .A1(n59), .A2(n168), .B1(n91), .B2(n165), .ZN(n2669) );
  OAI221_X2 U2143 ( .B1(n155), .B2(n162), .C1(n123), .C2(n31), .A(n2670), .ZN(
        n2668) );
  AOI22_X2 U2144 ( .A1(n28), .A2(\registers[7][5] ), .B1(n25), .B2(
        \registers[6][5] ), .ZN(n2670) );
  AOI221_X2 U2145 ( .B1(n22), .B2(\registers[13][5] ), .C1(n19), .C2(
        \registers[12][5] ), .A(n2671), .ZN(n2657) );
  OAI22_X2 U2146 ( .A1(n443), .A2(n16), .B1(n475), .B2(n13), .ZN(n2671) );
  AOI221_X2 U2147 ( .B1(n10), .B2(\registers[9][5] ), .C1(n7), .C2(
        \registers[8][5] ), .A(n2672), .ZN(n2656) );
  OAI22_X2 U2148 ( .A1(n315), .A2(n4), .B1(n347), .B2(n1), .ZN(n2672) );
  NAND4_X2 U2149 ( .A1(n2673), .A2(n2674), .A3(n2675), .A4(n2676), .ZN(N190)
         );
  NOR4_X2 U2150 ( .A1(n2677), .A2(n2678), .A3(n2679), .A4(n2680), .ZN(n2676)
         );
  OAI221_X2 U2151 ( .B1(n540), .B2(n219), .C1(n508), .C2(n216), .A(n2681), 
        .ZN(n2680) );
  AOI22_X2 U2152 ( .A1(n213), .A2(\registers[19][4] ), .B1(n210), .B2(
        \registers[18][4] ), .ZN(n2681) );
  OAI221_X2 U2153 ( .B1(n668), .B2(n207), .C1(n636), .C2(n204), .A(n2682), 
        .ZN(n2679) );
  AOI22_X2 U2154 ( .A1(n201), .A2(\registers[23][4] ), .B1(n198), .B2(
        \registers[22][4] ), .ZN(n2682) );
  OAI221_X2 U2155 ( .B1(n860), .B2(n195), .C1(n828), .C2(n192), .A(n2683), 
        .ZN(n2678) );
  AOI22_X2 U2156 ( .A1(n189), .A2(\registers[25][4] ), .B1(n186), .B2(
        \registers[24][4] ), .ZN(n2683) );
  OAI221_X2 U2157 ( .B1(n988), .B2(n183), .C1(n956), .C2(n180), .A(n2684), 
        .ZN(n2677) );
  AOI22_X2 U2158 ( .A1(n177), .A2(\registers[29][4] ), .B1(n174), .B2(
        \registers[28][4] ), .ZN(n2684) );
  AOI211_X2 U2159 ( .C1(n171), .C2(\registers[1][4] ), .A(n2685), .B(n2686), 
        .ZN(n2675) );
  OAI22_X2 U2160 ( .A1(n60), .A2(n168), .B1(n92), .B2(n165), .ZN(n2686) );
  OAI221_X2 U2161 ( .B1(n156), .B2(n162), .C1(n124), .C2(n31), .A(n2687), .ZN(
        n2685) );
  AOI22_X2 U2162 ( .A1(n28), .A2(\registers[7][4] ), .B1(n25), .B2(
        \registers[6][4] ), .ZN(n2687) );
  AOI221_X2 U2163 ( .B1(n22), .B2(\registers[13][4] ), .C1(n19), .C2(
        \registers[12][4] ), .A(n2688), .ZN(n2674) );
  OAI22_X2 U2164 ( .A1(n444), .A2(n16), .B1(n476), .B2(n13), .ZN(n2688) );
  AOI221_X2 U2165 ( .B1(n10), .B2(\registers[9][4] ), .C1(n7), .C2(
        \registers[8][4] ), .A(n2689), .ZN(n2673) );
  OAI22_X2 U2166 ( .A1(n316), .A2(n4), .B1(n348), .B2(n1), .ZN(n2689) );
  NAND4_X2 U2167 ( .A1(n2690), .A2(n2691), .A3(n2692), .A4(n2693), .ZN(N189)
         );
  NOR4_X2 U2168 ( .A1(n2694), .A2(n2695), .A3(n2696), .A4(n2697), .ZN(n2693)
         );
  OAI221_X2 U2169 ( .B1(n541), .B2(n219), .C1(n509), .C2(n216), .A(n2698), 
        .ZN(n2697) );
  AOI22_X2 U2170 ( .A1(n213), .A2(\registers[19][3] ), .B1(n210), .B2(
        \registers[18][3] ), .ZN(n2698) );
  OAI221_X2 U2171 ( .B1(n669), .B2(n207), .C1(n637), .C2(n204), .A(n2699), 
        .ZN(n2696) );
  AOI22_X2 U2172 ( .A1(n201), .A2(\registers[23][3] ), .B1(n198), .B2(
        \registers[22][3] ), .ZN(n2699) );
  OAI221_X2 U2173 ( .B1(n861), .B2(n195), .C1(n829), .C2(n192), .A(n2700), 
        .ZN(n2695) );
  AOI22_X2 U2174 ( .A1(n189), .A2(\registers[25][3] ), .B1(n186), .B2(
        \registers[24][3] ), .ZN(n2700) );
  OAI221_X2 U2175 ( .B1(n989), .B2(n183), .C1(n957), .C2(n180), .A(n2701), 
        .ZN(n2694) );
  AOI22_X2 U2176 ( .A1(n177), .A2(\registers[29][3] ), .B1(n174), .B2(
        \registers[28][3] ), .ZN(n2701) );
  AOI211_X2 U2177 ( .C1(n171), .C2(\registers[1][3] ), .A(n2702), .B(n2703), 
        .ZN(n2692) );
  OAI22_X2 U2178 ( .A1(n61), .A2(n168), .B1(n93), .B2(n165), .ZN(n2703) );
  OAI221_X2 U2179 ( .B1(n157), .B2(n162), .C1(n125), .C2(n31), .A(n2704), .ZN(
        n2702) );
  AOI22_X2 U2180 ( .A1(n28), .A2(\registers[7][3] ), .B1(n25), .B2(
        \registers[6][3] ), .ZN(n2704) );
  AOI221_X2 U2181 ( .B1(n22), .B2(\registers[13][3] ), .C1(n19), .C2(
        \registers[12][3] ), .A(n2705), .ZN(n2691) );
  OAI22_X2 U2182 ( .A1(n445), .A2(n16), .B1(n477), .B2(n13), .ZN(n2705) );
  AOI221_X2 U2183 ( .B1(n10), .B2(\registers[9][3] ), .C1(n7), .C2(
        \registers[8][3] ), .A(n2706), .ZN(n2690) );
  OAI22_X2 U2184 ( .A1(n317), .A2(n4), .B1(n349), .B2(n1), .ZN(n2706) );
  NAND4_X2 U2185 ( .A1(n2707), .A2(n2708), .A3(n2709), .A4(n2710), .ZN(N188)
         );
  NOR4_X2 U2186 ( .A1(n2711), .A2(n2712), .A3(n2713), .A4(n2714), .ZN(n2710)
         );
  OAI221_X2 U2187 ( .B1(n542), .B2(n219), .C1(n510), .C2(n216), .A(n2715), 
        .ZN(n2714) );
  AOI22_X2 U2188 ( .A1(n213), .A2(\registers[19][2] ), .B1(n210), .B2(
        \registers[18][2] ), .ZN(n2715) );
  OAI221_X2 U2189 ( .B1(n670), .B2(n207), .C1(n638), .C2(n204), .A(n2716), 
        .ZN(n2713) );
  AOI22_X2 U2190 ( .A1(n201), .A2(\registers[23][2] ), .B1(n198), .B2(
        \registers[22][2] ), .ZN(n2716) );
  OAI221_X2 U2191 ( .B1(n862), .B2(n195), .C1(n830), .C2(n192), .A(n2717), 
        .ZN(n2712) );
  AOI22_X2 U2192 ( .A1(n189), .A2(\registers[25][2] ), .B1(n186), .B2(
        \registers[24][2] ), .ZN(n2717) );
  OAI221_X2 U2193 ( .B1(n990), .B2(n183), .C1(n958), .C2(n180), .A(n2718), 
        .ZN(n2711) );
  AOI22_X2 U2194 ( .A1(n177), .A2(\registers[29][2] ), .B1(n174), .B2(
        \registers[28][2] ), .ZN(n2718) );
  AOI211_X2 U2195 ( .C1(n171), .C2(\registers[1][2] ), .A(n2719), .B(n2720), 
        .ZN(n2709) );
  OAI22_X2 U2196 ( .A1(n62), .A2(n168), .B1(n94), .B2(n165), .ZN(n2720) );
  OAI221_X2 U2197 ( .B1(n158), .B2(n162), .C1(n126), .C2(n31), .A(n2721), .ZN(
        n2719) );
  AOI22_X2 U2198 ( .A1(n28), .A2(\registers[7][2] ), .B1(n25), .B2(
        \registers[6][2] ), .ZN(n2721) );
  AOI221_X2 U2199 ( .B1(n22), .B2(\registers[13][2] ), .C1(n19), .C2(
        \registers[12][2] ), .A(n2722), .ZN(n2708) );
  OAI22_X2 U2200 ( .A1(n446), .A2(n16), .B1(n478), .B2(n13), .ZN(n2722) );
  AOI221_X2 U2201 ( .B1(n10), .B2(\registers[9][2] ), .C1(n7), .C2(
        \registers[8][2] ), .A(n2723), .ZN(n2707) );
  OAI22_X2 U2202 ( .A1(n318), .A2(n4), .B1(n350), .B2(n1), .ZN(n2723) );
  NAND4_X2 U2203 ( .A1(n2724), .A2(n2725), .A3(n2726), .A4(n2727), .ZN(N187)
         );
  NOR4_X2 U2204 ( .A1(n2728), .A2(n2729), .A3(n2730), .A4(n2731), .ZN(n2727)
         );
  OAI221_X2 U2205 ( .B1(n543), .B2(n219), .C1(n511), .C2(n216), .A(n2732), 
        .ZN(n2731) );
  AOI22_X2 U2206 ( .A1(n213), .A2(\registers[19][1] ), .B1(n210), .B2(
        \registers[18][1] ), .ZN(n2732) );
  OAI221_X2 U2207 ( .B1(n671), .B2(n207), .C1(n639), .C2(n204), .A(n2733), 
        .ZN(n2730) );
  AOI22_X2 U2208 ( .A1(n201), .A2(\registers[23][1] ), .B1(n198), .B2(
        \registers[22][1] ), .ZN(n2733) );
  OAI221_X2 U2209 ( .B1(n863), .B2(n195), .C1(n831), .C2(n192), .A(n2734), 
        .ZN(n2729) );
  AOI22_X2 U2210 ( .A1(n189), .A2(\registers[25][1] ), .B1(n186), .B2(
        \registers[24][1] ), .ZN(n2734) );
  OAI221_X2 U2211 ( .B1(n991), .B2(n183), .C1(n959), .C2(n180), .A(n2735), 
        .ZN(n2728) );
  AOI22_X2 U2212 ( .A1(n177), .A2(\registers[29][1] ), .B1(n174), .B2(
        \registers[28][1] ), .ZN(n2735) );
  AOI211_X2 U2213 ( .C1(n171), .C2(\registers[1][1] ), .A(n2736), .B(n2737), 
        .ZN(n2726) );
  OAI22_X2 U2214 ( .A1(n63), .A2(n168), .B1(n95), .B2(n165), .ZN(n2737) );
  OAI221_X2 U2215 ( .B1(n159), .B2(n162), .C1(n127), .C2(n31), .A(n2738), .ZN(
        n2736) );
  AOI22_X2 U2216 ( .A1(n28), .A2(\registers[7][1] ), .B1(n25), .B2(
        \registers[6][1] ), .ZN(n2738) );
  AOI221_X2 U2217 ( .B1(n22), .B2(\registers[13][1] ), .C1(n19), .C2(
        \registers[12][1] ), .A(n2739), .ZN(n2725) );
  OAI22_X2 U2218 ( .A1(n447), .A2(n16), .B1(n479), .B2(n13), .ZN(n2739) );
  AOI221_X2 U2219 ( .B1(n10), .B2(\registers[9][1] ), .C1(n7), .C2(
        \registers[8][1] ), .A(n2740), .ZN(n2724) );
  OAI22_X2 U2220 ( .A1(n319), .A2(n4), .B1(n351), .B2(n1), .ZN(n2740) );
  NAND4_X2 U2221 ( .A1(n2741), .A2(n2742), .A3(n2743), .A4(n2744), .ZN(N186)
         );
  NOR4_X2 U2222 ( .A1(n2745), .A2(n2746), .A3(n2747), .A4(n2748), .ZN(n2744)
         );
  OAI221_X2 U2223 ( .B1(n544), .B2(n219), .C1(n512), .C2(n216), .A(n2749), 
        .ZN(n2748) );
  AOI22_X2 U2224 ( .A1(n213), .A2(\registers[19][0] ), .B1(n210), .B2(
        \registers[18][0] ), .ZN(n2749) );
  AND2_X2 U2225 ( .A1(n2750), .A2(n2751), .ZN(n2195) );
  AND2_X2 U2226 ( .A1(n2752), .A2(n2751), .ZN(n2194) );
  NAND2_X2 U2227 ( .A1(n2750), .A2(n2753), .ZN(n2192) );
  NAND2_X2 U2228 ( .A1(n2752), .A2(n2753), .ZN(n2191) );
  OAI221_X2 U2229 ( .B1(n672), .B2(n207), .C1(n640), .C2(n204), .A(n2754), 
        .ZN(n2747) );
  AOI22_X2 U2230 ( .A1(n201), .A2(\registers[23][0] ), .B1(n198), .B2(
        \registers[22][0] ), .ZN(n2754) );
  AND2_X2 U2231 ( .A1(n2750), .A2(n2755), .ZN(n2200) );
  AND2_X2 U2232 ( .A1(n2752), .A2(n2755), .ZN(n2199) );
  NAND2_X2 U2233 ( .A1(n2750), .A2(n2756), .ZN(n2197) );
  AND2_X2 U2234 ( .A1(n2757), .A2(n3855), .ZN(n2750) );
  NAND2_X2 U2235 ( .A1(n2752), .A2(n2756), .ZN(n2196) );
  AND2_X2 U2236 ( .A1(n2757), .A2(ADD_RD1[0]), .ZN(n2752) );
  AND2_X2 U2237 ( .A1(ADD_RD1[4]), .A2(n3853), .ZN(n2757) );
  OAI221_X2 U2238 ( .B1(n864), .B2(n195), .C1(n832), .C2(n192), .A(n2758), 
        .ZN(n2746) );
  AOI22_X2 U2239 ( .A1(n189), .A2(\registers[25][0] ), .B1(n186), .B2(
        \registers[24][0] ), .ZN(n2758) );
  AND2_X2 U2240 ( .A1(n2753), .A2(n2759), .ZN(n2205) );
  AND2_X2 U2241 ( .A1(n2753), .A2(n2760), .ZN(n2204) );
  NAND2_X2 U2242 ( .A1(n2751), .A2(n2759), .ZN(n2202) );
  NAND2_X2 U2243 ( .A1(n2751), .A2(n2760), .ZN(n2201) );
  OAI221_X2 U2244 ( .B1(n992), .B2(n183), .C1(n960), .C2(n180), .A(n2761), 
        .ZN(n2745) );
  AOI22_X2 U2245 ( .A1(n177), .A2(\registers[29][0] ), .B1(n174), .B2(
        \registers[28][0] ), .ZN(n2761) );
  AND2_X2 U2246 ( .A1(n2756), .A2(n2759), .ZN(n2210) );
  AND2_X2 U2247 ( .A1(n2756), .A2(n2760), .ZN(n2209) );
  NAND2_X2 U2248 ( .A1(n2759), .A2(n2755), .ZN(n2207) );
  AND2_X2 U2249 ( .A1(n2762), .A2(n3855), .ZN(n2759) );
  NAND2_X2 U2250 ( .A1(n2755), .A2(n2760), .ZN(n2206) );
  AND2_X2 U2251 ( .A1(ADD_RD1[0]), .A2(n2762), .ZN(n2760) );
  AND2_X2 U2252 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2762) );
  AOI211_X2 U2253 ( .C1(n171), .C2(\registers[1][0] ), .A(n2763), .B(n2764), 
        .ZN(n2743) );
  OAI22_X2 U2254 ( .A1(n64), .A2(n168), .B1(n96), .B2(n165), .ZN(n2764) );
  NAND2_X2 U2255 ( .A1(n2765), .A2(n2751), .ZN(n2215) );
  NAND2_X2 U2256 ( .A1(n2766), .A2(n2751), .ZN(n2214) );
  OAI221_X2 U2257 ( .B1(n160), .B2(n162), .C1(n128), .C2(n31), .A(n2767), .ZN(
        n2763) );
  AOI22_X2 U2258 ( .A1(n28), .A2(\registers[7][0] ), .B1(n25), .B2(
        \registers[6][0] ), .ZN(n2767) );
  AND2_X2 U2259 ( .A1(n2766), .A2(n2755), .ZN(n2220) );
  AND2_X2 U2260 ( .A1(n2765), .A2(n2755), .ZN(n2219) );
  NAND2_X2 U2261 ( .A1(n2766), .A2(n2756), .ZN(n2217) );
  AND2_X2 U2262 ( .A1(n2768), .A2(n3855), .ZN(n2766) );
  NAND2_X2 U2263 ( .A1(n2765), .A2(n2756), .ZN(n2216) );
  AND2_X2 U2264 ( .A1(n2765), .A2(n2753), .ZN(n2211) );
  AND2_X2 U2265 ( .A1(n2768), .A2(ADD_RD1[0]), .ZN(n2765) );
  NOR2_X2 U2266 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n2768) );
  AOI221_X2 U2267 ( .B1(n22), .B2(\registers[13][0] ), .C1(n19), .C2(
        \registers[12][0] ), .A(n2769), .ZN(n2742) );
  OAI22_X2 U2268 ( .A1(n448), .A2(n16), .B1(n480), .B2(n13), .ZN(n2769) );
  NAND2_X2 U2269 ( .A1(n2770), .A2(n2755), .ZN(n2225) );
  NAND2_X2 U2270 ( .A1(n2771), .A2(n2755), .ZN(n2224) );
  AND2_X2 U2271 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n2755) );
  AND2_X2 U2272 ( .A1(n2771), .A2(n2756), .ZN(n2222) );
  AND2_X2 U2273 ( .A1(n2770), .A2(n2756), .ZN(n2221) );
  AND2_X2 U2274 ( .A1(ADD_RD1[2]), .A2(n3854), .ZN(n2756) );
  AOI221_X2 U2275 ( .B1(n10), .B2(\registers[9][0] ), .C1(n7), .C2(
        \registers[8][0] ), .A(n2772), .ZN(n2741) );
  OAI22_X2 U2276 ( .A1(n320), .A2(n4), .B1(n352), .B2(n1), .ZN(n2772) );
  NAND2_X2 U2277 ( .A1(n2770), .A2(n2751), .ZN(n2230) );
  NAND2_X2 U2278 ( .A1(n2771), .A2(n2751), .ZN(n2229) );
  NOR2_X2 U2279 ( .A1(n3854), .A2(ADD_RD1[2]), .ZN(n2751) );
  AND2_X2 U2280 ( .A1(n2771), .A2(n2753), .ZN(n2227) );
  AND2_X2 U2281 ( .A1(n2773), .A2(n3855), .ZN(n2771) );
  AND2_X2 U2282 ( .A1(n2770), .A2(n2753), .ZN(n2226) );
  NOR2_X2 U2283 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2753) );
  AND2_X2 U2284 ( .A1(n2773), .A2(ADD_RD1[0]), .ZN(n2770) );
  NOR2_X2 U2285 ( .A1(n3853), .A2(ADD_RD1[4]), .ZN(n2773) );
  BUF_X4 U2286 ( .A(n2230), .Z(n1) );
  BUF_X4 U2287 ( .A(n2230), .Z(n2) );
  BUF_X4 U2288 ( .A(n2229), .Z(n4) );
  BUF_X4 U2289 ( .A(n2229), .Z(n5) );
  BUF_X4 U2290 ( .A(n2225), .Z(n13) );
  BUF_X4 U2291 ( .A(n2225), .Z(n14) );
  BUF_X4 U2292 ( .A(n2224), .Z(n16) );
  BUF_X4 U2293 ( .A(n2224), .Z(n17) );
  BUF_X4 U2294 ( .A(n2217), .Z(n31) );
  BUF_X4 U2295 ( .A(n2217), .Z(n32) );
  BUF_X4 U2296 ( .A(n2216), .Z(n163) );
  BUF_X4 U2297 ( .A(n2215), .Z(n165) );
  BUF_X4 U2298 ( .A(n2215), .Z(n166) );
  BUF_X4 U2299 ( .A(n2214), .Z(n168) );
  BUF_X4 U2300 ( .A(n2214), .Z(n169) );
  BUF_X4 U2301 ( .A(n2207), .Z(n180) );
  BUF_X4 U2302 ( .A(n2207), .Z(n181) );
  BUF_X4 U2303 ( .A(n2206), .Z(n184) );
  BUF_X4 U2304 ( .A(n2202), .Z(n192) );
  BUF_X4 U2305 ( .A(n2202), .Z(n193) );
  BUF_X4 U2306 ( .A(n2201), .Z(n196) );
  BUF_X4 U2307 ( .A(n2197), .Z(n204) );
  BUF_X4 U2308 ( .A(n2197), .Z(n205) );
  BUF_X4 U2309 ( .A(n2196), .Z(n208) );
  BUF_X4 U2310 ( .A(n2192), .Z(n216) );
  BUF_X4 U2311 ( .A(n2192), .Z(n217) );
  BUF_X4 U2312 ( .A(n2191), .Z(n220) );
  BUF_X4 U2313 ( .A(n1639), .Z(n222) );
  BUF_X4 U2314 ( .A(n1639), .Z(n223) );
  BUF_X4 U2315 ( .A(n1638), .Z(n225) );
  BUF_X4 U2316 ( .A(n1638), .Z(n226) );
  BUF_X4 U2317 ( .A(n1634), .Z(n234) );
  BUF_X4 U2318 ( .A(n1634), .Z(n235) );
  BUF_X4 U2319 ( .A(n1633), .Z(n237) );
  BUF_X4 U2320 ( .A(n1633), .Z(n238) );
  BUF_X4 U2321 ( .A(n1626), .Z(n252) );
  BUF_X4 U2322 ( .A(n1626), .Z(n253) );
  BUF_X4 U2323 ( .A(n1625), .Z(n256) );
  BUF_X4 U2324 ( .A(n1624), .Z(n258) );
  BUF_X4 U2325 ( .A(n1624), .Z(n259) );
  BUF_X4 U2326 ( .A(n1623), .Z(n261) );
  BUF_X4 U2327 ( .A(n1623), .Z(n262) );
  BUF_X4 U2328 ( .A(n1616), .Z(n273) );
  BUF_X4 U2329 ( .A(n1616), .Z(n274) );
  BUF_X4 U2330 ( .A(n1615), .Z(n277) );
  BUF_X4 U2331 ( .A(n1611), .Z(n285) );
  BUF_X4 U2332 ( .A(n1611), .Z(n286) );
  BUF_X4 U2333 ( .A(n1610), .Z(n353) );
  BUF_X4 U2334 ( .A(n1606), .Z(n361) );
  BUF_X4 U2335 ( .A(n1606), .Z(n362) );
  BUF_X4 U2336 ( .A(n1605), .Z(n365) );
  BUF_X4 U2337 ( .A(n1601), .Z(n373) );
  BUF_X4 U2338 ( .A(n1601), .Z(n374) );
  BUF_X4 U2339 ( .A(n1600), .Z(n377) );
  INV_X2 U2340 ( .A(n388), .ZN(n379) );
  INV_X2 U2341 ( .A(n388), .ZN(n380) );
  INV_X2 U2342 ( .A(n398), .ZN(n389) );
  INV_X2 U2343 ( .A(n398), .ZN(n390) );
  INV_X2 U2344 ( .A(n409), .ZN(n400) );
  INV_X2 U2345 ( .A(n409), .ZN(n401) );
  INV_X2 U2346 ( .A(n548), .ZN(n411) );
  INV_X2 U2347 ( .A(n548), .ZN(n412) );
  INV_X2 U2348 ( .A(n559), .ZN(n550) );
  INV_X2 U2349 ( .A(n559), .ZN(n551) );
  INV_X2 U2350 ( .A(n570), .ZN(n561) );
  INV_X2 U2351 ( .A(n570), .ZN(n562) );
  INV_X2 U2352 ( .A(n580), .ZN(n571) );
  INV_X2 U2353 ( .A(n580), .ZN(n572) );
  INV_X2 U2354 ( .A(n590), .ZN(n581) );
  INV_X2 U2355 ( .A(n590), .ZN(n582) );
  INV_X2 U2356 ( .A(n600), .ZN(n591) );
  INV_X2 U2357 ( .A(n600), .ZN(n592) );
  INV_X2 U2358 ( .A(n674), .ZN(n601) );
  INV_X2 U2359 ( .A(n674), .ZN(n602) );
  INV_X2 U2360 ( .A(n685), .ZN(n676) );
  INV_X2 U2361 ( .A(n685), .ZN(n677) );
  INV_X2 U2362 ( .A(n696), .ZN(n687) );
  INV_X2 U2363 ( .A(n696), .ZN(n688) );
  INV_X2 U2364 ( .A(n706), .ZN(n697) );
  INV_X2 U2365 ( .A(n706), .ZN(n698) );
  INV_X2 U2366 ( .A(n716), .ZN(n707) );
  INV_X2 U2367 ( .A(n716), .ZN(n708) );
  INV_X2 U2368 ( .A(n727), .ZN(n718) );
  INV_X2 U2369 ( .A(n727), .ZN(n719) );
  INV_X2 U2370 ( .A(n738), .ZN(n729) );
  INV_X2 U2371 ( .A(n738), .ZN(n730) );
  INV_X2 U2372 ( .A(n749), .ZN(n740) );
  INV_X2 U2373 ( .A(n749), .ZN(n741) );
  INV_X2 U2374 ( .A(n760), .ZN(n751) );
  INV_X2 U2375 ( .A(n760), .ZN(n752) );
  INV_X2 U2376 ( .A(n770), .ZN(n761) );
  INV_X2 U2377 ( .A(n770), .ZN(n762) );
  INV_X2 U2378 ( .A(n780), .ZN(n771) );
  INV_X2 U2379 ( .A(n780), .ZN(n772) );
  INV_X2 U2380 ( .A(n791), .ZN(n782) );
  INV_X2 U2381 ( .A(n791), .ZN(n783) );
  INV_X2 U2382 ( .A(n866), .ZN(n793) );
  INV_X2 U2383 ( .A(n866), .ZN(n794) );
  INV_X2 U2384 ( .A(n876), .ZN(n867) );
  INV_X2 U2385 ( .A(n876), .ZN(n868) );
  INV_X2 U2386 ( .A(n886), .ZN(n877) );
  INV_X2 U2387 ( .A(n886), .ZN(n878) );
  INV_X2 U2388 ( .A(n896), .ZN(n887) );
  INV_X2 U2389 ( .A(n896), .ZN(n888) );
  INV_X2 U2390 ( .A(n906), .ZN(n897) );
  INV_X2 U2391 ( .A(n906), .ZN(n898) );
  INV_X2 U2392 ( .A(n917), .ZN(n908) );
  INV_X2 U2393 ( .A(n917), .ZN(n909) );
  INV_X2 U2394 ( .A(n928), .ZN(n919) );
  INV_X2 U2395 ( .A(n928), .ZN(n920) );
  INV_X2 U2396 ( .A(n1002), .ZN(n993) );
  INV_X2 U2397 ( .A(n1002), .ZN(n994) );
  INV_X2 U2398 ( .A(n1012), .ZN(n1003) );
  INV_X2 U2399 ( .A(n1012), .ZN(n1004) );
  INV_X2 U2400 ( .A(n1023), .ZN(n1014) );
  INV_X2 U2401 ( .A(n1023), .ZN(n1015) );
  INV_X2 U2402 ( .A(n1023), .ZN(n1016) );
  CLKBUF_X3 U2403 ( .A(n2230), .Z(n3) );
  CLKBUF_X3 U2404 ( .A(n2229), .Z(n6) );
  CLKBUF_X3 U2405 ( .A(n2227), .Z(n7) );
  CLKBUF_X3 U2406 ( .A(n2227), .Z(n8) );
  CLKBUF_X3 U2407 ( .A(n2227), .Z(n9) );
  CLKBUF_X3 U2408 ( .A(n2226), .Z(n10) );
  CLKBUF_X3 U2409 ( .A(n2226), .Z(n11) );
  CLKBUF_X3 U2410 ( .A(n2226), .Z(n12) );
  CLKBUF_X3 U2411 ( .A(n2225), .Z(n15) );
  CLKBUF_X3 U2412 ( .A(n2224), .Z(n18) );
  CLKBUF_X3 U2413 ( .A(n2222), .Z(n19) );
  CLKBUF_X3 U2414 ( .A(n2222), .Z(n20) );
  CLKBUF_X3 U2415 ( .A(n2222), .Z(n21) );
  CLKBUF_X3 U2416 ( .A(n2221), .Z(n22) );
  CLKBUF_X3 U2417 ( .A(n2221), .Z(n23) );
  CLKBUF_X3 U2418 ( .A(n2221), .Z(n24) );
  CLKBUF_X3 U2419 ( .A(n2220), .Z(n25) );
  CLKBUF_X3 U2420 ( .A(n2220), .Z(n26) );
  CLKBUF_X3 U2421 ( .A(n2220), .Z(n27) );
  CLKBUF_X3 U2422 ( .A(n2219), .Z(n28) );
  CLKBUF_X3 U2423 ( .A(n2219), .Z(n29) );
  CLKBUF_X3 U2424 ( .A(n2219), .Z(n30) );
  CLKBUF_X3 U2425 ( .A(n2217), .Z(n161) );
  CLKBUF_X3 U2426 ( .A(n2216), .Z(n162) );
  CLKBUF_X3 U2427 ( .A(n2216), .Z(n164) );
  CLKBUF_X3 U2428 ( .A(n2215), .Z(n167) );
  CLKBUF_X3 U2429 ( .A(n2214), .Z(n170) );
  CLKBUF_X3 U2430 ( .A(n2211), .Z(n171) );
  CLKBUF_X3 U2431 ( .A(n2211), .Z(n172) );
  CLKBUF_X3 U2432 ( .A(n2211), .Z(n173) );
  CLKBUF_X3 U2433 ( .A(n2210), .Z(n174) );
  CLKBUF_X3 U2434 ( .A(n2210), .Z(n175) );
  CLKBUF_X3 U2435 ( .A(n2210), .Z(n176) );
  CLKBUF_X3 U2436 ( .A(n2209), .Z(n177) );
  CLKBUF_X3 U2437 ( .A(n2209), .Z(n178) );
  CLKBUF_X3 U2438 ( .A(n2209), .Z(n179) );
  CLKBUF_X3 U2439 ( .A(n2207), .Z(n182) );
  CLKBUF_X3 U2440 ( .A(n2206), .Z(n183) );
  CLKBUF_X3 U2441 ( .A(n2206), .Z(n185) );
  CLKBUF_X3 U2442 ( .A(n2205), .Z(n186) );
  CLKBUF_X3 U2443 ( .A(n2205), .Z(n187) );
  CLKBUF_X3 U2444 ( .A(n2205), .Z(n188) );
  CLKBUF_X3 U2445 ( .A(n2204), .Z(n189) );
  CLKBUF_X3 U2446 ( .A(n2204), .Z(n190) );
  CLKBUF_X3 U2447 ( .A(n2204), .Z(n191) );
  CLKBUF_X3 U2448 ( .A(n2202), .Z(n194) );
  CLKBUF_X3 U2449 ( .A(n2201), .Z(n195) );
  CLKBUF_X3 U2450 ( .A(n2201), .Z(n197) );
  CLKBUF_X3 U2451 ( .A(n2200), .Z(n198) );
  CLKBUF_X3 U2452 ( .A(n2200), .Z(n199) );
  CLKBUF_X3 U2453 ( .A(n2200), .Z(n200) );
  CLKBUF_X3 U2454 ( .A(n2199), .Z(n201) );
  CLKBUF_X3 U2455 ( .A(n2199), .Z(n202) );
  CLKBUF_X3 U2456 ( .A(n2199), .Z(n203) );
  CLKBUF_X3 U2457 ( .A(n2197), .Z(n206) );
  CLKBUF_X3 U2458 ( .A(n2196), .Z(n207) );
  CLKBUF_X3 U2459 ( .A(n2196), .Z(n209) );
  CLKBUF_X3 U2460 ( .A(n2195), .Z(n210) );
  CLKBUF_X3 U2461 ( .A(n2195), .Z(n211) );
  CLKBUF_X3 U2462 ( .A(n2195), .Z(n212) );
  CLKBUF_X3 U2463 ( .A(n2194), .Z(n213) );
  CLKBUF_X3 U2464 ( .A(n2194), .Z(n214) );
  CLKBUF_X3 U2465 ( .A(n2194), .Z(n215) );
  CLKBUF_X3 U2466 ( .A(n2192), .Z(n218) );
  CLKBUF_X3 U2467 ( .A(n2191), .Z(n219) );
  CLKBUF_X3 U2468 ( .A(n2191), .Z(n221) );
  CLKBUF_X3 U2469 ( .A(n1639), .Z(n224) );
  CLKBUF_X3 U2470 ( .A(n1638), .Z(n227) );
  CLKBUF_X3 U2471 ( .A(n1636), .Z(n228) );
  CLKBUF_X3 U2472 ( .A(n1636), .Z(n229) );
  CLKBUF_X3 U2473 ( .A(n1636), .Z(n230) );
  CLKBUF_X3 U2474 ( .A(n1635), .Z(n231) );
  CLKBUF_X3 U2475 ( .A(n1635), .Z(n232) );
  CLKBUF_X3 U2476 ( .A(n1635), .Z(n233) );
  CLKBUF_X3 U2477 ( .A(n1634), .Z(n236) );
  CLKBUF_X3 U2478 ( .A(n1633), .Z(n239) );
  CLKBUF_X3 U2479 ( .A(n1631), .Z(n240) );
  CLKBUF_X3 U2480 ( .A(n1631), .Z(n241) );
  CLKBUF_X3 U2481 ( .A(n1631), .Z(n242) );
  CLKBUF_X3 U2482 ( .A(n1630), .Z(n243) );
  CLKBUF_X3 U2483 ( .A(n1630), .Z(n244) );
  CLKBUF_X3 U2484 ( .A(n1630), .Z(n245) );
  CLKBUF_X3 U2485 ( .A(n1629), .Z(n246) );
  CLKBUF_X3 U2486 ( .A(n1629), .Z(n247) );
  CLKBUF_X3 U2487 ( .A(n1629), .Z(n248) );
  CLKBUF_X3 U2488 ( .A(n1628), .Z(n249) );
  CLKBUF_X3 U2489 ( .A(n1628), .Z(n250) );
  CLKBUF_X3 U2490 ( .A(n1628), .Z(n251) );
  CLKBUF_X3 U2491 ( .A(n1626), .Z(n254) );
  CLKBUF_X3 U2492 ( .A(n1625), .Z(n255) );
  CLKBUF_X3 U2493 ( .A(n1625), .Z(n257) );
  CLKBUF_X3 U2494 ( .A(n1624), .Z(n260) );
  CLKBUF_X3 U2495 ( .A(n1623), .Z(n263) );
  CLKBUF_X3 U2496 ( .A(n1620), .Z(n264) );
  CLKBUF_X3 U2497 ( .A(n1620), .Z(n265) );
  CLKBUF_X3 U2498 ( .A(n1620), .Z(n266) );
  CLKBUF_X3 U2499 ( .A(n1619), .Z(n267) );
  CLKBUF_X3 U2500 ( .A(n1619), .Z(n268) );
  CLKBUF_X3 U2501 ( .A(n1619), .Z(n269) );
  CLKBUF_X3 U2502 ( .A(n1618), .Z(n270) );
  CLKBUF_X3 U2503 ( .A(n1618), .Z(n271) );
  CLKBUF_X3 U2504 ( .A(n1618), .Z(n272) );
  CLKBUF_X3 U2505 ( .A(n1616), .Z(n275) );
  CLKBUF_X3 U2506 ( .A(n1615), .Z(n276) );
  CLKBUF_X3 U2507 ( .A(n1615), .Z(n278) );
  CLKBUF_X3 U2508 ( .A(n1614), .Z(n279) );
  CLKBUF_X3 U2509 ( .A(n1614), .Z(n280) );
  CLKBUF_X3 U2510 ( .A(n1614), .Z(n281) );
  CLKBUF_X3 U2511 ( .A(n1613), .Z(n282) );
  CLKBUF_X3 U2512 ( .A(n1613), .Z(n283) );
  CLKBUF_X3 U2513 ( .A(n1613), .Z(n284) );
  CLKBUF_X3 U2514 ( .A(n1611), .Z(n287) );
  CLKBUF_X3 U2515 ( .A(n1610), .Z(n288) );
  CLKBUF_X3 U2516 ( .A(n1610), .Z(n354) );
  CLKBUF_X3 U2517 ( .A(n1609), .Z(n355) );
  CLKBUF_X3 U2518 ( .A(n1609), .Z(n356) );
  CLKBUF_X3 U2519 ( .A(n1609), .Z(n357) );
  CLKBUF_X3 U2520 ( .A(n1608), .Z(n358) );
  CLKBUF_X3 U2521 ( .A(n1608), .Z(n359) );
  CLKBUF_X3 U2522 ( .A(n1608), .Z(n360) );
  CLKBUF_X3 U2523 ( .A(n1606), .Z(n363) );
  CLKBUF_X3 U2524 ( .A(n1605), .Z(n364) );
  CLKBUF_X3 U2525 ( .A(n1605), .Z(n366) );
  CLKBUF_X3 U2526 ( .A(n1604), .Z(n367) );
  CLKBUF_X3 U2527 ( .A(n1604), .Z(n368) );
  CLKBUF_X3 U2528 ( .A(n1604), .Z(n369) );
  CLKBUF_X3 U2529 ( .A(n1603), .Z(n370) );
  CLKBUF_X3 U2530 ( .A(n1603), .Z(n371) );
  CLKBUF_X3 U2531 ( .A(n1603), .Z(n372) );
  CLKBUF_X3 U2532 ( .A(n1601), .Z(n375) );
  CLKBUF_X3 U2533 ( .A(n1600), .Z(n376) );
  CLKBUF_X3 U2534 ( .A(n1600), .Z(n378) );
  INV_X1 U2535 ( .A(n388), .ZN(n381) );
  CLKBUF_X3 U2536 ( .A(n1560), .Z(n382) );
  CLKBUF_X3 U2537 ( .A(n1560), .Z(n383) );
  CLKBUF_X3 U2538 ( .A(n1560), .Z(n384) );
  CLKBUF_X3 U2539 ( .A(n1560), .Z(n385) );
  CLKBUF_X3 U2540 ( .A(n1560), .Z(n386) );
  CLKBUF_X3 U2541 ( .A(n1560), .Z(n387) );
  CLKBUF_X3 U2542 ( .A(n1560), .Z(n388) );
  INV_X1 U2543 ( .A(n398), .ZN(n391) );
  CLKBUF_X3 U2544 ( .A(n399), .Z(n392) );
  CLKBUF_X3 U2545 ( .A(n399), .Z(n393) );
  CLKBUF_X3 U2546 ( .A(n399), .Z(n394) );
  CLKBUF_X3 U2547 ( .A(n399), .Z(n395) );
  CLKBUF_X3 U2548 ( .A(n399), .Z(n396) );
  CLKBUF_X3 U2549 ( .A(n399), .Z(n397) );
  CLKBUF_X3 U2550 ( .A(n399), .Z(n398) );
  INV_X16 U2551 ( .A(n1558), .ZN(n399) );
  INV_X1 U2552 ( .A(n409), .ZN(n402) );
  CLKBUF_X3 U2553 ( .A(n410), .Z(n403) );
  CLKBUF_X3 U2554 ( .A(n410), .Z(n404) );
  CLKBUF_X3 U2555 ( .A(n410), .Z(n405) );
  CLKBUF_X3 U2556 ( .A(n410), .Z(n406) );
  CLKBUF_X3 U2557 ( .A(n410), .Z(n407) );
  CLKBUF_X3 U2558 ( .A(n410), .Z(n408) );
  CLKBUF_X3 U2559 ( .A(n410), .Z(n409) );
  INV_X16 U2560 ( .A(n1557), .ZN(n410) );
  INV_X1 U2561 ( .A(n548), .ZN(n413) );
  CLKBUF_X3 U2562 ( .A(n549), .Z(n414) );
  CLKBUF_X3 U2563 ( .A(n549), .Z(n415) );
  CLKBUF_X3 U2564 ( .A(n549), .Z(n416) );
  CLKBUF_X3 U2565 ( .A(n549), .Z(n545) );
  CLKBUF_X3 U2566 ( .A(n549), .Z(n546) );
  CLKBUF_X3 U2567 ( .A(n549), .Z(n547) );
  CLKBUF_X3 U2568 ( .A(n549), .Z(n548) );
  INV_X16 U2569 ( .A(n1556), .ZN(n549) );
  INV_X1 U2570 ( .A(n559), .ZN(n552) );
  CLKBUF_X3 U2571 ( .A(n560), .Z(n553) );
  CLKBUF_X3 U2572 ( .A(n560), .Z(n554) );
  CLKBUF_X3 U2573 ( .A(n560), .Z(n555) );
  CLKBUF_X3 U2574 ( .A(n560), .Z(n556) );
  CLKBUF_X3 U2575 ( .A(n560), .Z(n557) );
  CLKBUF_X3 U2576 ( .A(n560), .Z(n558) );
  CLKBUF_X3 U2577 ( .A(n560), .Z(n559) );
  INV_X16 U2578 ( .A(n1555), .ZN(n560) );
  INV_X1 U2579 ( .A(n570), .ZN(n563) );
  CLKBUF_X3 U2580 ( .A(n1523), .Z(n564) );
  CLKBUF_X3 U2581 ( .A(n1523), .Z(n565) );
  CLKBUF_X3 U2582 ( .A(n1523), .Z(n566) );
  CLKBUF_X3 U2583 ( .A(n1523), .Z(n567) );
  CLKBUF_X3 U2584 ( .A(n1523), .Z(n568) );
  CLKBUF_X3 U2585 ( .A(n1523), .Z(n569) );
  CLKBUF_X3 U2586 ( .A(n1523), .Z(n570) );
  INV_X1 U2587 ( .A(n580), .ZN(n573) );
  CLKBUF_X3 U2588 ( .A(n1489), .Z(n574) );
  CLKBUF_X3 U2589 ( .A(n1489), .Z(n575) );
  CLKBUF_X3 U2590 ( .A(n1489), .Z(n576) );
  CLKBUF_X3 U2591 ( .A(n1489), .Z(n577) );
  CLKBUF_X3 U2592 ( .A(n1489), .Z(n578) );
  CLKBUF_X3 U2593 ( .A(n1489), .Z(n579) );
  CLKBUF_X3 U2594 ( .A(n1489), .Z(n580) );
  INV_X1 U2595 ( .A(n590), .ZN(n583) );
  CLKBUF_X3 U2596 ( .A(n1456), .Z(n584) );
  CLKBUF_X3 U2597 ( .A(n1456), .Z(n585) );
  CLKBUF_X3 U2598 ( .A(n1456), .Z(n586) );
  CLKBUF_X3 U2599 ( .A(n1456), .Z(n587) );
  CLKBUF_X3 U2600 ( .A(n1456), .Z(n588) );
  CLKBUF_X3 U2601 ( .A(n1456), .Z(n589) );
  CLKBUF_X3 U2602 ( .A(n1456), .Z(n590) );
  INV_X1 U2603 ( .A(n600), .ZN(n593) );
  CLKBUF_X3 U2604 ( .A(n1423), .Z(n594) );
  CLKBUF_X3 U2605 ( .A(n1423), .Z(n595) );
  CLKBUF_X3 U2606 ( .A(n1423), .Z(n596) );
  CLKBUF_X3 U2607 ( .A(n1423), .Z(n597) );
  CLKBUF_X3 U2608 ( .A(n1423), .Z(n598) );
  CLKBUF_X3 U2609 ( .A(n1423), .Z(n599) );
  CLKBUF_X3 U2610 ( .A(n1423), .Z(n600) );
  INV_X1 U2611 ( .A(n674), .ZN(n603) );
  CLKBUF_X3 U2612 ( .A(n675), .Z(n604) );
  CLKBUF_X3 U2613 ( .A(n675), .Z(n605) );
  CLKBUF_X3 U2614 ( .A(n675), .Z(n606) );
  CLKBUF_X3 U2615 ( .A(n675), .Z(n607) );
  CLKBUF_X3 U2616 ( .A(n675), .Z(n608) );
  CLKBUF_X3 U2617 ( .A(n675), .Z(n673) );
  CLKBUF_X3 U2618 ( .A(n675), .Z(n674) );
  INV_X16 U2619 ( .A(n1421), .ZN(n675) );
  INV_X1 U2620 ( .A(n685), .ZN(n678) );
  CLKBUF_X3 U2621 ( .A(n686), .Z(n679) );
  CLKBUF_X3 U2622 ( .A(n686), .Z(n680) );
  CLKBUF_X3 U2623 ( .A(n686), .Z(n681) );
  CLKBUF_X3 U2624 ( .A(n686), .Z(n682) );
  CLKBUF_X3 U2625 ( .A(n686), .Z(n683) );
  CLKBUF_X3 U2626 ( .A(n686), .Z(n684) );
  CLKBUF_X3 U2627 ( .A(n686), .Z(n685) );
  INV_X16 U2628 ( .A(n1420), .ZN(n686) );
  INV_X1 U2629 ( .A(n696), .ZN(n689) );
  CLKBUF_X3 U2630 ( .A(n1388), .Z(n690) );
  CLKBUF_X3 U2631 ( .A(n1388), .Z(n691) );
  CLKBUF_X3 U2632 ( .A(n1388), .Z(n692) );
  CLKBUF_X3 U2633 ( .A(n1388), .Z(n693) );
  CLKBUF_X3 U2634 ( .A(n1388), .Z(n694) );
  CLKBUF_X3 U2635 ( .A(n1388), .Z(n695) );
  CLKBUF_X3 U2636 ( .A(n1388), .Z(n696) );
  INV_X1 U2637 ( .A(n706), .ZN(n699) );
  CLKBUF_X3 U2638 ( .A(n1355), .Z(n700) );
  CLKBUF_X3 U2639 ( .A(n1355), .Z(n701) );
  CLKBUF_X3 U2640 ( .A(n1355), .Z(n702) );
  CLKBUF_X3 U2641 ( .A(n1355), .Z(n703) );
  CLKBUF_X3 U2642 ( .A(n1355), .Z(n704) );
  CLKBUF_X3 U2643 ( .A(n1355), .Z(n705) );
  CLKBUF_X3 U2644 ( .A(n1355), .Z(n706) );
  INV_X1 U2645 ( .A(n716), .ZN(n709) );
  CLKBUF_X3 U2646 ( .A(n717), .Z(n710) );
  CLKBUF_X3 U2647 ( .A(n717), .Z(n711) );
  CLKBUF_X3 U2648 ( .A(n717), .Z(n712) );
  CLKBUF_X3 U2649 ( .A(n717), .Z(n713) );
  CLKBUF_X3 U2650 ( .A(n717), .Z(n714) );
  CLKBUF_X3 U2651 ( .A(n717), .Z(n715) );
  CLKBUF_X3 U2652 ( .A(n717), .Z(n716) );
  INV_X16 U2653 ( .A(n1353), .ZN(n717) );
  INV_X1 U2654 ( .A(n727), .ZN(n720) );
  CLKBUF_X3 U2655 ( .A(n728), .Z(n721) );
  CLKBUF_X3 U2656 ( .A(n728), .Z(n722) );
  CLKBUF_X3 U2657 ( .A(n728), .Z(n723) );
  CLKBUF_X3 U2658 ( .A(n728), .Z(n724) );
  CLKBUF_X3 U2659 ( .A(n728), .Z(n725) );
  CLKBUF_X3 U2660 ( .A(n728), .Z(n726) );
  CLKBUF_X3 U2661 ( .A(n728), .Z(n727) );
  INV_X16 U2662 ( .A(n1351), .ZN(n728) );
  INV_X1 U2663 ( .A(n738), .ZN(n731) );
  CLKBUF_X3 U2664 ( .A(n739), .Z(n732) );
  CLKBUF_X3 U2665 ( .A(n739), .Z(n733) );
  CLKBUF_X3 U2666 ( .A(n739), .Z(n734) );
  CLKBUF_X3 U2667 ( .A(n739), .Z(n735) );
  CLKBUF_X3 U2668 ( .A(n739), .Z(n736) );
  CLKBUF_X3 U2669 ( .A(n739), .Z(n737) );
  CLKBUF_X3 U2670 ( .A(n739), .Z(n738) );
  INV_X16 U2671 ( .A(n1350), .ZN(n739) );
  INV_X1 U2672 ( .A(n749), .ZN(n742) );
  CLKBUF_X3 U2673 ( .A(n750), .Z(n743) );
  CLKBUF_X3 U2674 ( .A(n750), .Z(n744) );
  CLKBUF_X3 U2675 ( .A(n750), .Z(n745) );
  CLKBUF_X3 U2676 ( .A(n750), .Z(n746) );
  CLKBUF_X3 U2677 ( .A(n750), .Z(n747) );
  CLKBUF_X3 U2678 ( .A(n750), .Z(n748) );
  CLKBUF_X3 U2679 ( .A(n750), .Z(n749) );
  INV_X16 U2680 ( .A(n1349), .ZN(n750) );
  INV_X1 U2681 ( .A(n760), .ZN(n753) );
  CLKBUF_X3 U2682 ( .A(n1317), .Z(n754) );
  CLKBUF_X3 U2683 ( .A(n1317), .Z(n755) );
  CLKBUF_X3 U2684 ( .A(n1317), .Z(n756) );
  CLKBUF_X3 U2685 ( .A(n1317), .Z(n757) );
  CLKBUF_X3 U2686 ( .A(n1317), .Z(n758) );
  CLKBUF_X3 U2687 ( .A(n1317), .Z(n759) );
  CLKBUF_X3 U2688 ( .A(n1317), .Z(n760) );
  INV_X1 U2689 ( .A(n770), .ZN(n763) );
  CLKBUF_X3 U2690 ( .A(n1284), .Z(n764) );
  CLKBUF_X3 U2691 ( .A(n1284), .Z(n765) );
  CLKBUF_X3 U2692 ( .A(n1284), .Z(n766) );
  CLKBUF_X3 U2693 ( .A(n1284), .Z(n767) );
  CLKBUF_X3 U2694 ( .A(n1284), .Z(n768) );
  CLKBUF_X3 U2695 ( .A(n1284), .Z(n769) );
  CLKBUF_X3 U2696 ( .A(n1284), .Z(n770) );
  INV_X1 U2697 ( .A(n780), .ZN(n773) );
  CLKBUF_X3 U2698 ( .A(n781), .Z(n774) );
  CLKBUF_X3 U2699 ( .A(n781), .Z(n775) );
  CLKBUF_X3 U2700 ( .A(n781), .Z(n776) );
  CLKBUF_X3 U2701 ( .A(n781), .Z(n777) );
  CLKBUF_X3 U2702 ( .A(n781), .Z(n778) );
  CLKBUF_X3 U2703 ( .A(n781), .Z(n779) );
  CLKBUF_X3 U2704 ( .A(n781), .Z(n780) );
  INV_X16 U2705 ( .A(n1282), .ZN(n781) );
  INV_X1 U2706 ( .A(n791), .ZN(n784) );
  CLKBUF_X3 U2707 ( .A(n792), .Z(n785) );
  CLKBUF_X3 U2708 ( .A(n792), .Z(n786) );
  CLKBUF_X3 U2709 ( .A(n792), .Z(n787) );
  CLKBUF_X3 U2710 ( .A(n792), .Z(n788) );
  CLKBUF_X3 U2711 ( .A(n792), .Z(n789) );
  CLKBUF_X3 U2712 ( .A(n792), .Z(n790) );
  CLKBUF_X3 U2713 ( .A(n792), .Z(n791) );
  INV_X16 U2714 ( .A(n1281), .ZN(n792) );
  INV_X1 U2715 ( .A(n866), .ZN(n795) );
  CLKBUF_X3 U2716 ( .A(n1249), .Z(n796) );
  CLKBUF_X3 U2717 ( .A(n1249), .Z(n797) );
  CLKBUF_X3 U2718 ( .A(n1249), .Z(n798) );
  CLKBUF_X3 U2719 ( .A(n1249), .Z(n799) );
  CLKBUF_X3 U2720 ( .A(n1249), .Z(n800) );
  CLKBUF_X3 U2721 ( .A(n1249), .Z(n865) );
  CLKBUF_X3 U2722 ( .A(n1249), .Z(n866) );
  INV_X1 U2723 ( .A(n876), .ZN(n869) );
  CLKBUF_X3 U2724 ( .A(n1215), .Z(n870) );
  CLKBUF_X3 U2725 ( .A(n1215), .Z(n871) );
  CLKBUF_X3 U2726 ( .A(n1215), .Z(n872) );
  CLKBUF_X3 U2727 ( .A(n1215), .Z(n873) );
  CLKBUF_X3 U2728 ( .A(n1215), .Z(n874) );
  CLKBUF_X3 U2729 ( .A(n1215), .Z(n875) );
  CLKBUF_X3 U2730 ( .A(n1215), .Z(n876) );
  INV_X1 U2731 ( .A(n886), .ZN(n879) );
  CLKBUF_X3 U2732 ( .A(n1180), .Z(n880) );
  CLKBUF_X3 U2733 ( .A(n1180), .Z(n881) );
  CLKBUF_X3 U2734 ( .A(n1180), .Z(n882) );
  CLKBUF_X3 U2735 ( .A(n1180), .Z(n883) );
  CLKBUF_X3 U2736 ( .A(n1180), .Z(n884) );
  CLKBUF_X3 U2737 ( .A(n1180), .Z(n885) );
  CLKBUF_X3 U2738 ( .A(n1180), .Z(n886) );
  INV_X1 U2739 ( .A(n896), .ZN(n889) );
  CLKBUF_X3 U2740 ( .A(n1146), .Z(n890) );
  CLKBUF_X3 U2741 ( .A(n1146), .Z(n891) );
  CLKBUF_X3 U2742 ( .A(n1146), .Z(n892) );
  CLKBUF_X3 U2743 ( .A(n1146), .Z(n893) );
  CLKBUF_X3 U2744 ( .A(n1146), .Z(n894) );
  CLKBUF_X3 U2745 ( .A(n1146), .Z(n895) );
  CLKBUF_X3 U2746 ( .A(n1146), .Z(n896) );
  INV_X1 U2747 ( .A(n906), .ZN(n899) );
  CLKBUF_X3 U2748 ( .A(n907), .Z(n900) );
  CLKBUF_X3 U2749 ( .A(n907), .Z(n901) );
  CLKBUF_X3 U2750 ( .A(n907), .Z(n902) );
  CLKBUF_X3 U2751 ( .A(n907), .Z(n903) );
  CLKBUF_X3 U2752 ( .A(n907), .Z(n904) );
  CLKBUF_X3 U2753 ( .A(n907), .Z(n905) );
  CLKBUF_X3 U2754 ( .A(n907), .Z(n906) );
  INV_X16 U2755 ( .A(n1143), .ZN(n907) );
  INV_X1 U2756 ( .A(n917), .ZN(n910) );
  CLKBUF_X3 U2757 ( .A(n918), .Z(n911) );
  CLKBUF_X3 U2758 ( .A(n918), .Z(n912) );
  CLKBUF_X3 U2759 ( .A(n918), .Z(n913) );
  CLKBUF_X3 U2760 ( .A(n918), .Z(n914) );
  CLKBUF_X3 U2761 ( .A(n918), .Z(n915) );
  CLKBUF_X3 U2762 ( .A(n918), .Z(n916) );
  CLKBUF_X3 U2763 ( .A(n918), .Z(n917) );
  INV_X16 U2764 ( .A(n1141), .ZN(n918) );
  INV_X1 U2765 ( .A(n928), .ZN(n921) );
  CLKBUF_X3 U2766 ( .A(n1108), .Z(n922) );
  CLKBUF_X3 U2767 ( .A(n1108), .Z(n923) );
  CLKBUF_X3 U2768 ( .A(n1108), .Z(n924) );
  CLKBUF_X3 U2769 ( .A(n1108), .Z(n925) );
  CLKBUF_X3 U2770 ( .A(n1108), .Z(n926) );
  CLKBUF_X3 U2771 ( .A(n1108), .Z(n927) );
  CLKBUF_X3 U2772 ( .A(n1108), .Z(n928) );
  INV_X1 U2773 ( .A(n1002), .ZN(n995) );
  CLKBUF_X3 U2774 ( .A(n1074), .Z(n996) );
  CLKBUF_X3 U2775 ( .A(n1074), .Z(n997) );
  CLKBUF_X3 U2776 ( .A(n1074), .Z(n998) );
  CLKBUF_X3 U2777 ( .A(n1074), .Z(n999) );
  CLKBUF_X3 U2778 ( .A(n1074), .Z(n1000) );
  CLKBUF_X3 U2779 ( .A(n1074), .Z(n1001) );
  CLKBUF_X3 U2780 ( .A(n1074), .Z(n1002) );
  INV_X1 U2781 ( .A(n1012), .ZN(n1005) );
  CLKBUF_X3 U2782 ( .A(n1013), .Z(n1006) );
  CLKBUF_X3 U2783 ( .A(n1013), .Z(n1007) );
  CLKBUF_X3 U2784 ( .A(n1013), .Z(n1008) );
  CLKBUF_X3 U2785 ( .A(n1013), .Z(n1009) );
  CLKBUF_X3 U2786 ( .A(n1013), .Z(n1010) );
  CLKBUF_X3 U2787 ( .A(n1013), .Z(n1011) );
  CLKBUF_X3 U2788 ( .A(n1013), .Z(n1012) );
  INV_X16 U2789 ( .A(n1071), .ZN(n1013) );
  CLKBUF_X3 U2790 ( .A(n1068), .Z(n1017) );
  CLKBUF_X3 U2791 ( .A(n1068), .Z(n1018) );
  CLKBUF_X3 U2792 ( .A(n1068), .Z(n1019) );
  CLKBUF_X3 U2793 ( .A(n1068), .Z(n1020) );
  CLKBUF_X3 U2794 ( .A(n1068), .Z(n1021) );
  CLKBUF_X3 U2795 ( .A(n1068), .Z(n1022) );
  CLKBUF_X3 U2796 ( .A(n1068), .Z(n1023) );
  CLKBUF_X1 U2797 ( .A(N218), .Z(n1024) );
  CLKBUF_X1 U2798 ( .A(N218), .Z(n1025) );
  CLKBUF_X1 U2799 ( .A(N218), .Z(n1026) );
  CLKBUF_X1 U2800 ( .A(N218), .Z(n1027) );
  CLKBUF_X1 U2801 ( .A(N83), .Z(n1028) );
  CLKBUF_X1 U2802 ( .A(N83), .Z(n1029) );
  CLKBUF_X1 U2803 ( .A(N83), .Z(n1030) );
  CLKBUF_X1 U2804 ( .A(N83), .Z(n1031) );
  CLKBUF_X2 U2805 ( .A(n1042), .Z(n1032) );
  CLKBUF_X2 U2806 ( .A(n1042), .Z(n1033) );
  CLKBUF_X2 U2807 ( .A(n1041), .Z(n1034) );
  CLKBUF_X2 U2808 ( .A(n1041), .Z(n1035) );
  CLKBUF_X2 U2809 ( .A(n1041), .Z(n1036) );
  CLKBUF_X2 U2810 ( .A(n1040), .Z(n1037) );
  CLKBUF_X2 U2811 ( .A(n1040), .Z(n1038) );
  CLKBUF_X2 U2812 ( .A(n1040), .Z(n1039) );
  CLKBUF_X3 U2813 ( .A(RST_AN), .Z(n1040) );
  CLKBUF_X3 U2814 ( .A(RST_AN), .Z(n1041) );
  CLKBUF_X3 U2815 ( .A(RST_AN), .Z(n1042) );
  CLKBUF_X1 U2816 ( .A(n3367), .Z(n1043) );
  CLKBUF_X1 U2817 ( .A(n3366), .Z(n1044) );
  CLKBUF_X1 U2818 ( .A(n3366), .Z(n1045) );
  CLKBUF_X1 U2819 ( .A(n3366), .Z(n1046) );
  CLKBUF_X1 U2820 ( .A(n3366), .Z(n1047) );
  CLKBUF_X1 U2821 ( .A(n3366), .Z(n1048) );
  CLKBUF_X1 U2822 ( .A(n3366), .Z(n1049) );
  CLKBUF_X1 U2823 ( .A(n3365), .Z(n1050) );
  CLKBUF_X1 U2824 ( .A(n3365), .Z(n1051) );
  CLKBUF_X1 U2825 ( .A(n3365), .Z(n1052) );
  CLKBUF_X1 U2826 ( .A(n3365), .Z(n1053) );
  CLKBUF_X1 U2827 ( .A(n3365), .Z(n1054) );
  CLKBUF_X1 U2828 ( .A(n3365), .Z(n1055) );
  CLKBUF_X1 U2829 ( .A(n3364), .Z(n1056) );
  CLKBUF_X1 U2830 ( .A(n3364), .Z(n1057) );
  CLKBUF_X1 U2831 ( .A(n3364), .Z(n1058) );
  CLKBUF_X1 U2832 ( .A(n3364), .Z(n1059) );
  CLKBUF_X1 U2833 ( .A(n3364), .Z(n1060) );
  CLKBUF_X1 U2834 ( .A(n3364), .Z(n1061) );
  CLKBUF_X1 U2835 ( .A(n3363), .Z(n1062) );
  CLKBUF_X1 U2836 ( .A(n3363), .Z(n1063) );
  CLKBUF_X1 U2837 ( .A(n3363), .Z(n1064) );
  CLKBUF_X1 U2838 ( .A(n3363), .Z(n1065) );
  CLKBUF_X1 U2839 ( .A(n3363), .Z(n1066) );
  CLKBUF_X1 U2840 ( .A(n3363), .Z(n1067) );
  CLKBUF_X1 U2841 ( .A(n3362), .Z(n3286) );
  CLKBUF_X1 U2842 ( .A(n3362), .Z(n3287) );
  CLKBUF_X1 U2843 ( .A(n3362), .Z(n3288) );
  CLKBUF_X1 U2844 ( .A(n3362), .Z(n3289) );
  CLKBUF_X1 U2845 ( .A(n3362), .Z(n3290) );
  CLKBUF_X1 U2846 ( .A(n3362), .Z(n3291) );
  CLKBUF_X1 U2847 ( .A(n3361), .Z(n3292) );
  CLKBUF_X1 U2848 ( .A(n3361), .Z(n3293) );
  CLKBUF_X1 U2849 ( .A(n3361), .Z(n3294) );
  CLKBUF_X1 U2850 ( .A(n3361), .Z(n3295) );
  CLKBUF_X1 U2851 ( .A(n3361), .Z(n3296) );
  CLKBUF_X1 U2852 ( .A(n3361), .Z(n3297) );
  CLKBUF_X1 U2853 ( .A(n3360), .Z(n3298) );
  CLKBUF_X1 U2854 ( .A(n3360), .Z(n3299) );
  CLKBUF_X1 U2855 ( .A(n3360), .Z(n3300) );
  CLKBUF_X1 U2856 ( .A(n3360), .Z(n3301) );
  CLKBUF_X1 U2857 ( .A(n3360), .Z(n3302) );
  CLKBUF_X1 U2858 ( .A(n3360), .Z(n3303) );
  CLKBUF_X1 U2859 ( .A(n3359), .Z(n3304) );
  CLKBUF_X1 U2860 ( .A(n3359), .Z(n3305) );
  CLKBUF_X1 U2861 ( .A(n3359), .Z(n3306) );
  CLKBUF_X1 U2862 ( .A(n3359), .Z(n3307) );
  CLKBUF_X1 U2863 ( .A(n3359), .Z(n3308) );
  CLKBUF_X1 U2864 ( .A(n3359), .Z(n3309) );
  CLKBUF_X1 U2865 ( .A(n3358), .Z(n3310) );
  CLKBUF_X1 U2866 ( .A(n3358), .Z(n3311) );
  CLKBUF_X1 U2867 ( .A(n3358), .Z(n3312) );
  CLKBUF_X1 U2868 ( .A(n3358), .Z(n3313) );
  CLKBUF_X1 U2869 ( .A(n3358), .Z(n3314) );
  CLKBUF_X1 U2870 ( .A(n3358), .Z(n3315) );
  CLKBUF_X1 U2871 ( .A(n3357), .Z(n3316) );
  CLKBUF_X1 U2872 ( .A(n3357), .Z(n3317) );
  CLKBUF_X1 U2873 ( .A(n3357), .Z(n3318) );
  CLKBUF_X1 U2874 ( .A(n3357), .Z(n3319) );
  CLKBUF_X1 U2875 ( .A(n3357), .Z(n3320) );
  CLKBUF_X1 U2876 ( .A(n3357), .Z(n3321) );
  CLKBUF_X1 U2877 ( .A(n3356), .Z(n3322) );
  CLKBUF_X1 U2878 ( .A(n3356), .Z(n3323) );
  CLKBUF_X1 U2879 ( .A(n3356), .Z(n3324) );
  CLKBUF_X1 U2880 ( .A(n3356), .Z(n3325) );
  CLKBUF_X1 U2881 ( .A(n3356), .Z(n3326) );
  CLKBUF_X1 U2882 ( .A(n3356), .Z(n3327) );
  CLKBUF_X1 U2883 ( .A(n3355), .Z(n3328) );
  CLKBUF_X1 U2884 ( .A(n3355), .Z(n3329) );
  CLKBUF_X1 U2885 ( .A(n3355), .Z(n3330) );
  CLKBUF_X1 U2886 ( .A(n3355), .Z(n3331) );
  CLKBUF_X1 U2887 ( .A(n3355), .Z(n3332) );
  CLKBUF_X1 U2888 ( .A(n3355), .Z(n3333) );
  CLKBUF_X1 U2889 ( .A(n3354), .Z(n3334) );
  CLKBUF_X1 U2890 ( .A(n3354), .Z(n3335) );
  CLKBUF_X1 U2891 ( .A(n3354), .Z(n3336) );
  CLKBUF_X1 U2892 ( .A(n3354), .Z(n3337) );
  CLKBUF_X1 U2893 ( .A(n3354), .Z(n3338) );
  CLKBUF_X1 U2894 ( .A(n3354), .Z(n3339) );
  CLKBUF_X1 U2895 ( .A(n3353), .Z(n3340) );
  CLKBUF_X1 U2896 ( .A(n3353), .Z(n3341) );
  CLKBUF_X1 U2897 ( .A(n3353), .Z(n3342) );
  CLKBUF_X1 U2898 ( .A(n3353), .Z(n3343) );
  CLKBUF_X1 U2899 ( .A(n3353), .Z(n3344) );
  CLKBUF_X1 U2900 ( .A(n3353), .Z(n3345) );
  CLKBUF_X1 U2901 ( .A(n3352), .Z(n3346) );
  CLKBUF_X1 U2902 ( .A(n3352), .Z(n3347) );
  CLKBUF_X1 U2903 ( .A(n3352), .Z(n3348) );
  CLKBUF_X1 U2904 ( .A(n3352), .Z(n3349) );
  CLKBUF_X1 U2905 ( .A(n3352), .Z(n3350) );
  CLKBUF_X1 U2906 ( .A(n3352), .Z(n3351) );
  CLKBUF_X3 U2907 ( .A(n1032), .Z(n3352) );
  CLKBUF_X3 U2908 ( .A(n1032), .Z(n3353) );
  CLKBUF_X3 U2909 ( .A(n1033), .Z(n3354) );
  CLKBUF_X3 U2910 ( .A(n1033), .Z(n3355) );
  CLKBUF_X3 U2911 ( .A(n1034), .Z(n3356) );
  CLKBUF_X3 U2912 ( .A(n1034), .Z(n3357) );
  CLKBUF_X3 U2913 ( .A(n1035), .Z(n3358) );
  CLKBUF_X3 U2914 ( .A(n1035), .Z(n3359) );
  CLKBUF_X3 U2915 ( .A(n1036), .Z(n3360) );
  CLKBUF_X3 U2916 ( .A(n1036), .Z(n3361) );
  CLKBUF_X3 U2917 ( .A(n1037), .Z(n3362) );
  CLKBUF_X3 U2918 ( .A(n1037), .Z(n3363) );
  CLKBUF_X3 U2919 ( .A(n1038), .Z(n3364) );
  CLKBUF_X3 U2920 ( .A(n1038), .Z(n3365) );
  CLKBUF_X3 U2921 ( .A(n1039), .Z(n3366) );
  CLKBUF_X3 U2922 ( .A(n1039), .Z(n3367) );
  INV_X2 U2923 ( .A(n1455), .ZN(n3368) );
  INV_X2 U2924 ( .A(n1457), .ZN(n3369) );
  INV_X2 U2925 ( .A(n1458), .ZN(n3370) );
  INV_X2 U2926 ( .A(n1459), .ZN(n3371) );
  INV_X2 U2927 ( .A(n1460), .ZN(n3372) );
  INV_X2 U2928 ( .A(n1461), .ZN(n3373) );
  INV_X2 U2929 ( .A(n1462), .ZN(n3374) );
  INV_X2 U2930 ( .A(n1463), .ZN(n3375) );
  INV_X2 U2931 ( .A(n1464), .ZN(n3376) );
  INV_X2 U2932 ( .A(n1465), .ZN(n3377) );
  INV_X2 U2933 ( .A(n1466), .ZN(n3378) );
  INV_X2 U2934 ( .A(n1467), .ZN(n3379) );
  INV_X2 U2935 ( .A(n1468), .ZN(n3380) );
  INV_X2 U2936 ( .A(n1469), .ZN(n3381) );
  INV_X2 U2937 ( .A(n1470), .ZN(n3382) );
  INV_X2 U2938 ( .A(n1471), .ZN(n3383) );
  INV_X2 U2939 ( .A(n1472), .ZN(n3384) );
  INV_X2 U2940 ( .A(n1473), .ZN(n3385) );
  INV_X2 U2941 ( .A(n1474), .ZN(n3386) );
  INV_X2 U2942 ( .A(n1475), .ZN(n3387) );
  INV_X2 U2943 ( .A(n1476), .ZN(n3388) );
  INV_X2 U2944 ( .A(n1477), .ZN(n3389) );
  INV_X2 U2945 ( .A(n1478), .ZN(n3390) );
  INV_X2 U2946 ( .A(n1479), .ZN(n3391) );
  INV_X2 U2947 ( .A(n1480), .ZN(n3392) );
  INV_X2 U2948 ( .A(n1481), .ZN(n3393) );
  INV_X2 U2949 ( .A(n1482), .ZN(n3394) );
  INV_X2 U2950 ( .A(n1483), .ZN(n3395) );
  INV_X2 U2951 ( .A(n1484), .ZN(n3396) );
  INV_X2 U2952 ( .A(n1485), .ZN(n3397) );
  INV_X2 U2953 ( .A(n1486), .ZN(n3398) );
  INV_X2 U2954 ( .A(n1487), .ZN(n3399) );
  INV_X2 U2955 ( .A(n1422), .ZN(n3400) );
  INV_X2 U2956 ( .A(n1424), .ZN(n3401) );
  INV_X2 U2957 ( .A(n1425), .ZN(n3402) );
  INV_X2 U2958 ( .A(n1426), .ZN(n3403) );
  INV_X2 U2959 ( .A(n1427), .ZN(n3404) );
  INV_X2 U2960 ( .A(n1428), .ZN(n3405) );
  INV_X2 U2961 ( .A(n1429), .ZN(n3406) );
  INV_X2 U2962 ( .A(n1430), .ZN(n3407) );
  INV_X2 U2963 ( .A(n1431), .ZN(n3408) );
  INV_X2 U2964 ( .A(n1432), .ZN(n3409) );
  INV_X2 U2965 ( .A(n1433), .ZN(n3410) );
  INV_X2 U2966 ( .A(n1434), .ZN(n3411) );
  INV_X2 U2967 ( .A(n1435), .ZN(n3412) );
  INV_X2 U2968 ( .A(n1436), .ZN(n3413) );
  INV_X2 U2969 ( .A(n1437), .ZN(n3414) );
  INV_X2 U2970 ( .A(n1438), .ZN(n3415) );
  INV_X2 U2971 ( .A(n1439), .ZN(n3416) );
  INV_X2 U2972 ( .A(n1440), .ZN(n3417) );
  INV_X2 U2973 ( .A(n1441), .ZN(n3418) );
  INV_X2 U2974 ( .A(n1442), .ZN(n3419) );
  INV_X2 U2975 ( .A(n1443), .ZN(n3420) );
  INV_X2 U2976 ( .A(n1444), .ZN(n3421) );
  INV_X2 U2977 ( .A(n1445), .ZN(n3422) );
  INV_X2 U2978 ( .A(n1446), .ZN(n3423) );
  INV_X2 U2979 ( .A(n1447), .ZN(n3424) );
  INV_X2 U2980 ( .A(n1448), .ZN(n3425) );
  INV_X2 U2981 ( .A(n1449), .ZN(n3426) );
  INV_X2 U2982 ( .A(n1450), .ZN(n3427) );
  INV_X2 U2983 ( .A(n1451), .ZN(n3428) );
  INV_X2 U2984 ( .A(n1452), .ZN(n3429) );
  INV_X2 U2985 ( .A(n1453), .ZN(n3430) );
  INV_X2 U2986 ( .A(n1454), .ZN(n3431) );
  INV_X2 U2987 ( .A(n1387), .ZN(n3432) );
  INV_X2 U2988 ( .A(n1389), .ZN(n3433) );
  INV_X2 U2989 ( .A(n1390), .ZN(n3434) );
  INV_X2 U2990 ( .A(n1391), .ZN(n3435) );
  INV_X2 U2991 ( .A(n1392), .ZN(n3436) );
  INV_X2 U2992 ( .A(n1393), .ZN(n3437) );
  INV_X2 U2993 ( .A(n1394), .ZN(n3438) );
  INV_X2 U2994 ( .A(n1395), .ZN(n3439) );
  INV_X2 U2995 ( .A(n1396), .ZN(n3440) );
  INV_X2 U2996 ( .A(n1397), .ZN(n3441) );
  INV_X2 U2997 ( .A(n1398), .ZN(n3442) );
  INV_X2 U2998 ( .A(n1399), .ZN(n3443) );
  INV_X2 U2999 ( .A(n1400), .ZN(n3444) );
  INV_X2 U3000 ( .A(n1401), .ZN(n3445) );
  INV_X2 U3001 ( .A(n1402), .ZN(n3446) );
  INV_X2 U3002 ( .A(n1403), .ZN(n3447) );
  INV_X2 U3003 ( .A(n1404), .ZN(n3448) );
  INV_X2 U3004 ( .A(n1405), .ZN(n3449) );
  INV_X2 U3005 ( .A(n1406), .ZN(n3450) );
  INV_X2 U3006 ( .A(n1407), .ZN(n3451) );
  INV_X2 U3007 ( .A(n1408), .ZN(n3452) );
  INV_X2 U3008 ( .A(n1409), .ZN(n3453) );
  INV_X2 U3009 ( .A(n1410), .ZN(n3454) );
  INV_X2 U3010 ( .A(n1411), .ZN(n3455) );
  INV_X2 U3011 ( .A(n1412), .ZN(n3456) );
  INV_X2 U3012 ( .A(n1413), .ZN(n3457) );
  INV_X2 U3013 ( .A(n1414), .ZN(n3458) );
  INV_X2 U3014 ( .A(n1415), .ZN(n3459) );
  INV_X2 U3015 ( .A(n1416), .ZN(n3460) );
  INV_X2 U3016 ( .A(n1417), .ZN(n3461) );
  INV_X2 U3017 ( .A(n1418), .ZN(n3462) );
  INV_X2 U3018 ( .A(n1419), .ZN(n3463) );
  INV_X2 U3019 ( .A(n1354), .ZN(n3464) );
  INV_X2 U3020 ( .A(n1356), .ZN(n3465) );
  INV_X2 U3021 ( .A(n1357), .ZN(n3466) );
  INV_X2 U3022 ( .A(n1358), .ZN(n3467) );
  INV_X2 U3023 ( .A(n1359), .ZN(n3468) );
  INV_X2 U3024 ( .A(n1360), .ZN(n3469) );
  INV_X2 U3025 ( .A(n1361), .ZN(n3470) );
  INV_X2 U3026 ( .A(n1362), .ZN(n3471) );
  INV_X2 U3027 ( .A(n1363), .ZN(n3472) );
  INV_X2 U3028 ( .A(n1364), .ZN(n3473) );
  INV_X2 U3029 ( .A(n1365), .ZN(n3474) );
  INV_X2 U3030 ( .A(n1366), .ZN(n3475) );
  INV_X2 U3031 ( .A(n1367), .ZN(n3476) );
  INV_X2 U3032 ( .A(n1368), .ZN(n3477) );
  INV_X2 U3033 ( .A(n1369), .ZN(n3478) );
  INV_X2 U3034 ( .A(n1370), .ZN(n3479) );
  INV_X2 U3035 ( .A(n1371), .ZN(n3480) );
  INV_X2 U3036 ( .A(n1372), .ZN(n3481) );
  INV_X2 U3037 ( .A(n1373), .ZN(n3482) );
  INV_X2 U3038 ( .A(n1374), .ZN(n3483) );
  INV_X2 U3039 ( .A(n1375), .ZN(n3484) );
  INV_X2 U3040 ( .A(n1376), .ZN(n3485) );
  INV_X2 U3041 ( .A(n1377), .ZN(n3486) );
  INV_X2 U3042 ( .A(n1378), .ZN(n3487) );
  INV_X2 U3043 ( .A(n1379), .ZN(n3488) );
  INV_X2 U3044 ( .A(n1380), .ZN(n3489) );
  INV_X2 U3045 ( .A(n1381), .ZN(n3490) );
  INV_X2 U3046 ( .A(n1382), .ZN(n3491) );
  INV_X2 U3047 ( .A(n1383), .ZN(n3492) );
  INV_X2 U3048 ( .A(n1384), .ZN(n3493) );
  INV_X2 U3049 ( .A(n1385), .ZN(n3494) );
  INV_X2 U3050 ( .A(n1386), .ZN(n3495) );
  INV_X2 U3051 ( .A(n1559), .ZN(n3496) );
  INV_X2 U3052 ( .A(n1561), .ZN(n3497) );
  INV_X2 U3053 ( .A(n1562), .ZN(n3498) );
  INV_X2 U3054 ( .A(n1563), .ZN(n3499) );
  INV_X2 U3055 ( .A(n1564), .ZN(n3500) );
  INV_X2 U3056 ( .A(n1565), .ZN(n3501) );
  INV_X2 U3057 ( .A(n1566), .ZN(n3502) );
  INV_X2 U3058 ( .A(n1567), .ZN(n3503) );
  INV_X2 U3059 ( .A(n1568), .ZN(n3504) );
  INV_X2 U3060 ( .A(n1569), .ZN(n3505) );
  INV_X2 U3061 ( .A(n1570), .ZN(n3506) );
  INV_X2 U3062 ( .A(n1571), .ZN(n3507) );
  INV_X2 U3063 ( .A(n1572), .ZN(n3508) );
  INV_X2 U3064 ( .A(n1573), .ZN(n3509) );
  INV_X2 U3065 ( .A(n1574), .ZN(n3510) );
  INV_X2 U3066 ( .A(n1575), .ZN(n3511) );
  INV_X2 U3067 ( .A(n1576), .ZN(n3512) );
  INV_X2 U3068 ( .A(n1577), .ZN(n3513) );
  INV_X2 U3069 ( .A(n1578), .ZN(n3514) );
  INV_X2 U3070 ( .A(n1579), .ZN(n3515) );
  INV_X2 U3071 ( .A(n1580), .ZN(n3516) );
  INV_X2 U3072 ( .A(n1581), .ZN(n3517) );
  INV_X2 U3073 ( .A(n1582), .ZN(n3518) );
  INV_X2 U3074 ( .A(n1583), .ZN(n3519) );
  INV_X2 U3075 ( .A(n1584), .ZN(n3520) );
  INV_X2 U3076 ( .A(n1585), .ZN(n3521) );
  INV_X2 U3077 ( .A(n1586), .ZN(n3522) );
  INV_X2 U3078 ( .A(n1587), .ZN(n3523) );
  INV_X2 U3079 ( .A(n1588), .ZN(n3524) );
  INV_X2 U3080 ( .A(n1589), .ZN(n3525) );
  INV_X2 U3081 ( .A(n1590), .ZN(n3526) );
  INV_X2 U3082 ( .A(n1591), .ZN(n3527) );
  INV_X2 U3083 ( .A(n1522), .ZN(n3528) );
  INV_X2 U3084 ( .A(n1524), .ZN(n3529) );
  INV_X2 U3085 ( .A(n1525), .ZN(n3530) );
  INV_X2 U3086 ( .A(n1526), .ZN(n3531) );
  INV_X2 U3087 ( .A(n1527), .ZN(n3532) );
  INV_X2 U3088 ( .A(n1528), .ZN(n3533) );
  INV_X2 U3089 ( .A(n1529), .ZN(n3534) );
  INV_X2 U3090 ( .A(n1530), .ZN(n3535) );
  INV_X2 U3091 ( .A(n1531), .ZN(n3536) );
  INV_X2 U3092 ( .A(n1532), .ZN(n3537) );
  INV_X2 U3093 ( .A(n1533), .ZN(n3538) );
  INV_X2 U3094 ( .A(n1534), .ZN(n3539) );
  INV_X2 U3095 ( .A(n1535), .ZN(n3540) );
  INV_X2 U3096 ( .A(n1536), .ZN(n3541) );
  INV_X2 U3097 ( .A(n1537), .ZN(n3542) );
  INV_X2 U3098 ( .A(n1538), .ZN(n3543) );
  INV_X2 U3099 ( .A(n1539), .ZN(n3544) );
  INV_X2 U3100 ( .A(n1540), .ZN(n3545) );
  INV_X2 U3101 ( .A(n1541), .ZN(n3546) );
  INV_X2 U3102 ( .A(n1542), .ZN(n3547) );
  INV_X2 U3103 ( .A(n1543), .ZN(n3548) );
  INV_X2 U3104 ( .A(n1544), .ZN(n3549) );
  INV_X2 U3105 ( .A(n1545), .ZN(n3550) );
  INV_X2 U3106 ( .A(n1546), .ZN(n3551) );
  INV_X2 U3107 ( .A(n1547), .ZN(n3552) );
  INV_X2 U3108 ( .A(n1548), .ZN(n3553) );
  INV_X2 U3109 ( .A(n1549), .ZN(n3554) );
  INV_X2 U3110 ( .A(n1550), .ZN(n3555) );
  INV_X2 U3111 ( .A(n1551), .ZN(n3556) );
  INV_X2 U3112 ( .A(n1552), .ZN(n3557) );
  INV_X2 U3113 ( .A(n1553), .ZN(n3558) );
  INV_X2 U3114 ( .A(n1554), .ZN(n3559) );
  INV_X2 U3115 ( .A(n1488), .ZN(n3560) );
  INV_X2 U3116 ( .A(n1490), .ZN(n3561) );
  INV_X2 U3117 ( .A(n1491), .ZN(n3562) );
  INV_X2 U3118 ( .A(n1492), .ZN(n3563) );
  INV_X2 U3119 ( .A(n1493), .ZN(n3564) );
  INV_X2 U3120 ( .A(n1494), .ZN(n3565) );
  INV_X2 U3121 ( .A(n1495), .ZN(n3566) );
  INV_X2 U3122 ( .A(n1496), .ZN(n3567) );
  INV_X2 U3123 ( .A(n1497), .ZN(n3568) );
  INV_X2 U3124 ( .A(n1498), .ZN(n3569) );
  INV_X2 U3125 ( .A(n1499), .ZN(n3570) );
  INV_X2 U3126 ( .A(n1500), .ZN(n3571) );
  INV_X2 U3127 ( .A(n1501), .ZN(n3572) );
  INV_X2 U3128 ( .A(n1502), .ZN(n3573) );
  INV_X2 U3129 ( .A(n1503), .ZN(n3574) );
  INV_X2 U3130 ( .A(n1504), .ZN(n3575) );
  INV_X2 U3131 ( .A(n1505), .ZN(n3576) );
  INV_X2 U3132 ( .A(n1506), .ZN(n3577) );
  INV_X2 U3133 ( .A(n1507), .ZN(n3578) );
  INV_X2 U3134 ( .A(n1508), .ZN(n3579) );
  INV_X2 U3135 ( .A(n1509), .ZN(n3580) );
  INV_X2 U3136 ( .A(n1510), .ZN(n3581) );
  INV_X2 U3137 ( .A(n1511), .ZN(n3582) );
  INV_X2 U3138 ( .A(n1512), .ZN(n3583) );
  INV_X2 U3139 ( .A(n1513), .ZN(n3584) );
  INV_X2 U3140 ( .A(n1514), .ZN(n3585) );
  INV_X2 U3141 ( .A(n1515), .ZN(n3586) );
  INV_X2 U3142 ( .A(n1516), .ZN(n3587) );
  INV_X2 U3143 ( .A(n1517), .ZN(n3588) );
  INV_X2 U3144 ( .A(n1518), .ZN(n3589) );
  INV_X2 U3145 ( .A(n1519), .ZN(n3590) );
  INV_X2 U3146 ( .A(n1520), .ZN(n3591) );
  INV_X2 U3147 ( .A(ADD_WR[4]), .ZN(n3592) );
  INV_X2 U3148 ( .A(n1316), .ZN(n3593) );
  INV_X2 U3149 ( .A(n1318), .ZN(n3594) );
  INV_X2 U3150 ( .A(n1319), .ZN(n3595) );
  INV_X2 U3151 ( .A(n1320), .ZN(n3596) );
  INV_X2 U3152 ( .A(n1321), .ZN(n3597) );
  INV_X2 U3153 ( .A(n1322), .ZN(n3598) );
  INV_X2 U3154 ( .A(n1323), .ZN(n3599) );
  INV_X2 U3155 ( .A(n1324), .ZN(n3600) );
  INV_X2 U3156 ( .A(n1325), .ZN(n3601) );
  INV_X2 U3157 ( .A(n1326), .ZN(n3602) );
  INV_X2 U3158 ( .A(n1327), .ZN(n3603) );
  INV_X2 U3159 ( .A(n1328), .ZN(n3604) );
  INV_X2 U3160 ( .A(n1329), .ZN(n3605) );
  INV_X2 U3161 ( .A(n1330), .ZN(n3606) );
  INV_X2 U3162 ( .A(n1331), .ZN(n3607) );
  INV_X2 U3163 ( .A(n1332), .ZN(n3608) );
  INV_X2 U3164 ( .A(n1333), .ZN(n3609) );
  INV_X2 U3165 ( .A(n1334), .ZN(n3610) );
  INV_X2 U3166 ( .A(n1335), .ZN(n3611) );
  INV_X2 U3167 ( .A(n1336), .ZN(n3612) );
  INV_X2 U3168 ( .A(n1337), .ZN(n3613) );
  INV_X2 U3169 ( .A(n1338), .ZN(n3614) );
  INV_X2 U3170 ( .A(n1339), .ZN(n3615) );
  INV_X2 U3171 ( .A(n1340), .ZN(n3616) );
  INV_X2 U3172 ( .A(n1341), .ZN(n3617) );
  INV_X2 U3173 ( .A(n1342), .ZN(n3618) );
  INV_X2 U3174 ( .A(n1343), .ZN(n3619) );
  INV_X2 U3175 ( .A(n1344), .ZN(n3620) );
  INV_X2 U3176 ( .A(n1345), .ZN(n3621) );
  INV_X2 U3177 ( .A(n1346), .ZN(n3622) );
  INV_X2 U3178 ( .A(n1347), .ZN(n3623) );
  INV_X2 U3179 ( .A(n1348), .ZN(n3624) );
  INV_X2 U3180 ( .A(n1283), .ZN(n3625) );
  INV_X2 U3181 ( .A(n1285), .ZN(n3626) );
  INV_X2 U3182 ( .A(n1286), .ZN(n3627) );
  INV_X2 U3183 ( .A(n1287), .ZN(n3628) );
  INV_X2 U3184 ( .A(n1288), .ZN(n3629) );
  INV_X2 U3185 ( .A(n1289), .ZN(n3630) );
  INV_X2 U3186 ( .A(n1290), .ZN(n3631) );
  INV_X2 U3187 ( .A(n1291), .ZN(n3632) );
  INV_X2 U3188 ( .A(n1292), .ZN(n3633) );
  INV_X2 U3189 ( .A(n1293), .ZN(n3634) );
  INV_X2 U3190 ( .A(n1294), .ZN(n3635) );
  INV_X2 U3191 ( .A(n1295), .ZN(n3636) );
  INV_X2 U3192 ( .A(n1296), .ZN(n3637) );
  INV_X2 U3193 ( .A(n1297), .ZN(n3638) );
  INV_X2 U3194 ( .A(n1298), .ZN(n3639) );
  INV_X2 U3195 ( .A(n1299), .ZN(n3640) );
  INV_X2 U3196 ( .A(n1300), .ZN(n3641) );
  INV_X2 U3197 ( .A(n1301), .ZN(n3642) );
  INV_X2 U3198 ( .A(n1302), .ZN(n3643) );
  INV_X2 U3199 ( .A(n1303), .ZN(n3644) );
  INV_X2 U3200 ( .A(n1304), .ZN(n3645) );
  INV_X2 U3201 ( .A(n1305), .ZN(n3646) );
  INV_X2 U3202 ( .A(n1306), .ZN(n3647) );
  INV_X2 U3203 ( .A(n1307), .ZN(n3648) );
  INV_X2 U3204 ( .A(n1308), .ZN(n3649) );
  INV_X2 U3205 ( .A(n1309), .ZN(n3650) );
  INV_X2 U3206 ( .A(n1310), .ZN(n3651) );
  INV_X2 U3207 ( .A(n1311), .ZN(n3652) );
  INV_X2 U3208 ( .A(n1312), .ZN(n3653) );
  INV_X2 U3209 ( .A(n1313), .ZN(n3654) );
  INV_X2 U3210 ( .A(n1314), .ZN(n3655) );
  INV_X2 U3211 ( .A(n1315), .ZN(n3656) );
  INV_X2 U3212 ( .A(n1248), .ZN(n3657) );
  INV_X2 U3213 ( .A(n1250), .ZN(n3658) );
  INV_X2 U3214 ( .A(n1251), .ZN(n3659) );
  INV_X2 U3215 ( .A(n1252), .ZN(n3660) );
  INV_X2 U3216 ( .A(n1253), .ZN(n3661) );
  INV_X2 U3217 ( .A(n1254), .ZN(n3662) );
  INV_X2 U3218 ( .A(n1255), .ZN(n3663) );
  INV_X2 U3219 ( .A(n1256), .ZN(n3664) );
  INV_X2 U3220 ( .A(n1257), .ZN(n3665) );
  INV_X2 U3221 ( .A(n1258), .ZN(n3666) );
  INV_X2 U3222 ( .A(n1259), .ZN(n3667) );
  INV_X2 U3223 ( .A(n1260), .ZN(n3668) );
  INV_X2 U3224 ( .A(n1261), .ZN(n3669) );
  INV_X2 U3225 ( .A(n1262), .ZN(n3670) );
  INV_X2 U3226 ( .A(n1263), .ZN(n3671) );
  INV_X2 U3227 ( .A(n1264), .ZN(n3672) );
  INV_X2 U3228 ( .A(n1265), .ZN(n3673) );
  INV_X2 U3229 ( .A(n1266), .ZN(n3674) );
  INV_X2 U3230 ( .A(n1267), .ZN(n3675) );
  INV_X2 U3231 ( .A(n1268), .ZN(n3676) );
  INV_X2 U3232 ( .A(n1269), .ZN(n3677) );
  INV_X2 U3233 ( .A(n1270), .ZN(n3678) );
  INV_X2 U3234 ( .A(n1271), .ZN(n3679) );
  INV_X2 U3235 ( .A(n1272), .ZN(n3680) );
  INV_X2 U3236 ( .A(n1273), .ZN(n3681) );
  INV_X2 U3237 ( .A(n1274), .ZN(n3682) );
  INV_X2 U3238 ( .A(n1275), .ZN(n3683) );
  INV_X2 U3239 ( .A(n1276), .ZN(n3684) );
  INV_X2 U3240 ( .A(n1277), .ZN(n3685) );
  INV_X2 U3241 ( .A(n1278), .ZN(n3686) );
  INV_X2 U3242 ( .A(n1279), .ZN(n3687) );
  INV_X2 U3243 ( .A(n1280), .ZN(n3688) );
  INV_X2 U3244 ( .A(n1214), .ZN(n3689) );
  INV_X2 U3245 ( .A(n1216), .ZN(n3690) );
  INV_X2 U3246 ( .A(n1217), .ZN(n3691) );
  INV_X2 U3247 ( .A(n1218), .ZN(n3692) );
  INV_X2 U3248 ( .A(n1219), .ZN(n3693) );
  INV_X2 U3249 ( .A(n1220), .ZN(n3694) );
  INV_X2 U3250 ( .A(n1221), .ZN(n3695) );
  INV_X2 U3251 ( .A(n1222), .ZN(n3696) );
  INV_X2 U3252 ( .A(n1223), .ZN(n3697) );
  INV_X2 U3253 ( .A(n1224), .ZN(n3698) );
  INV_X2 U3254 ( .A(n1225), .ZN(n3699) );
  INV_X2 U3255 ( .A(n1226), .ZN(n3700) );
  INV_X2 U3256 ( .A(n1227), .ZN(n3701) );
  INV_X2 U3257 ( .A(n1228), .ZN(n3702) );
  INV_X2 U3258 ( .A(n1229), .ZN(n3703) );
  INV_X2 U3259 ( .A(n1230), .ZN(n3704) );
  INV_X2 U3260 ( .A(n1231), .ZN(n3705) );
  INV_X2 U3261 ( .A(n1232), .ZN(n3706) );
  INV_X2 U3262 ( .A(n1233), .ZN(n3707) );
  INV_X2 U3263 ( .A(n1234), .ZN(n3708) );
  INV_X2 U3264 ( .A(n1235), .ZN(n3709) );
  INV_X2 U3265 ( .A(n1236), .ZN(n3710) );
  INV_X2 U3266 ( .A(n1237), .ZN(n3711) );
  INV_X2 U3267 ( .A(n1238), .ZN(n3712) );
  INV_X2 U3268 ( .A(n1239), .ZN(n3713) );
  INV_X2 U3269 ( .A(n1240), .ZN(n3714) );
  INV_X2 U3270 ( .A(n1241), .ZN(n3715) );
  INV_X2 U3271 ( .A(n1242), .ZN(n3716) );
  INV_X2 U3272 ( .A(n1243), .ZN(n3717) );
  INV_X2 U3273 ( .A(n1244), .ZN(n3718) );
  INV_X2 U3274 ( .A(n1245), .ZN(n3719) );
  INV_X2 U3275 ( .A(n1246), .ZN(n3720) );
  INV_X2 U3276 ( .A(n1179), .ZN(n3721) );
  INV_X2 U3277 ( .A(n1181), .ZN(n3722) );
  INV_X2 U3278 ( .A(n1182), .ZN(n3723) );
  INV_X2 U3279 ( .A(n1183), .ZN(n3724) );
  INV_X2 U3280 ( .A(n1184), .ZN(n3725) );
  INV_X2 U3281 ( .A(n1185), .ZN(n3726) );
  INV_X2 U3282 ( .A(n1186), .ZN(n3727) );
  INV_X2 U3283 ( .A(n1187), .ZN(n3728) );
  INV_X2 U3284 ( .A(n1188), .ZN(n3729) );
  INV_X2 U3285 ( .A(n1189), .ZN(n3730) );
  INV_X2 U3286 ( .A(n1190), .ZN(n3731) );
  INV_X2 U3287 ( .A(n1191), .ZN(n3732) );
  INV_X2 U3288 ( .A(n1192), .ZN(n3733) );
  INV_X2 U3289 ( .A(n1193), .ZN(n3734) );
  INV_X2 U3290 ( .A(n1194), .ZN(n3735) );
  INV_X2 U3291 ( .A(n1195), .ZN(n3736) );
  INV_X2 U3292 ( .A(n1196), .ZN(n3737) );
  INV_X2 U3293 ( .A(n1197), .ZN(n3738) );
  INV_X2 U3294 ( .A(n1198), .ZN(n3739) );
  INV_X2 U3295 ( .A(n1199), .ZN(n3740) );
  INV_X2 U3296 ( .A(n1200), .ZN(n3741) );
  INV_X2 U3297 ( .A(n1201), .ZN(n3742) );
  INV_X2 U3298 ( .A(n1202), .ZN(n3743) );
  INV_X2 U3299 ( .A(n1203), .ZN(n3744) );
  INV_X2 U3300 ( .A(n1204), .ZN(n3745) );
  INV_X2 U3301 ( .A(n1205), .ZN(n3746) );
  INV_X2 U3302 ( .A(n1206), .ZN(n3747) );
  INV_X2 U3303 ( .A(n1207), .ZN(n3748) );
  INV_X2 U3304 ( .A(n1208), .ZN(n3749) );
  INV_X2 U3305 ( .A(n1209), .ZN(n3750) );
  INV_X2 U3306 ( .A(n1210), .ZN(n3751) );
  INV_X2 U3307 ( .A(n1211), .ZN(n3752) );
  INV_X2 U3308 ( .A(n1145), .ZN(n3753) );
  INV_X2 U3309 ( .A(n1147), .ZN(n3754) );
  INV_X2 U3310 ( .A(n1148), .ZN(n3755) );
  INV_X2 U3311 ( .A(n1149), .ZN(n3756) );
  INV_X2 U3312 ( .A(n1150), .ZN(n3757) );
  INV_X2 U3313 ( .A(n1151), .ZN(n3758) );
  INV_X2 U3314 ( .A(n1152), .ZN(n3759) );
  INV_X2 U3315 ( .A(n1153), .ZN(n3760) );
  INV_X2 U3316 ( .A(n1154), .ZN(n3761) );
  INV_X2 U3317 ( .A(n1155), .ZN(n3762) );
  INV_X2 U3318 ( .A(n1156), .ZN(n3763) );
  INV_X2 U3319 ( .A(n1157), .ZN(n3764) );
  INV_X2 U3320 ( .A(n1158), .ZN(n3765) );
  INV_X2 U3321 ( .A(n1159), .ZN(n3766) );
  INV_X2 U3322 ( .A(n1160), .ZN(n3767) );
  INV_X2 U3323 ( .A(n1161), .ZN(n3768) );
  INV_X2 U3324 ( .A(n1162), .ZN(n3769) );
  INV_X2 U3325 ( .A(n1163), .ZN(n3770) );
  INV_X2 U3326 ( .A(n1164), .ZN(n3771) );
  INV_X2 U3327 ( .A(n1165), .ZN(n3772) );
  INV_X2 U3328 ( .A(n1166), .ZN(n3773) );
  INV_X2 U3329 ( .A(n1167), .ZN(n3774) );
  INV_X2 U3330 ( .A(n1168), .ZN(n3775) );
  INV_X2 U3331 ( .A(n1169), .ZN(n3776) );
  INV_X2 U3332 ( .A(n1170), .ZN(n3777) );
  INV_X2 U3333 ( .A(n1171), .ZN(n3778) );
  INV_X2 U3334 ( .A(n1172), .ZN(n3779) );
  INV_X2 U3335 ( .A(n1173), .ZN(n3780) );
  INV_X2 U3336 ( .A(n1174), .ZN(n3781) );
  INV_X2 U3337 ( .A(n1175), .ZN(n3782) );
  INV_X2 U3338 ( .A(n1176), .ZN(n3783) );
  INV_X2 U3339 ( .A(n1177), .ZN(n3784) );
  INV_X2 U3340 ( .A(n1107), .ZN(n3785) );
  INV_X2 U3341 ( .A(n1109), .ZN(n3786) );
  INV_X2 U3342 ( .A(n1110), .ZN(n3787) );
  INV_X2 U3343 ( .A(n1111), .ZN(n3788) );
  INV_X2 U3344 ( .A(n1112), .ZN(n3789) );
  INV_X2 U3345 ( .A(n1113), .ZN(n3790) );
  INV_X2 U3346 ( .A(n1114), .ZN(n3791) );
  INV_X2 U3347 ( .A(n1115), .ZN(n3792) );
  INV_X2 U3348 ( .A(n1116), .ZN(n3793) );
  INV_X2 U3349 ( .A(n1117), .ZN(n3794) );
  INV_X2 U3350 ( .A(n1118), .ZN(n3795) );
  INV_X2 U3351 ( .A(n1119), .ZN(n3796) );
  INV_X2 U3352 ( .A(n1120), .ZN(n3797) );
  INV_X2 U3353 ( .A(n1121), .ZN(n3798) );
  INV_X2 U3354 ( .A(n1122), .ZN(n3799) );
  INV_X2 U3355 ( .A(n1123), .ZN(n3800) );
  INV_X2 U3356 ( .A(n1124), .ZN(n3801) );
  INV_X2 U3357 ( .A(n1125), .ZN(n3802) );
  INV_X2 U3358 ( .A(n1126), .ZN(n3803) );
  INV_X2 U3359 ( .A(n1127), .ZN(n3804) );
  INV_X2 U3360 ( .A(n1128), .ZN(n3805) );
  INV_X2 U3361 ( .A(n1129), .ZN(n3806) );
  INV_X2 U3362 ( .A(n1130), .ZN(n3807) );
  INV_X2 U3363 ( .A(n1131), .ZN(n3808) );
  INV_X2 U3364 ( .A(n1132), .ZN(n3809) );
  INV_X2 U3365 ( .A(n1133), .ZN(n3810) );
  INV_X2 U3366 ( .A(n1134), .ZN(n3811) );
  INV_X2 U3367 ( .A(n1135), .ZN(n3812) );
  INV_X2 U3368 ( .A(n1136), .ZN(n3813) );
  INV_X2 U3369 ( .A(n1137), .ZN(n3814) );
  INV_X2 U3370 ( .A(n1138), .ZN(n3815) );
  INV_X2 U3371 ( .A(n1139), .ZN(n3816) );
  INV_X2 U3372 ( .A(n1073), .ZN(n3817) );
  INV_X2 U3373 ( .A(n1075), .ZN(n3818) );
  INV_X2 U3374 ( .A(n1076), .ZN(n3819) );
  INV_X2 U3375 ( .A(n1077), .ZN(n3820) );
  INV_X2 U3376 ( .A(n1078), .ZN(n3821) );
  INV_X2 U3377 ( .A(n1079), .ZN(n3822) );
  INV_X2 U3378 ( .A(n1080), .ZN(n3823) );
  INV_X2 U3379 ( .A(n1081), .ZN(n3824) );
  INV_X2 U3380 ( .A(n1082), .ZN(n3825) );
  INV_X2 U3381 ( .A(n1083), .ZN(n3826) );
  INV_X2 U3382 ( .A(n1084), .ZN(n3827) );
  INV_X2 U3383 ( .A(n1085), .ZN(n3828) );
  INV_X2 U3384 ( .A(n1086), .ZN(n3829) );
  INV_X2 U3385 ( .A(n1087), .ZN(n3830) );
  INV_X2 U3386 ( .A(n1088), .ZN(n3831) );
  INV_X2 U3387 ( .A(n1089), .ZN(n3832) );
  INV_X2 U3388 ( .A(n1090), .ZN(n3833) );
  INV_X2 U3389 ( .A(n1091), .ZN(n3834) );
  INV_X2 U3390 ( .A(n1092), .ZN(n3835) );
  INV_X2 U3391 ( .A(n1093), .ZN(n3836) );
  INV_X2 U3392 ( .A(n1094), .ZN(n3837) );
  INV_X2 U3393 ( .A(n1095), .ZN(n3838) );
  INV_X2 U3394 ( .A(n1096), .ZN(n3839) );
  INV_X2 U3395 ( .A(n1097), .ZN(n3840) );
  INV_X2 U3396 ( .A(n1098), .ZN(n3841) );
  INV_X2 U3397 ( .A(n1099), .ZN(n3842) );
  INV_X2 U3398 ( .A(n1100), .ZN(n3843) );
  INV_X2 U3399 ( .A(n1101), .ZN(n3844) );
  INV_X2 U3400 ( .A(n1102), .ZN(n3845) );
  INV_X2 U3401 ( .A(n1103), .ZN(n3846) );
  INV_X2 U3402 ( .A(n1104), .ZN(n3847) );
  INV_X2 U3403 ( .A(n1105), .ZN(n3848) );
  INV_X2 U3404 ( .A(ADD_WR[3]), .ZN(n3849) );
  INV_X2 U3405 ( .A(ADD_WR[2]), .ZN(n3850) );
  INV_X2 U3406 ( .A(ADD_WR[1]), .ZN(n3851) );
  INV_X2 U3407 ( .A(ADD_WR[0]), .ZN(n3852) );
  INV_X2 U3408 ( .A(ADD_RD1[3]), .ZN(n3853) );
  INV_X2 U3409 ( .A(ADD_RD1[1]), .ZN(n3854) );
  INV_X2 U3410 ( .A(ADD_RD1[0]), .ZN(n3855) );
  INV_X2 U3411 ( .A(ADD_RD2[3]), .ZN(n3856) );
  INV_X2 U3412 ( .A(ADD_RD2[1]), .ZN(n3857) );
  INV_X2 U3413 ( .A(ADD_RD2[0]), .ZN(n3858) );
  INV_X2 U3414 ( .A(DATAIN[31]), .ZN(n3859) );
  INV_X2 U3415 ( .A(DATAIN[30]), .ZN(n3860) );
  INV_X2 U3416 ( .A(DATAIN[29]), .ZN(n3861) );
  INV_X2 U3417 ( .A(DATAIN[28]), .ZN(n3862) );
  INV_X2 U3418 ( .A(DATAIN[27]), .ZN(n3863) );
  INV_X2 U3419 ( .A(DATAIN[26]), .ZN(n3864) );
  INV_X2 U3420 ( .A(DATAIN[25]), .ZN(n3865) );
  INV_X2 U3421 ( .A(DATAIN[24]), .ZN(n3866) );
  INV_X2 U3422 ( .A(DATAIN[23]), .ZN(n3867) );
  INV_X2 U3423 ( .A(DATAIN[22]), .ZN(n3868) );
  INV_X2 U3424 ( .A(DATAIN[21]), .ZN(n3869) );
  INV_X2 U3425 ( .A(DATAIN[20]), .ZN(n3870) );
  INV_X2 U3426 ( .A(DATAIN[19]), .ZN(n3871) );
  INV_X2 U3427 ( .A(DATAIN[18]), .ZN(n3872) );
  INV_X2 U3428 ( .A(DATAIN[17]), .ZN(n3873) );
  INV_X2 U3429 ( .A(DATAIN[16]), .ZN(n3874) );
  INV_X2 U3430 ( .A(DATAIN[15]), .ZN(n3875) );
  INV_X2 U3431 ( .A(DATAIN[14]), .ZN(n3876) );
  INV_X2 U3432 ( .A(DATAIN[13]), .ZN(n3877) );
  INV_X2 U3433 ( .A(DATAIN[12]), .ZN(n3878) );
  INV_X2 U3434 ( .A(DATAIN[11]), .ZN(n3879) );
  INV_X2 U3435 ( .A(DATAIN[10]), .ZN(n3880) );
  INV_X2 U3436 ( .A(DATAIN[9]), .ZN(n3881) );
  INV_X2 U3437 ( .A(DATAIN[8]), .ZN(n3882) );
  INV_X2 U3438 ( .A(DATAIN[7]), .ZN(n3883) );
  INV_X2 U3439 ( .A(DATAIN[6]), .ZN(n3884) );
  INV_X2 U3440 ( .A(DATAIN[5]), .ZN(n3885) );
  INV_X2 U3441 ( .A(DATAIN[4]), .ZN(n3886) );
  INV_X2 U3442 ( .A(DATAIN[3]), .ZN(n3887) );
  INV_X2 U3443 ( .A(DATAIN[2]), .ZN(n3888) );
  INV_X2 U3444 ( .A(DATAIN[1]), .ZN(n3889) );
  INV_X2 U3445 ( .A(DATAIN[0]), .ZN(n3890) );
  INV_X2 U3446 ( .A(CLK), .ZN(n3891) );
endmodule


module REG_PIPO_6_00_00_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n4, n5, n6, n7, n8, n3, n9, n10, n11, n12, n13, n14;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  AOI22_X2 U3 ( .A1(DIN[0]), .A2(n2), .B1(n14), .B2(DOUT[0]), .ZN(n1) );
  AOI22_X2 U5 ( .A1(DIN[1]), .A2(n2), .B1(n14), .B2(DOUT[1]), .ZN(n4) );
  AOI22_X2 U7 ( .A1(DIN[2]), .A2(n2), .B1(n14), .B2(DOUT[2]), .ZN(n5) );
  AOI22_X2 U9 ( .A1(DIN[3]), .A2(n2), .B1(n14), .B2(DOUT[3]), .ZN(n6) );
  AOI22_X2 U11 ( .A1(DIN[4]), .A2(n2), .B1(n14), .B2(DOUT[4]), .ZN(n7) );
  AOI22_X2 U13 ( .A1(DIN[5]), .A2(n2), .B1(n14), .B2(DOUT[5]), .ZN(n8) );
  NOR2_X2 U14 ( .A1(INIT), .A2(n14), .ZN(n2) );
  INV_X2 U2 ( .A(n8), .ZN(n3) );
  INV_X2 U4 ( .A(n7), .ZN(n9) );
  INV_X2 U6 ( .A(n6), .ZN(n10) );
  INV_X2 U8 ( .A(n5), .ZN(n11) );
  INV_X2 U10 ( .A(n4), .ZN(n12) );
  INV_X2 U12 ( .A(n1), .ZN(n13) );
  INV_X2 U15 ( .A(EN), .ZN(n14) );
endmodule


module REG_PIPO_32_00000000_00000000_10 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_9 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_8 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_7 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n9), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n10), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n11), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n13), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n14), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n15), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[25]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[26]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[27]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[29]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[30]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[31]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_5_00_00_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n4, n5, n6, n7, n3, n8, n9, n10, n11, n12;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  AOI22_X2 U3 ( .A1(DIN[0]), .A2(n2), .B1(n12), .B2(DOUT[0]), .ZN(n1) );
  AOI22_X2 U5 ( .A1(DIN[1]), .A2(n2), .B1(n12), .B2(DOUT[1]), .ZN(n4) );
  AOI22_X2 U7 ( .A1(DIN[2]), .A2(n2), .B1(n12), .B2(DOUT[2]), .ZN(n5) );
  AOI22_X2 U9 ( .A1(DIN[3]), .A2(n2), .B1(n12), .B2(DOUT[3]), .ZN(n6) );
  AOI22_X2 U11 ( .A1(DIN[4]), .A2(n2), .B1(n12), .B2(DOUT[4]), .ZN(n7) );
  NOR2_X2 U12 ( .A1(INIT), .A2(n12), .ZN(n2) );
  INV_X2 U2 ( .A(n7), .ZN(n3) );
  INV_X2 U4 ( .A(n6), .ZN(n8) );
  INV_X2 U6 ( .A(n5), .ZN(n9) );
  INV_X2 U8 ( .A(n4), .ZN(n10) );
  INV_X2 U10 ( .A(n1), .ZN(n11) );
  INV_X2 U13 ( .A(EN), .ZN(n12) );
endmodule


module REG_PIPO_5_00_00_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  AOI22_X2 U3 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  AOI22_X2 U5 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  AOI22_X2 U7 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  AOI22_X2 U9 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  AOI22_X2 U11 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  NOR2_X2 U12 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X2 U2 ( .A(n13), .ZN(n3) );
  INV_X2 U4 ( .A(n14), .ZN(n8) );
  INV_X2 U6 ( .A(n15), .ZN(n9) );
  INV_X2 U8 ( .A(n16), .ZN(n10) );
  INV_X2 U10 ( .A(n18), .ZN(n11) );
  INV_X2 U13 ( .A(EN), .ZN(n12) );
endmodule


module ALU_DATA_W32_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189;

  INV_X2 U1 ( .A(n142), .ZN(GE) );
  INV_X2 U2 ( .A(n52), .ZN(n2) );
  INV_X2 U3 ( .A(n143), .ZN(n3) );
  INV_X2 U4 ( .A(B[29]), .ZN(n4) );
  INV_X2 U5 ( .A(n63), .ZN(n5) );
  INV_X2 U6 ( .A(B[28]), .ZN(n6) );
  INV_X2 U7 ( .A(n64), .ZN(n7) );
  INV_X2 U8 ( .A(B[27]), .ZN(n8) );
  INV_X2 U9 ( .A(B[26]), .ZN(n9) );
  INV_X2 U10 ( .A(B[25]), .ZN(n10) );
  INV_X2 U11 ( .A(n73), .ZN(n11) );
  INV_X2 U12 ( .A(B[24]), .ZN(n12) );
  INV_X2 U13 ( .A(n74), .ZN(n13) );
  INV_X2 U14 ( .A(B[23]), .ZN(n14) );
  INV_X2 U15 ( .A(B[22]), .ZN(n15) );
  INV_X2 U16 ( .A(B[21]), .ZN(n16) );
  INV_X2 U17 ( .A(n83), .ZN(n17) );
  INV_X2 U18 ( .A(B[20]), .ZN(n18) );
  INV_X2 U19 ( .A(n84), .ZN(n19) );
  INV_X2 U20 ( .A(B[19]), .ZN(n20) );
  INV_X2 U21 ( .A(B[18]), .ZN(n21) );
  INV_X2 U22 ( .A(B[17]), .ZN(n22) );
  INV_X2 U23 ( .A(n93), .ZN(n23) );
  INV_X2 U24 ( .A(B[16]), .ZN(n24) );
  INV_X2 U25 ( .A(n94), .ZN(n25) );
  INV_X2 U26 ( .A(B[15]), .ZN(n26) );
  INV_X2 U27 ( .A(B[14]), .ZN(n27) );
  INV_X2 U28 ( .A(B[13]), .ZN(n28) );
  INV_X2 U29 ( .A(n103), .ZN(n29) );
  INV_X2 U30 ( .A(B[12]), .ZN(n30) );
  INV_X2 U31 ( .A(n104), .ZN(n31) );
  INV_X2 U32 ( .A(B[11]), .ZN(n32) );
  INV_X2 U33 ( .A(B[10]), .ZN(n33) );
  INV_X2 U34 ( .A(B[9]), .ZN(n34) );
  INV_X2 U35 ( .A(n113), .ZN(n35) );
  INV_X2 U36 ( .A(B[8]), .ZN(n36) );
  INV_X2 U37 ( .A(n114), .ZN(n37) );
  INV_X2 U38 ( .A(B[7]), .ZN(n38) );
  INV_X2 U39 ( .A(B[6]), .ZN(n39) );
  INV_X2 U40 ( .A(B[5]), .ZN(n40) );
  INV_X2 U41 ( .A(n123), .ZN(n41) );
  INV_X2 U42 ( .A(B[4]), .ZN(n42) );
  INV_X2 U43 ( .A(n124), .ZN(n43) );
  INV_X2 U44 ( .A(B[3]), .ZN(n44) );
  INV_X2 U45 ( .A(B[2]), .ZN(n45) );
  INV_X2 U46 ( .A(n189), .ZN(n46) );
  INV_X2 U47 ( .A(n127), .ZN(n47) );
  INV_X2 U48 ( .A(B[0]), .ZN(n48) );
  INV_X2 U49 ( .A(A[31]), .ZN(n49) );
  INV_X2 U50 ( .A(A[30]), .ZN(n50) );
  INV_X2 U51 ( .A(A[1]), .ZN(n51) );
  NAND2_X1 U52 ( .A1(GE), .A2(LE), .ZN(NE) );
  AOI21_X1 U53 ( .B1(n52), .B2(A[31]), .A(n53), .ZN(LE) );
  AOI21_X1 U54 ( .B1(n49), .B2(n2), .A(B[31]), .ZN(n53) );
  OAI21_X1 U55 ( .B1(B[30]), .B2(n50), .A(n54), .ZN(n52) );
  OAI211_X1 U56 ( .C1(n55), .C2(n56), .A(n57), .B(n58), .ZN(n54) );
  NAND2_X1 U57 ( .A1(n59), .A2(n60), .ZN(n56) );
  AOI211_X1 U58 ( .C1(n61), .C2(n62), .A(n63), .B(n64), .ZN(n55) );
  OAI211_X1 U59 ( .C1(n65), .C2(n66), .A(n67), .B(n68), .ZN(n62) );
  NAND2_X1 U60 ( .A1(n69), .A2(n70), .ZN(n66) );
  AOI211_X1 U61 ( .C1(n71), .C2(n72), .A(n73), .B(n74), .ZN(n65) );
  OAI211_X1 U62 ( .C1(n75), .C2(n76), .A(n77), .B(n78), .ZN(n72) );
  NAND2_X1 U63 ( .A1(n79), .A2(n80), .ZN(n76) );
  AOI211_X1 U64 ( .C1(n81), .C2(n82), .A(n83), .B(n84), .ZN(n75) );
  OAI211_X1 U65 ( .C1(n85), .C2(n86), .A(n87), .B(n88), .ZN(n82) );
  NAND2_X1 U66 ( .A1(n89), .A2(n90), .ZN(n86) );
  AOI211_X1 U67 ( .C1(n91), .C2(n92), .A(n93), .B(n94), .ZN(n85) );
  OAI211_X1 U68 ( .C1(n95), .C2(n96), .A(n97), .B(n98), .ZN(n92) );
  NAND2_X1 U69 ( .A1(n99), .A2(n100), .ZN(n96) );
  AOI211_X1 U70 ( .C1(n101), .C2(n102), .A(n103), .B(n104), .ZN(n95) );
  OAI211_X1 U71 ( .C1(n105), .C2(n106), .A(n107), .B(n108), .ZN(n102) );
  NAND2_X1 U72 ( .A1(n109), .A2(n110), .ZN(n106) );
  AOI211_X1 U73 ( .C1(n111), .C2(n112), .A(n113), .B(n114), .ZN(n105) );
  OAI211_X1 U74 ( .C1(n115), .C2(n116), .A(n117), .B(n118), .ZN(n112) );
  NAND2_X1 U75 ( .A1(n119), .A2(n120), .ZN(n116) );
  AOI211_X1 U76 ( .C1(n121), .C2(n122), .A(n123), .B(n124), .ZN(n115) );
  OAI211_X1 U77 ( .C1(A[1]), .C2(n47), .A(n125), .B(n126), .ZN(n122) );
  OAI21_X1 U78 ( .B1(n51), .B2(n127), .A(B[1]), .ZN(n125) );
  NAND2_X1 U79 ( .A1(A[0]), .A2(n48), .ZN(n127) );
  AND2_X1 U80 ( .A1(n128), .A2(n129), .ZN(n121) );
  AND2_X1 U81 ( .A1(n130), .A2(n131), .ZN(n111) );
  AND2_X1 U82 ( .A1(n132), .A2(n133), .ZN(n101) );
  AND2_X1 U83 ( .A1(n134), .A2(n135), .ZN(n91) );
  AND2_X1 U84 ( .A1(n136), .A2(n137), .ZN(n81) );
  AND2_X1 U85 ( .A1(n138), .A2(n139), .ZN(n71) );
  AND2_X1 U86 ( .A1(n140), .A2(n141), .ZN(n61) );
  OAI21_X1 U87 ( .B1(A[31]), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U88 ( .B1(n3), .B2(n49), .A(B[31]), .ZN(n144) );
  AOI21_X1 U89 ( .B1(n50), .B2(B[30]), .A(n145), .ZN(n143) );
  AND3_X1 U90 ( .A1(n146), .A2(n59), .A3(n58), .ZN(n145) );
  XOR2_X1 U91 ( .A(n50), .B(B[30]), .Z(n58) );
  NAND2_X1 U92 ( .A1(A[29]), .A2(n4), .ZN(n59) );
  NAND3_X1 U93 ( .A1(n147), .A2(n148), .A3(n57), .ZN(n146) );
  OR2_X1 U94 ( .A1(n4), .A2(A[29]), .ZN(n57) );
  NAND3_X1 U95 ( .A1(n149), .A2(n141), .A3(n5), .ZN(n147) );
  NAND2_X1 U96 ( .A1(n148), .A2(n60), .ZN(n63) );
  NAND2_X1 U97 ( .A1(A[28]), .A2(n6), .ZN(n60) );
  OR2_X1 U98 ( .A1(n6), .A2(A[28]), .ZN(n148) );
  NAND2_X1 U99 ( .A1(A[27]), .A2(n8), .ZN(n141) );
  NAND3_X1 U100 ( .A1(n150), .A2(n151), .A3(n7), .ZN(n149) );
  NOR2_X1 U101 ( .A1(n8), .A2(A[27]), .ZN(n64) );
  NAND3_X1 U102 ( .A1(n152), .A2(n69), .A3(n68), .ZN(n150) );
  AND2_X1 U103 ( .A1(n151), .A2(n140), .ZN(n68) );
  NAND2_X1 U104 ( .A1(A[26]), .A2(n9), .ZN(n140) );
  OR2_X1 U105 ( .A1(n9), .A2(A[26]), .ZN(n151) );
  NAND2_X1 U106 ( .A1(A[25]), .A2(n10), .ZN(n69) );
  NAND3_X1 U107 ( .A1(n153), .A2(n154), .A3(n67), .ZN(n152) );
  OR2_X1 U108 ( .A1(n10), .A2(A[25]), .ZN(n67) );
  NAND3_X1 U109 ( .A1(n155), .A2(n139), .A3(n11), .ZN(n153) );
  NAND2_X1 U110 ( .A1(n154), .A2(n70), .ZN(n73) );
  NAND2_X1 U111 ( .A1(A[24]), .A2(n12), .ZN(n70) );
  OR2_X1 U112 ( .A1(n12), .A2(A[24]), .ZN(n154) );
  NAND2_X1 U113 ( .A1(A[23]), .A2(n14), .ZN(n139) );
  NAND3_X1 U114 ( .A1(n156), .A2(n157), .A3(n13), .ZN(n155) );
  NOR2_X1 U115 ( .A1(n14), .A2(A[23]), .ZN(n74) );
  NAND3_X1 U116 ( .A1(n158), .A2(n79), .A3(n78), .ZN(n156) );
  AND2_X1 U117 ( .A1(n157), .A2(n138), .ZN(n78) );
  NAND2_X1 U118 ( .A1(A[22]), .A2(n15), .ZN(n138) );
  OR2_X1 U119 ( .A1(n15), .A2(A[22]), .ZN(n157) );
  NAND2_X1 U120 ( .A1(A[21]), .A2(n16), .ZN(n79) );
  NAND3_X1 U121 ( .A1(n159), .A2(n160), .A3(n77), .ZN(n158) );
  OR2_X1 U122 ( .A1(n16), .A2(A[21]), .ZN(n77) );
  NAND3_X1 U123 ( .A1(n161), .A2(n137), .A3(n17), .ZN(n159) );
  NAND2_X1 U124 ( .A1(n160), .A2(n80), .ZN(n83) );
  NAND2_X1 U125 ( .A1(A[20]), .A2(n18), .ZN(n80) );
  OR2_X1 U126 ( .A1(n18), .A2(A[20]), .ZN(n160) );
  NAND2_X1 U127 ( .A1(A[19]), .A2(n20), .ZN(n137) );
  NAND3_X1 U128 ( .A1(n162), .A2(n163), .A3(n19), .ZN(n161) );
  NOR2_X1 U129 ( .A1(n20), .A2(A[19]), .ZN(n84) );
  NAND3_X1 U130 ( .A1(n164), .A2(n89), .A3(n88), .ZN(n162) );
  AND2_X1 U131 ( .A1(n163), .A2(n136), .ZN(n88) );
  NAND2_X1 U132 ( .A1(A[18]), .A2(n21), .ZN(n136) );
  OR2_X1 U133 ( .A1(n21), .A2(A[18]), .ZN(n163) );
  NAND2_X1 U134 ( .A1(A[17]), .A2(n22), .ZN(n89) );
  NAND3_X1 U135 ( .A1(n165), .A2(n166), .A3(n87), .ZN(n164) );
  OR2_X1 U136 ( .A1(n22), .A2(A[17]), .ZN(n87) );
  NAND3_X1 U137 ( .A1(n167), .A2(n135), .A3(n23), .ZN(n165) );
  NAND2_X1 U138 ( .A1(n166), .A2(n90), .ZN(n93) );
  NAND2_X1 U139 ( .A1(A[16]), .A2(n24), .ZN(n90) );
  OR2_X1 U140 ( .A1(n24), .A2(A[16]), .ZN(n166) );
  NAND2_X1 U141 ( .A1(A[15]), .A2(n26), .ZN(n135) );
  NAND3_X1 U142 ( .A1(n168), .A2(n169), .A3(n25), .ZN(n167) );
  NOR2_X1 U143 ( .A1(n26), .A2(A[15]), .ZN(n94) );
  NAND3_X1 U144 ( .A1(n170), .A2(n99), .A3(n98), .ZN(n168) );
  AND2_X1 U145 ( .A1(n169), .A2(n134), .ZN(n98) );
  NAND2_X1 U146 ( .A1(A[14]), .A2(n27), .ZN(n134) );
  OR2_X1 U147 ( .A1(n27), .A2(A[14]), .ZN(n169) );
  NAND2_X1 U148 ( .A1(A[13]), .A2(n28), .ZN(n99) );
  NAND3_X1 U149 ( .A1(n171), .A2(n172), .A3(n97), .ZN(n170) );
  OR2_X1 U150 ( .A1(n28), .A2(A[13]), .ZN(n97) );
  NAND3_X1 U151 ( .A1(n173), .A2(n133), .A3(n29), .ZN(n171) );
  NAND2_X1 U152 ( .A1(n172), .A2(n100), .ZN(n103) );
  NAND2_X1 U153 ( .A1(A[12]), .A2(n30), .ZN(n100) );
  OR2_X1 U154 ( .A1(n30), .A2(A[12]), .ZN(n172) );
  NAND2_X1 U155 ( .A1(A[11]), .A2(n32), .ZN(n133) );
  NAND3_X1 U156 ( .A1(n174), .A2(n175), .A3(n31), .ZN(n173) );
  NOR2_X1 U157 ( .A1(n32), .A2(A[11]), .ZN(n104) );
  NAND3_X1 U158 ( .A1(n176), .A2(n109), .A3(n108), .ZN(n174) );
  AND2_X1 U159 ( .A1(n175), .A2(n132), .ZN(n108) );
  NAND2_X1 U160 ( .A1(A[10]), .A2(n33), .ZN(n132) );
  OR2_X1 U161 ( .A1(n33), .A2(A[10]), .ZN(n175) );
  NAND2_X1 U162 ( .A1(A[9]), .A2(n34), .ZN(n109) );
  NAND3_X1 U163 ( .A1(n177), .A2(n178), .A3(n107), .ZN(n176) );
  OR2_X1 U164 ( .A1(n34), .A2(A[9]), .ZN(n107) );
  NAND3_X1 U165 ( .A1(n179), .A2(n131), .A3(n35), .ZN(n177) );
  NAND2_X1 U166 ( .A1(n178), .A2(n110), .ZN(n113) );
  NAND2_X1 U167 ( .A1(A[8]), .A2(n36), .ZN(n110) );
  OR2_X1 U168 ( .A1(n36), .A2(A[8]), .ZN(n178) );
  NAND2_X1 U169 ( .A1(A[7]), .A2(n38), .ZN(n131) );
  NAND3_X1 U170 ( .A1(n180), .A2(n181), .A3(n37), .ZN(n179) );
  NOR2_X1 U171 ( .A1(n38), .A2(A[7]), .ZN(n114) );
  NAND3_X1 U172 ( .A1(n182), .A2(n119), .A3(n118), .ZN(n180) );
  AND2_X1 U173 ( .A1(n181), .A2(n130), .ZN(n118) );
  NAND2_X1 U174 ( .A1(A[6]), .A2(n39), .ZN(n130) );
  OR2_X1 U175 ( .A1(n39), .A2(A[6]), .ZN(n181) );
  NAND2_X1 U176 ( .A1(A[5]), .A2(n40), .ZN(n119) );
  NAND3_X1 U177 ( .A1(n183), .A2(n184), .A3(n117), .ZN(n182) );
  OR2_X1 U178 ( .A1(n40), .A2(A[5]), .ZN(n117) );
  NAND3_X1 U179 ( .A1(n185), .A2(n129), .A3(n41), .ZN(n183) );
  NAND2_X1 U180 ( .A1(n184), .A2(n120), .ZN(n123) );
  NAND2_X1 U181 ( .A1(A[4]), .A2(n42), .ZN(n120) );
  OR2_X1 U182 ( .A1(n42), .A2(A[4]), .ZN(n184) );
  NAND2_X1 U183 ( .A1(A[3]), .A2(n44), .ZN(n129) );
  NAND3_X1 U184 ( .A1(n186), .A2(n187), .A3(n43), .ZN(n185) );
  NOR2_X1 U185 ( .A1(n44), .A2(A[3]), .ZN(n124) );
  OAI211_X1 U186 ( .C1(n188), .C2(n51), .A(n46), .B(n126), .ZN(n186) );
  AND2_X1 U187 ( .A1(n187), .A2(n128), .ZN(n126) );
  NAND2_X1 U188 ( .A1(A[2]), .A2(n45), .ZN(n128) );
  OR2_X1 U189 ( .A1(n45), .A2(A[2]), .ZN(n187) );
  AOI21_X1 U190 ( .B1(n51), .B2(n188), .A(B[1]), .ZN(n189) );
  NOR2_X1 U191 ( .A1(n48), .A2(A[0]), .ZN(n188) );
endmodule


module ALU_DATA_W32_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301;

  INV_X2 U3 ( .A(n167), .ZN(n165) );
  INV_X2 U4 ( .A(n287), .ZN(n283) );
  XNOR2_X1 U5 ( .A(n1), .B(n2), .ZN(DIFF[9]) );
  INV_X2 U6 ( .A(n3), .ZN(n2) );
  NAND2_X2 U7 ( .A1(n4), .A2(n5), .ZN(n3) );
  XNOR2_X1 U8 ( .A(n6), .B(n7), .ZN(DIFF[8]) );
  NAND2_X2 U9 ( .A1(n8), .A2(n9), .ZN(n6) );
  XNOR2_X2 U10 ( .A(n10), .B(n11), .ZN(DIFF[7]) );
  INV_X2 U11 ( .A(n12), .ZN(n11) );
  NAND2_X2 U12 ( .A1(n13), .A2(n14), .ZN(n12) );
  AOI21_X2 U13 ( .B1(n15), .B2(n16), .A(n17), .ZN(n10) );
  XNOR2_X2 U14 ( .A(n18), .B(n16), .ZN(DIFF[6]) );
  OAI21_X2 U15 ( .B1(n19), .B2(n20), .A(n21), .ZN(n16) );
  INV_X1 U16 ( .A(n22), .ZN(n20) );
  INV_X1 U17 ( .A(n23), .ZN(n19) );
  NAND2_X2 U18 ( .A1(n15), .A2(n24), .ZN(n18) );
  XNOR2_X1 U19 ( .A(n25), .B(n23), .ZN(DIFF[5]) );
  OAI21_X2 U20 ( .B1(n26), .B2(n27), .A(n28), .ZN(n23) );
  INV_X1 U21 ( .A(n29), .ZN(n26) );
  NAND2_X2 U22 ( .A1(n22), .A2(n21), .ZN(n25) );
  XNOR2_X2 U23 ( .A(n30), .B(n31), .ZN(DIFF[4]) );
  NAND2_X2 U24 ( .A1(n28), .A2(n29), .ZN(n30) );
  XNOR2_X2 U25 ( .A(n32), .B(n33), .ZN(DIFF[3]) );
  NAND2_X2 U26 ( .A1(n34), .A2(n35), .ZN(n33) );
  NAND2_X2 U27 ( .A1(n36), .A2(n37), .ZN(n32) );
  NAND2_X2 U28 ( .A1(n38), .A2(n39), .ZN(n37) );
  XNOR2_X2 U29 ( .A(n40), .B(n41), .ZN(DIFF[31]) );
  XNOR2_X2 U30 ( .A(B[31]), .B(A[31]), .ZN(n41) );
  AOI21_X1 U31 ( .B1(n42), .B2(n43), .A(n44), .ZN(n40) );
  XNOR2_X2 U32 ( .A(n45), .B(n46), .ZN(DIFF[30]) );
  NOR2_X2 U33 ( .A1(n47), .A2(n44), .ZN(n46) );
  INV_X1 U34 ( .A(n48), .ZN(n44) );
  NAND2_X2 U35 ( .A1(A[30]), .A2(n49), .ZN(n48) );
  INV_X2 U36 ( .A(B[30]), .ZN(n49) );
  INV_X1 U37 ( .A(n43), .ZN(n47) );
  NAND2_X2 U38 ( .A1(B[30]), .A2(n50), .ZN(n43) );
  INV_X2 U39 ( .A(A[30]), .ZN(n50) );
  INV_X1 U40 ( .A(n42), .ZN(n45) );
  OAI21_X2 U41 ( .B1(n51), .B2(n52), .A(n53), .ZN(n42) );
  INV_X1 U42 ( .A(n54), .ZN(n51) );
  XNOR2_X2 U43 ( .A(n55), .B(n38), .ZN(DIFF[2]) );
  NAND2_X2 U44 ( .A1(n56), .A2(n57), .ZN(n38) );
  NAND2_X2 U45 ( .A1(n58), .A2(n59), .ZN(n56) );
  NAND2_X2 U46 ( .A1(n39), .A2(n36), .ZN(n55) );
  XNOR2_X2 U47 ( .A(n60), .B(n61), .ZN(DIFF[29]) );
  INV_X2 U48 ( .A(n52), .ZN(n61) );
  AND2_X2 U49 ( .A1(n62), .A2(n63), .ZN(n52) );
  NAND2_X2 U50 ( .A1(n64), .A2(n65), .ZN(n62) );
  NAND2_X2 U51 ( .A1(n53), .A2(n54), .ZN(n60) );
  NAND2_X2 U52 ( .A1(B[29]), .A2(n66), .ZN(n54) );
  INV_X2 U53 ( .A(A[29]), .ZN(n66) );
  NAND2_X2 U54 ( .A1(A[29]), .A2(n67), .ZN(n53) );
  INV_X2 U55 ( .A(B[29]), .ZN(n67) );
  XNOR2_X2 U56 ( .A(n68), .B(n69), .ZN(DIFF[28]) );
  NOR2_X2 U57 ( .A1(n70), .A2(n71), .ZN(n69) );
  INV_X1 U58 ( .A(n63), .ZN(n71) );
  NAND2_X2 U59 ( .A1(A[28]), .A2(n72), .ZN(n63) );
  INV_X2 U60 ( .A(B[28]), .ZN(n72) );
  INV_X1 U61 ( .A(n65), .ZN(n70) );
  NAND2_X2 U62 ( .A1(B[28]), .A2(n73), .ZN(n65) );
  INV_X2 U63 ( .A(A[28]), .ZN(n73) );
  INV_X1 U64 ( .A(n64), .ZN(n68) );
  OAI21_X2 U65 ( .B1(n74), .B2(n75), .A(n76), .ZN(n64) );
  AOI21_X2 U66 ( .B1(n77), .B2(n78), .A(n79), .ZN(n76) );
  OAI21_X2 U67 ( .B1(n80), .B2(n81), .A(n82), .ZN(n78) );
  INV_X1 U68 ( .A(n83), .ZN(n81) );
  AOI21_X2 U69 ( .B1(n84), .B2(n85), .A(n86), .ZN(n80) );
  INV_X1 U70 ( .A(n87), .ZN(n86) );
  INV_X1 U71 ( .A(n88), .ZN(n84) );
  NAND3_X1 U72 ( .A1(n83), .A2(n77), .A3(n85), .ZN(n75) );
  XNOR2_X2 U73 ( .A(n89), .B(n90), .ZN(DIFF[27]) );
  NOR2_X1 U74 ( .A1(n91), .A2(n79), .ZN(n90) );
  INV_X1 U75 ( .A(n92), .ZN(n79) );
  NAND2_X2 U76 ( .A1(A[27]), .A2(n93), .ZN(n92) );
  INV_X2 U77 ( .A(B[27]), .ZN(n93) );
  INV_X1 U78 ( .A(n77), .ZN(n91) );
  NAND2_X2 U79 ( .A1(B[27]), .A2(n94), .ZN(n77) );
  INV_X2 U80 ( .A(A[27]), .ZN(n94) );
  AOI21_X2 U81 ( .B1(n83), .B2(n95), .A(n96), .ZN(n89) );
  INV_X1 U82 ( .A(n82), .ZN(n96) );
  XNOR2_X2 U83 ( .A(n95), .B(n97), .ZN(DIFF[26]) );
  NAND2_X2 U84 ( .A1(n82), .A2(n83), .ZN(n97) );
  NAND2_X2 U85 ( .A1(B[26]), .A2(n98), .ZN(n83) );
  INV_X2 U86 ( .A(A[26]), .ZN(n98) );
  NAND2_X2 U87 ( .A1(A[26]), .A2(n99), .ZN(n82) );
  INV_X2 U88 ( .A(B[26]), .ZN(n99) );
  NAND2_X2 U89 ( .A1(n100), .A2(n87), .ZN(n95) );
  NAND2_X2 U90 ( .A1(n85), .A2(n101), .ZN(n100) );
  XNOR2_X2 U91 ( .A(n102), .B(n101), .ZN(DIFF[25]) );
  NAND2_X2 U92 ( .A1(n74), .A2(n88), .ZN(n101) );
  NAND2_X2 U93 ( .A1(n103), .A2(n104), .ZN(n74) );
  NAND2_X2 U94 ( .A1(n87), .A2(n85), .ZN(n102) );
  NAND2_X2 U95 ( .A1(B[25]), .A2(n105), .ZN(n85) );
  INV_X2 U96 ( .A(A[25]), .ZN(n105) );
  NAND2_X2 U97 ( .A1(A[25]), .A2(n106), .ZN(n87) );
  INV_X2 U98 ( .A(B[25]), .ZN(n106) );
  XNOR2_X2 U99 ( .A(n107), .B(n108), .ZN(DIFF[24]) );
  INV_X2 U100 ( .A(n109), .ZN(n108) );
  NAND2_X2 U101 ( .A1(n88), .A2(n104), .ZN(n109) );
  NAND2_X2 U102 ( .A1(B[24]), .A2(n110), .ZN(n104) );
  INV_X2 U103 ( .A(A[24]), .ZN(n110) );
  NAND2_X2 U104 ( .A1(A[24]), .A2(n111), .ZN(n88) );
  INV_X2 U105 ( .A(B[24]), .ZN(n111) );
  INV_X1 U106 ( .A(n103), .ZN(n107) );
  OAI21_X2 U107 ( .B1(n112), .B2(n113), .A(n114), .ZN(n103) );
  AOI21_X2 U108 ( .B1(n115), .B2(n116), .A(n117), .ZN(n114) );
  OAI21_X2 U109 ( .B1(n118), .B2(n119), .A(n120), .ZN(n116) );
  INV_X1 U110 ( .A(n121), .ZN(n119) );
  AOI21_X2 U111 ( .B1(n122), .B2(n123), .A(n124), .ZN(n118) );
  INV_X1 U112 ( .A(n125), .ZN(n124) );
  INV_X1 U113 ( .A(n126), .ZN(n122) );
  NAND3_X1 U114 ( .A1(n121), .A2(n115), .A3(n123), .ZN(n113) );
  XNOR2_X2 U115 ( .A(n127), .B(n128), .ZN(DIFF[23]) );
  NOR2_X1 U116 ( .A1(n129), .A2(n117), .ZN(n128) );
  INV_X1 U117 ( .A(n130), .ZN(n117) );
  NAND2_X2 U118 ( .A1(A[23]), .A2(n131), .ZN(n130) );
  INV_X2 U119 ( .A(B[23]), .ZN(n131) );
  INV_X1 U120 ( .A(n115), .ZN(n129) );
  NAND2_X2 U121 ( .A1(B[23]), .A2(n132), .ZN(n115) );
  INV_X2 U122 ( .A(A[23]), .ZN(n132) );
  AOI21_X2 U123 ( .B1(n121), .B2(n133), .A(n134), .ZN(n127) );
  INV_X1 U124 ( .A(n120), .ZN(n134) );
  XNOR2_X2 U125 ( .A(n133), .B(n135), .ZN(DIFF[22]) );
  NAND2_X2 U126 ( .A1(n120), .A2(n121), .ZN(n135) );
  NAND2_X2 U127 ( .A1(B[22]), .A2(n136), .ZN(n121) );
  INV_X2 U128 ( .A(A[22]), .ZN(n136) );
  NAND2_X2 U129 ( .A1(A[22]), .A2(n137), .ZN(n120) );
  INV_X2 U130 ( .A(B[22]), .ZN(n137) );
  NAND2_X2 U131 ( .A1(n138), .A2(n125), .ZN(n133) );
  NAND2_X2 U132 ( .A1(n123), .A2(n139), .ZN(n138) );
  XNOR2_X2 U133 ( .A(n140), .B(n139), .ZN(DIFF[21]) );
  NAND2_X2 U134 ( .A1(n112), .A2(n126), .ZN(n139) );
  NAND2_X2 U135 ( .A1(n141), .A2(n142), .ZN(n112) );
  NAND2_X2 U136 ( .A1(n125), .A2(n123), .ZN(n140) );
  NAND2_X2 U137 ( .A1(B[21]), .A2(n143), .ZN(n123) );
  INV_X2 U138 ( .A(A[21]), .ZN(n143) );
  NAND2_X2 U139 ( .A1(A[21]), .A2(n144), .ZN(n125) );
  INV_X2 U140 ( .A(B[21]), .ZN(n144) );
  XNOR2_X1 U141 ( .A(n145), .B(n141), .ZN(DIFF[20]) );
  OAI21_X2 U142 ( .B1(n146), .B2(n147), .A(n148), .ZN(n141) );
  AOI21_X2 U143 ( .B1(n149), .B2(n150), .A(n151), .ZN(n148) );
  INV_X1 U144 ( .A(n152), .ZN(n151) );
  OAI21_X2 U145 ( .B1(n153), .B2(n154), .A(n155), .ZN(n150) );
  AOI21_X2 U146 ( .B1(n156), .B2(n157), .A(n158), .ZN(n153) );
  INV_X1 U147 ( .A(n159), .ZN(n158) );
  INV_X1 U148 ( .A(n160), .ZN(n156) );
  NAND3_X1 U149 ( .A1(n161), .A2(n149), .A3(n157), .ZN(n147) );
  NAND2_X2 U150 ( .A1(n126), .A2(n142), .ZN(n145) );
  NAND2_X2 U151 ( .A1(B[20]), .A2(n162), .ZN(n142) );
  INV_X2 U152 ( .A(A[20]), .ZN(n162) );
  NAND2_X2 U153 ( .A1(A[20]), .A2(n163), .ZN(n126) );
  INV_X2 U154 ( .A(B[20]), .ZN(n163) );
  XNOR2_X2 U155 ( .A(n164), .B(n59), .ZN(DIFF[1]) );
  NAND2_X2 U156 ( .A1(n165), .A2(n166), .ZN(n59) );
  NAND2_X2 U157 ( .A1(n58), .A2(n57), .ZN(n164) );
  XNOR2_X2 U158 ( .A(n168), .B(n169), .ZN(DIFF[19]) );
  OAI21_X2 U159 ( .B1(n170), .B2(n154), .A(n155), .ZN(n169) );
  INV_X1 U160 ( .A(n161), .ZN(n154) );
  INV_X1 U161 ( .A(n171), .ZN(n170) );
  NAND2_X2 U162 ( .A1(n152), .A2(n149), .ZN(n168) );
  NAND2_X2 U163 ( .A1(B[19]), .A2(n172), .ZN(n149) );
  INV_X2 U164 ( .A(A[19]), .ZN(n172) );
  NAND2_X2 U165 ( .A1(A[19]), .A2(n173), .ZN(n152) );
  INV_X2 U166 ( .A(B[19]), .ZN(n173) );
  XNOR2_X2 U167 ( .A(n174), .B(n171), .ZN(DIFF[18]) );
  NAND2_X2 U168 ( .A1(n175), .A2(n159), .ZN(n171) );
  NAND2_X2 U169 ( .A1(n157), .A2(n176), .ZN(n175) );
  NAND2_X2 U170 ( .A1(n155), .A2(n161), .ZN(n174) );
  NAND2_X2 U171 ( .A1(B[18]), .A2(n177), .ZN(n161) );
  INV_X2 U172 ( .A(A[18]), .ZN(n177) );
  NAND2_X2 U173 ( .A1(A[18]), .A2(n178), .ZN(n155) );
  INV_X2 U174 ( .A(B[18]), .ZN(n178) );
  XNOR2_X2 U175 ( .A(n179), .B(n176), .ZN(DIFF[17]) );
  NAND2_X2 U176 ( .A1(n146), .A2(n160), .ZN(n176) );
  NAND2_X2 U177 ( .A1(n180), .A2(n181), .ZN(n146) );
  NAND2_X2 U178 ( .A1(n159), .A2(n157), .ZN(n179) );
  NAND2_X2 U179 ( .A1(B[17]), .A2(n182), .ZN(n157) );
  INV_X2 U180 ( .A(A[17]), .ZN(n182) );
  NAND2_X2 U181 ( .A1(A[17]), .A2(n183), .ZN(n159) );
  INV_X2 U182 ( .A(B[17]), .ZN(n183) );
  XNOR2_X2 U183 ( .A(n180), .B(n184), .ZN(DIFF[16]) );
  NAND2_X2 U184 ( .A1(n160), .A2(n181), .ZN(n184) );
  NAND2_X2 U185 ( .A1(B[16]), .A2(n185), .ZN(n181) );
  INV_X2 U186 ( .A(A[16]), .ZN(n185) );
  NAND2_X2 U187 ( .A1(A[16]), .A2(n186), .ZN(n160) );
  INV_X2 U188 ( .A(B[16]), .ZN(n186) );
  NAND2_X2 U189 ( .A1(n187), .A2(n188), .ZN(n180) );
  OAI21_X2 U190 ( .B1(n189), .B2(n190), .A(n191), .ZN(n188) );
  NOR2_X2 U191 ( .A1(n192), .A2(n193), .ZN(n189) );
  AOI21_X2 U192 ( .B1(n194), .B2(n195), .A(n196), .ZN(n192) );
  NOR2_X2 U193 ( .A1(n197), .A2(n198), .ZN(n187) );
  NAND2_X2 U194 ( .A1(n199), .A2(n200), .ZN(n198) );
  OAI21_X2 U195 ( .B1(n201), .B2(n202), .A(n203), .ZN(n199) );
  NOR2_X2 U196 ( .A1(n204), .A2(n205), .ZN(n202) );
  AOI21_X2 U197 ( .B1(n206), .B2(n207), .A(n208), .ZN(n204) );
  INV_X1 U198 ( .A(n209), .ZN(n208) );
  INV_X1 U199 ( .A(n210), .ZN(n206) );
  INV_X1 U200 ( .A(n211), .ZN(n201) );
  NOR2_X2 U201 ( .A1(n212), .A2(n213), .ZN(n197) );
  NAND2_X1 U202 ( .A1(n214), .A2(n191), .ZN(n213) );
  INV_X1 U203 ( .A(n215), .ZN(n191) );
  NAND4_X2 U204 ( .A1(n216), .A2(n207), .A3(n217), .A4(n203), .ZN(n215) );
  INV_X1 U205 ( .A(n193), .ZN(n214) );
  NAND2_X1 U206 ( .A1(n218), .A2(n194), .ZN(n212) );
  INV_X1 U207 ( .A(n219), .ZN(n194) );
  INV_X1 U208 ( .A(n220), .ZN(n218) );
  XNOR2_X2 U209 ( .A(n221), .B(n222), .ZN(DIFF[15]) );
  OAI21_X2 U210 ( .B1(n223), .B2(n205), .A(n211), .ZN(n222) );
  INV_X1 U211 ( .A(n217), .ZN(n205) );
  INV_X1 U212 ( .A(n224), .ZN(n223) );
  NAND2_X2 U213 ( .A1(n200), .A2(n203), .ZN(n221) );
  NAND2_X2 U214 ( .A1(B[15]), .A2(n225), .ZN(n203) );
  INV_X2 U215 ( .A(A[15]), .ZN(n225) );
  NAND2_X2 U216 ( .A1(A[15]), .A2(n226), .ZN(n200) );
  INV_X2 U217 ( .A(B[15]), .ZN(n226) );
  XNOR2_X2 U218 ( .A(n227), .B(n224), .ZN(DIFF[14]) );
  OAI21_X2 U219 ( .B1(n228), .B2(n229), .A(n209), .ZN(n224) );
  INV_X1 U220 ( .A(n207), .ZN(n229) );
  INV_X1 U221 ( .A(n230), .ZN(n228) );
  NAND2_X2 U222 ( .A1(n211), .A2(n217), .ZN(n227) );
  NAND2_X2 U223 ( .A1(B[14]), .A2(n231), .ZN(n217) );
  INV_X2 U224 ( .A(A[14]), .ZN(n231) );
  NAND2_X2 U225 ( .A1(A[14]), .A2(n232), .ZN(n211) );
  INV_X2 U226 ( .A(B[14]), .ZN(n232) );
  XNOR2_X1 U227 ( .A(n233), .B(n230), .ZN(DIFF[13]) );
  OAI21_X2 U228 ( .B1(n234), .B2(n235), .A(n210), .ZN(n230) );
  INV_X1 U229 ( .A(n236), .ZN(n235) );
  INV_X1 U230 ( .A(n216), .ZN(n234) );
  NAND2_X2 U231 ( .A1(n209), .A2(n207), .ZN(n233) );
  NAND2_X2 U232 ( .A1(B[13]), .A2(n237), .ZN(n207) );
  INV_X2 U233 ( .A(A[13]), .ZN(n237) );
  NAND2_X2 U234 ( .A1(A[13]), .A2(n238), .ZN(n209) );
  INV_X2 U235 ( .A(B[13]), .ZN(n238) );
  XNOR2_X2 U236 ( .A(n239), .B(n236), .ZN(DIFF[12]) );
  OAI21_X2 U237 ( .B1(n240), .B2(n193), .A(n241), .ZN(n236) );
  INV_X1 U238 ( .A(n190), .ZN(n241) );
  NAND2_X2 U239 ( .A1(n242), .A2(n243), .ZN(n190) );
  OAI21_X2 U240 ( .B1(n244), .B2(n245), .A(n246), .ZN(n242) );
  INV_X2 U241 ( .A(n247), .ZN(n245) );
  AOI21_X2 U242 ( .B1(n5), .B2(n248), .A(n249), .ZN(n244) );
  NAND2_X2 U243 ( .A1(n250), .A2(n4), .ZN(n248) );
  INV_X2 U244 ( .A(n8), .ZN(n250) );
  NAND4_X2 U245 ( .A1(n246), .A2(n251), .A3(n4), .A4(n9), .ZN(n193) );
  INV_X1 U246 ( .A(n7), .ZN(n240) );
  NAND2_X2 U247 ( .A1(n210), .A2(n216), .ZN(n239) );
  NAND2_X2 U248 ( .A1(B[12]), .A2(n252), .ZN(n216) );
  INV_X2 U249 ( .A(A[12]), .ZN(n252) );
  NAND2_X2 U250 ( .A1(A[12]), .A2(n253), .ZN(n210) );
  INV_X2 U251 ( .A(B[12]), .ZN(n253) );
  XNOR2_X1 U252 ( .A(n254), .B(n255), .ZN(DIFF[11]) );
  OAI21_X2 U253 ( .B1(n256), .B2(n249), .A(n247), .ZN(n255) );
  INV_X1 U254 ( .A(n251), .ZN(n249) );
  NAND2_X2 U255 ( .A1(n243), .A2(n246), .ZN(n254) );
  NAND2_X2 U256 ( .A1(B[11]), .A2(n257), .ZN(n246) );
  INV_X2 U257 ( .A(A[11]), .ZN(n257) );
  NAND2_X2 U258 ( .A1(A[11]), .A2(n258), .ZN(n243) );
  INV_X2 U259 ( .A(B[11]), .ZN(n258) );
  XNOR2_X1 U260 ( .A(n256), .B(n259), .ZN(DIFF[10]) );
  INV_X2 U261 ( .A(n260), .ZN(n259) );
  NAND2_X2 U262 ( .A1(n247), .A2(n251), .ZN(n260) );
  NAND2_X2 U263 ( .A1(B[10]), .A2(n261), .ZN(n251) );
  INV_X2 U264 ( .A(A[10]), .ZN(n261) );
  NAND2_X2 U265 ( .A1(A[10]), .A2(n262), .ZN(n247) );
  INV_X2 U266 ( .A(B[10]), .ZN(n262) );
  INV_X1 U267 ( .A(n263), .ZN(n256) );
  OAI21_X2 U268 ( .B1(n264), .B2(n1), .A(n5), .ZN(n263) );
  NAND2_X2 U269 ( .A1(A[9]), .A2(n265), .ZN(n5) );
  INV_X2 U270 ( .A(B[9]), .ZN(n265) );
  AND2_X2 U271 ( .A1(n266), .A2(n8), .ZN(n1) );
  NAND2_X2 U272 ( .A1(A[8]), .A2(n267), .ZN(n8) );
  INV_X2 U273 ( .A(B[8]), .ZN(n267) );
  NAND2_X2 U274 ( .A1(n7), .A2(n9), .ZN(n266) );
  NAND2_X2 U275 ( .A1(B[8]), .A2(n268), .ZN(n9) );
  INV_X2 U276 ( .A(A[8]), .ZN(n268) );
  OAI21_X2 U277 ( .B1(n27), .B2(n219), .A(n269), .ZN(n7) );
  INV_X1 U278 ( .A(n196), .ZN(n269) );
  NAND2_X2 U279 ( .A1(n270), .A2(n271), .ZN(n196) );
  NAND4_X2 U280 ( .A1(n272), .A2(n22), .A3(n15), .A4(n13), .ZN(n271) );
  NAND2_X2 U281 ( .A1(n21), .A2(n28), .ZN(n272) );
  NAND2_X2 U282 ( .A1(A[4]), .A2(n273), .ZN(n28) );
  INV_X2 U283 ( .A(B[4]), .ZN(n273) );
  NAND2_X2 U284 ( .A1(A[5]), .A2(n274), .ZN(n21) );
  INV_X2 U285 ( .A(B[5]), .ZN(n274) );
  AOI21_X2 U286 ( .B1(n17), .B2(n13), .A(n275), .ZN(n270) );
  INV_X1 U287 ( .A(n14), .ZN(n275) );
  NAND2_X2 U288 ( .A1(A[7]), .A2(n276), .ZN(n14) );
  INV_X2 U289 ( .A(B[7]), .ZN(n276) );
  INV_X1 U290 ( .A(n24), .ZN(n17) );
  NAND2_X2 U291 ( .A1(A[6]), .A2(n277), .ZN(n24) );
  INV_X2 U292 ( .A(B[6]), .ZN(n277) );
  NAND4_X2 U293 ( .A1(n29), .A2(n22), .A3(n15), .A4(n13), .ZN(n219) );
  NAND2_X2 U294 ( .A1(B[7]), .A2(n278), .ZN(n13) );
  INV_X2 U295 ( .A(A[7]), .ZN(n278) );
  NAND2_X2 U296 ( .A1(B[6]), .A2(n279), .ZN(n15) );
  INV_X2 U297 ( .A(A[6]), .ZN(n279) );
  NAND2_X2 U298 ( .A1(B[5]), .A2(n280), .ZN(n22) );
  INV_X2 U299 ( .A(A[5]), .ZN(n280) );
  NAND2_X2 U300 ( .A1(B[4]), .A2(n281), .ZN(n29) );
  INV_X2 U301 ( .A(A[4]), .ZN(n281) );
  INV_X1 U302 ( .A(n31), .ZN(n27) );
  NAND2_X2 U303 ( .A1(n282), .A2(n220), .ZN(n31) );
  NAND3_X1 U304 ( .A1(n283), .A2(n39), .A3(n284), .ZN(n220) );
  NOR2_X1 U305 ( .A1(n285), .A2(n286), .ZN(n284) );
  INV_X1 U306 ( .A(n167), .ZN(n286) );
  INV_X1 U307 ( .A(n58), .ZN(n285) );
  INV_X1 U308 ( .A(n34), .ZN(n287) );
  INV_X1 U309 ( .A(n195), .ZN(n282) );
  NAND2_X2 U310 ( .A1(n288), .A2(n289), .ZN(n195) );
  NAND4_X2 U311 ( .A1(n290), .A2(n58), .A3(n39), .A4(n34), .ZN(n289) );
  NAND2_X2 U312 ( .A1(B[2]), .A2(n291), .ZN(n39) );
  INV_X2 U313 ( .A(A[2]), .ZN(n291) );
  NAND2_X2 U314 ( .A1(B[1]), .A2(n292), .ZN(n58) );
  INV_X2 U315 ( .A(A[1]), .ZN(n292) );
  NAND2_X2 U316 ( .A1(n57), .A2(n166), .ZN(n290) );
  NAND2_X2 U317 ( .A1(A[1]), .A2(n293), .ZN(n57) );
  INV_X2 U318 ( .A(B[1]), .ZN(n293) );
  AOI21_X2 U319 ( .B1(n294), .B2(n34), .A(n295), .ZN(n288) );
  INV_X1 U320 ( .A(n35), .ZN(n295) );
  NAND2_X2 U321 ( .A1(A[3]), .A2(n296), .ZN(n35) );
  INV_X2 U322 ( .A(B[3]), .ZN(n296) );
  NAND2_X2 U323 ( .A1(B[3]), .A2(n297), .ZN(n34) );
  INV_X2 U324 ( .A(A[3]), .ZN(n297) );
  INV_X1 U325 ( .A(n36), .ZN(n294) );
  NAND2_X2 U326 ( .A1(A[2]), .A2(n298), .ZN(n36) );
  INV_X2 U327 ( .A(B[2]), .ZN(n298) );
  INV_X1 U328 ( .A(n4), .ZN(n264) );
  NAND2_X2 U329 ( .A1(B[9]), .A2(n299), .ZN(n4) );
  INV_X2 U330 ( .A(A[9]), .ZN(n299) );
  NAND2_X2 U331 ( .A1(n166), .A2(n167), .ZN(DIFF[0]) );
  NAND2_X2 U332 ( .A1(B[0]), .A2(n300), .ZN(n167) );
  INV_X2 U333 ( .A(A[0]), .ZN(n300) );
  NAND2_X2 U334 ( .A1(A[0]), .A2(n301), .ZN(n166) );
  INV_X2 U335 ( .A(B[0]), .ZN(n301) );
endmodule


module ALU_DATA_W32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282;

  INV_X2 U2 ( .A(n201), .ZN(n26) );
  INV_X2 U3 ( .A(n163), .ZN(n57) );
  INV_X2 U4 ( .A(n184), .ZN(n183) );
  INV_X2 U5 ( .A(n280), .ZN(SUM[0]) );
  XNOR2_X2 U6 ( .A(n1), .B(n2), .ZN(SUM[9]) );
  NAND2_X2 U7 ( .A1(n3), .A2(n4), .ZN(n1) );
  XNOR2_X2 U8 ( .A(n5), .B(n6), .ZN(SUM[8]) );
  NAND2_X2 U9 ( .A1(n7), .A2(n8), .ZN(n5) );
  XNOR2_X2 U10 ( .A(n9), .B(n10), .ZN(SUM[7]) );
  NAND2_X2 U11 ( .A1(n11), .A2(n12), .ZN(n10) );
  NAND2_X2 U12 ( .A1(n13), .A2(n14), .ZN(n11) );
  NAND2_X2 U13 ( .A1(n15), .A2(n16), .ZN(n9) );
  XNOR2_X2 U14 ( .A(n17), .B(n14), .ZN(SUM[6]) );
  OAI21_X2 U15 ( .B1(n18), .B2(n19), .A(n20), .ZN(n14) );
  INV_X1 U16 ( .A(n21), .ZN(n19) );
  INV_X1 U17 ( .A(n22), .ZN(n18) );
  NAND2_X2 U18 ( .A1(n13), .A2(n12), .ZN(n17) );
  XNOR2_X2 U19 ( .A(n23), .B(n22), .ZN(SUM[5]) );
  NAND2_X2 U20 ( .A1(n24), .A2(n25), .ZN(n22) );
  NAND2_X2 U21 ( .A1(n26), .A2(n27), .ZN(n24) );
  NAND2_X2 U22 ( .A1(n21), .A2(n20), .ZN(n23) );
  XNOR2_X2 U23 ( .A(n28), .B(n26), .ZN(SUM[4]) );
  NAND2_X2 U24 ( .A1(n25), .A2(n27), .ZN(n28) );
  XNOR2_X2 U25 ( .A(n29), .B(n30), .ZN(SUM[3]) );
  OAI21_X2 U26 ( .B1(n31), .B2(n32), .A(n33), .ZN(n30) );
  INV_X1 U27 ( .A(n34), .ZN(n31) );
  NAND2_X2 U28 ( .A1(n35), .A2(n36), .ZN(n29) );
  XNOR2_X2 U29 ( .A(n37), .B(n38), .ZN(SUM[31]) );
  INV_X2 U30 ( .A(n39), .ZN(n38) );
  XNOR2_X2 U31 ( .A(B[31]), .B(A[31]), .ZN(n39) );
  AOI21_X1 U32 ( .B1(n40), .B2(n41), .A(n42), .ZN(n37) );
  INV_X1 U33 ( .A(n43), .ZN(n42) );
  XNOR2_X2 U34 ( .A(n44), .B(n45), .ZN(SUM[30]) );
  INV_X2 U35 ( .A(n46), .ZN(n45) );
  NAND2_X2 U36 ( .A1(n43), .A2(n41), .ZN(n46) );
  NAND2_X2 U37 ( .A1(n47), .A2(n48), .ZN(n41) );
  INV_X2 U38 ( .A(A[30]), .ZN(n48) );
  INV_X2 U39 ( .A(B[30]), .ZN(n47) );
  NAND2_X2 U40 ( .A1(B[30]), .A2(A[30]), .ZN(n43) );
  INV_X1 U41 ( .A(n40), .ZN(n44) );
  OAI21_X2 U42 ( .B1(n49), .B2(n50), .A(n51), .ZN(n40) );
  INV_X1 U43 ( .A(n52), .ZN(n49) );
  XNOR2_X2 U44 ( .A(n53), .B(n34), .ZN(SUM[2]) );
  NAND2_X2 U45 ( .A1(n54), .A2(n55), .ZN(n34) );
  NAND2_X2 U46 ( .A1(n56), .A2(n57), .ZN(n54) );
  NAND2_X2 U47 ( .A1(n58), .A2(n33), .ZN(n53) );
  XNOR2_X2 U48 ( .A(n59), .B(n60), .ZN(SUM[29]) );
  INV_X2 U49 ( .A(n50), .ZN(n60) );
  AND2_X2 U50 ( .A1(n61), .A2(n62), .ZN(n50) );
  NAND2_X2 U51 ( .A1(n63), .A2(n64), .ZN(n61) );
  NAND2_X2 U52 ( .A1(n51), .A2(n52), .ZN(n59) );
  NAND2_X2 U53 ( .A1(n65), .A2(n66), .ZN(n52) );
  INV_X2 U54 ( .A(A[29]), .ZN(n66) );
  INV_X2 U55 ( .A(B[29]), .ZN(n65) );
  NAND2_X2 U56 ( .A1(B[29]), .A2(A[29]), .ZN(n51) );
  XNOR2_X2 U57 ( .A(n67), .B(n68), .ZN(SUM[28]) );
  INV_X2 U58 ( .A(n69), .ZN(n68) );
  NAND2_X2 U59 ( .A1(n62), .A2(n64), .ZN(n69) );
  NAND2_X2 U60 ( .A1(n70), .A2(n71), .ZN(n64) );
  INV_X2 U61 ( .A(A[28]), .ZN(n71) );
  INV_X2 U62 ( .A(B[28]), .ZN(n70) );
  NAND2_X2 U63 ( .A1(B[28]), .A2(A[28]), .ZN(n62) );
  INV_X1 U64 ( .A(n63), .ZN(n67) );
  OAI21_X2 U65 ( .B1(n72), .B2(n73), .A(n74), .ZN(n63) );
  NOR2_X2 U66 ( .A1(n75), .A2(n76), .ZN(n74) );
  AOI21_X2 U67 ( .B1(n77), .B2(n78), .A(n79), .ZN(n76) );
  NAND2_X2 U68 ( .A1(n80), .A2(n81), .ZN(n77) );
  OAI21_X2 U69 ( .B1(n82), .B2(n83), .A(n84), .ZN(n81) );
  INV_X1 U70 ( .A(n85), .ZN(n82) );
  NAND3_X1 U71 ( .A1(n80), .A2(n86), .A3(n85), .ZN(n73) );
  XNOR2_X2 U72 ( .A(n87), .B(n88), .ZN(SUM[27]) );
  NOR2_X2 U73 ( .A1(n79), .A2(n75), .ZN(n88) );
  INV_X1 U74 ( .A(n89), .ZN(n75) );
  NAND2_X2 U75 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U76 ( .A(n86), .ZN(n79) );
  NAND2_X2 U77 ( .A1(n90), .A2(n91), .ZN(n86) );
  INV_X2 U78 ( .A(A[27]), .ZN(n91) );
  INV_X2 U79 ( .A(B[27]), .ZN(n90) );
  AOI21_X2 U80 ( .B1(n80), .B2(n92), .A(n93), .ZN(n87) );
  INV_X1 U81 ( .A(n78), .ZN(n93) );
  XNOR2_X2 U82 ( .A(n92), .B(n94), .ZN(SUM[26]) );
  NAND2_X2 U83 ( .A1(n78), .A2(n80), .ZN(n94) );
  NAND2_X2 U84 ( .A1(n95), .A2(n96), .ZN(n80) );
  INV_X2 U85 ( .A(A[26]), .ZN(n96) );
  INV_X2 U86 ( .A(B[26]), .ZN(n95) );
  NAND2_X2 U87 ( .A1(B[26]), .A2(A[26]), .ZN(n78) );
  NAND2_X2 U88 ( .A1(n97), .A2(n84), .ZN(n92) );
  NAND2_X2 U89 ( .A1(n85), .A2(n98), .ZN(n97) );
  XNOR2_X2 U90 ( .A(n99), .B(n98), .ZN(SUM[25]) );
  NAND2_X2 U91 ( .A1(n72), .A2(n83), .ZN(n98) );
  NAND2_X2 U92 ( .A1(n100), .A2(n101), .ZN(n72) );
  NAND2_X2 U93 ( .A1(n84), .A2(n85), .ZN(n99) );
  NAND2_X2 U94 ( .A1(n102), .A2(n103), .ZN(n85) );
  INV_X2 U95 ( .A(A[25]), .ZN(n103) );
  INV_X2 U96 ( .A(B[25]), .ZN(n102) );
  NAND2_X2 U97 ( .A1(B[25]), .A2(A[25]), .ZN(n84) );
  XNOR2_X2 U98 ( .A(n104), .B(n105), .ZN(SUM[24]) );
  INV_X2 U99 ( .A(n106), .ZN(n105) );
  NAND2_X2 U100 ( .A1(n83), .A2(n101), .ZN(n106) );
  NAND2_X2 U101 ( .A1(n107), .A2(n108), .ZN(n101) );
  INV_X2 U102 ( .A(A[24]), .ZN(n108) );
  INV_X2 U103 ( .A(B[24]), .ZN(n107) );
  NAND2_X2 U104 ( .A1(B[24]), .A2(A[24]), .ZN(n83) );
  INV_X1 U105 ( .A(n100), .ZN(n104) );
  OAI21_X2 U106 ( .B1(n109), .B2(n110), .A(n111), .ZN(n100) );
  NOR2_X2 U107 ( .A1(n112), .A2(n113), .ZN(n111) );
  AOI21_X2 U108 ( .B1(n114), .B2(n115), .A(n116), .ZN(n113) );
  NAND2_X2 U109 ( .A1(n117), .A2(n118), .ZN(n114) );
  OAI21_X2 U110 ( .B1(n119), .B2(n120), .A(n121), .ZN(n118) );
  INV_X1 U111 ( .A(n122), .ZN(n119) );
  NAND3_X1 U112 ( .A1(n117), .A2(n123), .A3(n122), .ZN(n110) );
  XNOR2_X2 U113 ( .A(n124), .B(n125), .ZN(SUM[23]) );
  NOR2_X2 U114 ( .A1(n116), .A2(n112), .ZN(n125) );
  INV_X1 U115 ( .A(n126), .ZN(n112) );
  NAND2_X2 U116 ( .A1(B[23]), .A2(A[23]), .ZN(n126) );
  INV_X1 U117 ( .A(n123), .ZN(n116) );
  NAND2_X2 U118 ( .A1(n127), .A2(n128), .ZN(n123) );
  INV_X2 U119 ( .A(A[23]), .ZN(n128) );
  INV_X2 U120 ( .A(B[23]), .ZN(n127) );
  AOI21_X2 U121 ( .B1(n117), .B2(n129), .A(n130), .ZN(n124) );
  INV_X1 U122 ( .A(n115), .ZN(n130) );
  XNOR2_X2 U123 ( .A(n129), .B(n131), .ZN(SUM[22]) );
  NAND2_X2 U124 ( .A1(n115), .A2(n117), .ZN(n131) );
  NAND2_X2 U125 ( .A1(n132), .A2(n133), .ZN(n117) );
  INV_X2 U126 ( .A(A[22]), .ZN(n133) );
  INV_X2 U127 ( .A(B[22]), .ZN(n132) );
  NAND2_X2 U128 ( .A1(B[22]), .A2(A[22]), .ZN(n115) );
  NAND2_X2 U129 ( .A1(n134), .A2(n121), .ZN(n129) );
  NAND2_X2 U130 ( .A1(n122), .A2(n135), .ZN(n134) );
  XNOR2_X2 U131 ( .A(n136), .B(n135), .ZN(SUM[21]) );
  NAND2_X2 U132 ( .A1(n109), .A2(n120), .ZN(n135) );
  NAND2_X2 U133 ( .A1(n137), .A2(n138), .ZN(n109) );
  NAND2_X2 U134 ( .A1(n121), .A2(n122), .ZN(n136) );
  NAND2_X2 U135 ( .A1(n139), .A2(n140), .ZN(n122) );
  INV_X2 U136 ( .A(A[21]), .ZN(n140) );
  INV_X2 U137 ( .A(B[21]), .ZN(n139) );
  NAND2_X2 U138 ( .A1(B[21]), .A2(A[21]), .ZN(n121) );
  XNOR2_X1 U139 ( .A(n141), .B(n142), .ZN(SUM[20]) );
  INV_X2 U140 ( .A(n143), .ZN(n142) );
  NAND2_X2 U141 ( .A1(n120), .A2(n138), .ZN(n143) );
  NAND2_X2 U142 ( .A1(n144), .A2(n145), .ZN(n138) );
  INV_X2 U143 ( .A(A[20]), .ZN(n145) );
  INV_X2 U144 ( .A(B[20]), .ZN(n144) );
  NAND2_X2 U145 ( .A1(B[20]), .A2(A[20]), .ZN(n120) );
  INV_X1 U146 ( .A(n137), .ZN(n141) );
  OAI21_X2 U147 ( .B1(n146), .B2(n147), .A(n148), .ZN(n137) );
  NOR2_X2 U148 ( .A1(n149), .A2(n150), .ZN(n148) );
  AOI21_X2 U149 ( .B1(n151), .B2(n152), .A(n153), .ZN(n150) );
  INV_X1 U150 ( .A(n154), .ZN(n153) );
  NAND2_X2 U151 ( .A1(n155), .A2(n156), .ZN(n151) );
  OAI21_X2 U152 ( .B1(n157), .B2(n158), .A(n159), .ZN(n156) );
  INV_X1 U153 ( .A(n160), .ZN(n157) );
  INV_X1 U154 ( .A(n161), .ZN(n149) );
  NAND3_X1 U155 ( .A1(n155), .A2(n154), .A3(n160), .ZN(n147) );
  XNOR2_X2 U156 ( .A(n162), .B(n57), .ZN(SUM[1]) );
  NAND2_X2 U157 ( .A1(n56), .A2(n55), .ZN(n162) );
  XNOR2_X2 U158 ( .A(n164), .B(n165), .ZN(SUM[19]) );
  NAND2_X2 U159 ( .A1(n161), .A2(n154), .ZN(n165) );
  NAND2_X2 U160 ( .A1(n166), .A2(n167), .ZN(n154) );
  INV_X2 U161 ( .A(A[19]), .ZN(n167) );
  INV_X2 U162 ( .A(B[19]), .ZN(n166) );
  NAND2_X2 U163 ( .A1(B[19]), .A2(A[19]), .ZN(n161) );
  NAND2_X2 U164 ( .A1(n152), .A2(n168), .ZN(n164) );
  NAND2_X2 U165 ( .A1(n169), .A2(n155), .ZN(n168) );
  XNOR2_X2 U166 ( .A(n170), .B(n169), .ZN(SUM[18]) );
  NAND2_X2 U167 ( .A1(n171), .A2(n159), .ZN(n169) );
  NAND2_X2 U168 ( .A1(n160), .A2(n172), .ZN(n171) );
  NAND2_X2 U169 ( .A1(n152), .A2(n155), .ZN(n170) );
  NAND2_X2 U170 ( .A1(n173), .A2(n174), .ZN(n155) );
  INV_X2 U171 ( .A(A[18]), .ZN(n174) );
  INV_X2 U172 ( .A(B[18]), .ZN(n173) );
  NAND2_X2 U173 ( .A1(B[18]), .A2(A[18]), .ZN(n152) );
  XNOR2_X2 U174 ( .A(n175), .B(n172), .ZN(SUM[17]) );
  NAND2_X2 U175 ( .A1(n146), .A2(n158), .ZN(n172) );
  NAND2_X2 U176 ( .A1(n176), .A2(n177), .ZN(n146) );
  NAND2_X2 U177 ( .A1(n159), .A2(n160), .ZN(n175) );
  NAND2_X2 U178 ( .A1(n178), .A2(n179), .ZN(n160) );
  INV_X2 U179 ( .A(A[17]), .ZN(n179) );
  INV_X2 U180 ( .A(B[17]), .ZN(n178) );
  NAND2_X2 U181 ( .A1(B[17]), .A2(A[17]), .ZN(n159) );
  XNOR2_X1 U182 ( .A(n180), .B(n176), .ZN(SUM[16]) );
  OAI21_X2 U183 ( .B1(n181), .B2(n182), .A(n183), .ZN(n176) );
  OAI21_X2 U184 ( .B1(n185), .B2(n186), .A(n187), .ZN(n184) );
  AOI21_X2 U185 ( .B1(n188), .B2(n189), .A(n190), .ZN(n185) );
  OAI21_X2 U186 ( .B1(n191), .B2(n192), .A(n193), .ZN(n189) );
  NAND4_X2 U187 ( .A1(n196), .A2(n197), .A3(n188), .A4(n198), .ZN(n182) );
  AOI21_X2 U188 ( .B1(n194), .B2(n199), .A(n200), .ZN(n181) );
  OAI21_X2 U189 ( .B1(n201), .B2(n195), .A(n202), .ZN(n199) );
  INV_X1 U190 ( .A(n203), .ZN(n194) );
  NAND2_X2 U191 ( .A1(n158), .A2(n177), .ZN(n180) );
  NAND2_X2 U192 ( .A1(n204), .A2(n205), .ZN(n177) );
  INV_X2 U193 ( .A(A[16]), .ZN(n205) );
  INV_X2 U194 ( .A(B[16]), .ZN(n204) );
  NAND2_X2 U195 ( .A1(B[16]), .A2(A[16]), .ZN(n158) );
  XNOR2_X2 U196 ( .A(n206), .B(n207), .ZN(SUM[15]) );
  NOR2_X2 U197 ( .A1(n186), .A2(n208), .ZN(n207) );
  INV_X1 U198 ( .A(n187), .ZN(n208) );
  NAND2_X2 U199 ( .A1(B[15]), .A2(A[15]), .ZN(n187) );
  INV_X1 U200 ( .A(n198), .ZN(n186) );
  NAND2_X2 U201 ( .A1(n209), .A2(n210), .ZN(n198) );
  INV_X2 U202 ( .A(A[15]), .ZN(n210) );
  INV_X2 U203 ( .A(B[15]), .ZN(n209) );
  AOI21_X2 U204 ( .B1(n188), .B2(n211), .A(n190), .ZN(n206) );
  INV_X1 U205 ( .A(n212), .ZN(n190) );
  XNOR2_X2 U206 ( .A(n213), .B(n211), .ZN(SUM[14]) );
  OAI21_X2 U207 ( .B1(n214), .B2(n191), .A(n193), .ZN(n211) );
  INV_X1 U208 ( .A(n197), .ZN(n191) );
  INV_X1 U209 ( .A(n215), .ZN(n214) );
  NAND2_X2 U210 ( .A1(n212), .A2(n188), .ZN(n213) );
  NAND2_X2 U211 ( .A1(n216), .A2(n217), .ZN(n188) );
  INV_X2 U212 ( .A(A[14]), .ZN(n217) );
  INV_X2 U213 ( .A(B[14]), .ZN(n216) );
  NAND2_X2 U214 ( .A1(B[14]), .A2(A[14]), .ZN(n212) );
  XNOR2_X2 U215 ( .A(n218), .B(n215), .ZN(SUM[13]) );
  NAND2_X2 U216 ( .A1(n219), .A2(n192), .ZN(n215) );
  NAND2_X2 U217 ( .A1(n220), .A2(n196), .ZN(n219) );
  NAND2_X2 U218 ( .A1(n193), .A2(n197), .ZN(n218) );
  NAND2_X2 U219 ( .A1(n221), .A2(n222), .ZN(n197) );
  INV_X2 U220 ( .A(A[13]), .ZN(n222) );
  INV_X2 U221 ( .A(B[13]), .ZN(n221) );
  NAND2_X2 U222 ( .A1(B[13]), .A2(A[13]), .ZN(n193) );
  XNOR2_X2 U223 ( .A(n223), .B(n220), .ZN(SUM[12]) );
  OAI21_X2 U224 ( .B1(n224), .B2(n203), .A(n225), .ZN(n220) );
  INV_X1 U225 ( .A(n200), .ZN(n225) );
  OAI21_X2 U226 ( .B1(n226), .B2(n227), .A(n228), .ZN(n200) );
  INV_X1 U227 ( .A(n229), .ZN(n227) );
  AOI21_X2 U228 ( .B1(n230), .B2(n231), .A(n232), .ZN(n226) );
  INV_X1 U229 ( .A(n233), .ZN(n232) );
  OAI21_X2 U230 ( .B1(n234), .B2(n7), .A(n4), .ZN(n231) );
  NAND4_X2 U231 ( .A1(n229), .A2(n230), .A3(n3), .A4(n8), .ZN(n203) );
  INV_X1 U232 ( .A(n6), .ZN(n224) );
  NAND2_X2 U233 ( .A1(n192), .A2(n196), .ZN(n223) );
  NAND2_X2 U234 ( .A1(n235), .A2(n236), .ZN(n196) );
  INV_X2 U235 ( .A(A[12]), .ZN(n236) );
  INV_X2 U236 ( .A(B[12]), .ZN(n235) );
  NAND2_X2 U237 ( .A1(B[12]), .A2(A[12]), .ZN(n192) );
  XNOR2_X2 U238 ( .A(n237), .B(n238), .ZN(SUM[11]) );
  NAND2_X2 U239 ( .A1(n228), .A2(n229), .ZN(n238) );
  NAND2_X2 U240 ( .A1(n239), .A2(n240), .ZN(n229) );
  INV_X2 U241 ( .A(A[11]), .ZN(n240) );
  INV_X2 U242 ( .A(B[11]), .ZN(n239) );
  NAND2_X2 U243 ( .A1(B[11]), .A2(A[11]), .ZN(n228) );
  NAND2_X2 U244 ( .A1(n233), .A2(n241), .ZN(n237) );
  NAND2_X2 U245 ( .A1(n242), .A2(n230), .ZN(n241) );
  XNOR2_X2 U246 ( .A(n243), .B(n242), .ZN(SUM[10]) );
  OAI21_X2 U247 ( .B1(n234), .B2(n244), .A(n4), .ZN(n242) );
  NAND2_X2 U248 ( .A1(B[9]), .A2(A[9]), .ZN(n4) );
  INV_X1 U249 ( .A(n2), .ZN(n244) );
  NAND2_X2 U250 ( .A1(n245), .A2(n7), .ZN(n2) );
  NAND2_X2 U251 ( .A1(B[8]), .A2(A[8]), .ZN(n7) );
  NAND2_X2 U252 ( .A1(n6), .A2(n8), .ZN(n245) );
  NAND2_X2 U253 ( .A1(n246), .A2(n247), .ZN(n8) );
  INV_X2 U254 ( .A(A[8]), .ZN(n247) );
  INV_X2 U255 ( .A(B[8]), .ZN(n246) );
  OAI21_X2 U256 ( .B1(n248), .B2(n195), .A(n202), .ZN(n6) );
  INV_X1 U257 ( .A(n249), .ZN(n202) );
  NAND2_X2 U258 ( .A1(n250), .A2(n251), .ZN(n249) );
  NAND4_X2 U259 ( .A1(n252), .A2(n21), .A3(n13), .A4(n15), .ZN(n251) );
  NAND2_X2 U260 ( .A1(n20), .A2(n25), .ZN(n252) );
  NAND2_X2 U261 ( .A1(B[4]), .A2(A[4]), .ZN(n25) );
  NAND2_X2 U262 ( .A1(B[5]), .A2(A[5]), .ZN(n20) );
  AOI21_X2 U263 ( .B1(n253), .B2(n15), .A(n254), .ZN(n250) );
  INV_X1 U264 ( .A(n16), .ZN(n254) );
  NAND2_X2 U265 ( .A1(B[7]), .A2(A[7]), .ZN(n16) );
  INV_X1 U266 ( .A(n12), .ZN(n253) );
  NAND2_X2 U267 ( .A1(B[6]), .A2(A[6]), .ZN(n12) );
  NAND4_X2 U268 ( .A1(n27), .A2(n21), .A3(n13), .A4(n15), .ZN(n195) );
  NAND2_X2 U269 ( .A1(n255), .A2(n256), .ZN(n15) );
  INV_X2 U270 ( .A(A[7]), .ZN(n256) );
  INV_X2 U271 ( .A(B[7]), .ZN(n255) );
  NAND2_X2 U272 ( .A1(n257), .A2(n258), .ZN(n13) );
  INV_X2 U273 ( .A(A[6]), .ZN(n258) );
  INV_X2 U274 ( .A(B[6]), .ZN(n257) );
  NAND2_X2 U275 ( .A1(n259), .A2(n260), .ZN(n21) );
  INV_X2 U276 ( .A(A[5]), .ZN(n260) );
  INV_X2 U277 ( .A(B[5]), .ZN(n259) );
  NAND2_X2 U278 ( .A1(n261), .A2(n262), .ZN(n27) );
  INV_X2 U279 ( .A(A[4]), .ZN(n262) );
  INV_X2 U280 ( .A(B[4]), .ZN(n261) );
  INV_X1 U281 ( .A(n26), .ZN(n248) );
  INV_X1 U282 ( .A(n58), .ZN(n32) );
  NOR2_X2 U283 ( .A1(n264), .A2(n265), .ZN(n201) );
  OAI21_X2 U284 ( .B1(n266), .B2(n33), .A(n36), .ZN(n265) );
  NAND2_X2 U285 ( .A1(B[3]), .A2(A[3]), .ZN(n36) );
  NAND2_X2 U286 ( .A1(B[2]), .A2(A[2]), .ZN(n33) );
  INV_X2 U287 ( .A(n35), .ZN(n266) );
  NOR2_X2 U288 ( .A1(n267), .A2(n268), .ZN(n264) );
  NAND2_X2 U289 ( .A1(n56), .A2(n269), .ZN(n268) );
  NAND2_X2 U290 ( .A1(n55), .A2(n163), .ZN(n269) );
  NAND2_X2 U291 ( .A1(B[1]), .A2(A[1]), .ZN(n55) );
  NAND2_X2 U292 ( .A1(n270), .A2(n271), .ZN(n56) );
  INV_X2 U293 ( .A(A[1]), .ZN(n271) );
  INV_X2 U294 ( .A(B[1]), .ZN(n270) );
  NAND2_X2 U295 ( .A1(n58), .A2(n35), .ZN(n267) );
  NAND2_X2 U296 ( .A1(n272), .A2(n273), .ZN(n35) );
  INV_X2 U297 ( .A(A[3]), .ZN(n273) );
  INV_X2 U298 ( .A(B[3]), .ZN(n272) );
  NAND2_X2 U299 ( .A1(n274), .A2(n275), .ZN(n58) );
  INV_X2 U300 ( .A(A[2]), .ZN(n275) );
  INV_X2 U301 ( .A(B[2]), .ZN(n274) );
  INV_X1 U302 ( .A(n3), .ZN(n234) );
  NAND2_X2 U303 ( .A1(n276), .A2(n277), .ZN(n3) );
  INV_X2 U304 ( .A(A[9]), .ZN(n277) );
  INV_X2 U305 ( .A(B[9]), .ZN(n276) );
  NAND2_X2 U306 ( .A1(n233), .A2(n230), .ZN(n243) );
  NAND2_X2 U307 ( .A1(n278), .A2(n279), .ZN(n230) );
  INV_X2 U308 ( .A(A[10]), .ZN(n279) );
  INV_X2 U309 ( .A(B[10]), .ZN(n278) );
  NAND2_X2 U310 ( .A1(B[10]), .A2(A[10]), .ZN(n233) );
  NAND2_X2 U311 ( .A1(n163), .A2(n263), .ZN(n280) );
  NAND2_X2 U312 ( .A1(n281), .A2(n282), .ZN(n263) );
  INV_X2 U313 ( .A(A[0]), .ZN(n282) );
  INV_X2 U314 ( .A(B[0]), .ZN(n281) );
  NAND2_X2 U315 ( .A1(B[0]), .A2(A[0]), .ZN(n163) );
endmodule


module ALU_DATA_W32 ( .FUNC({\FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), A, 
        B, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   N19, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N794, N795, N796, n121, n123, n124, n127, n130, n131, n136,
         n146, n148, n150, n151, n157, n159, n162, n163, n170, n172, n175,
         n176, n183, n184, n186, n192, n195, n196, n197, n198, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n213, n214, n217,
         n218, n219, n220, n232, n235, n239, n247, n253, n254, n258, n259,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n279,
         n285, n295, n302, n338, n339, n378, n401, n402, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n454, n455,
         n465, n474, n480, n482, n483, n484, n485, n487, n488, n489, n496,
         n497, n503, n504, n506, n507, n508, n509, n512, n513, n518, n519,
         n520, n521, n522, n523, n524, n527, n528, n529, n530, n534, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n547, n549,
         n550, n551, n552, n553, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n19, n20, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n122,
         n125, n126, n128, n129, n132, n133, n134, n135, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n147, n149, n152, n153, n154,
         n155, n156, n158, n160, n161, n164, n165, n166, n167, n168, n169,
         n171, n173, n174, n177, n178, n179, n180, n181, n182, n185, n187,
         n188, n189, n190, n191, n193, n194, n199, n200, n201, n212, n215,
         n216, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n233, n234, n236, n237, n238, n240, n241, n242, n243, n244,
         n245, n246, n248, n249, n250, n251, n252, n255, n256, n257, n260,
         n261, n262, n273, n274, n275, n276, n277, n278, n280, n281, n282,
         n283, n284, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n296, n297, n298, n299, n300, n301, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n403, n404, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n466, n467, n468, n469, n470,
         n471, n472, n473, n475, n476, n477, n478, n479, n481, n486, n490,
         n491, n492, n493, n494, n495, n498, n499, n500, n501, n502, n505,
         n510, n511, n514, n515, n516, n517, n525, n526, n531, n532, n533,
         n535, n546, n548, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748;
  wire   [3:0] FUNC;

  OAI21_X2 U17 ( .B1(B[9]), .B2(n57), .A(n53), .ZN(n121) );
  OAI221_X2 U19 ( .B1(A[9]), .B2(n58), .C1(n735), .C2(n49), .A(n52), .ZN(n127)
         );
  OAI21_X2 U24 ( .B1(B[8]), .B2(n57), .A(n52), .ZN(n146) );
  OAI221_X2 U26 ( .B1(A[8]), .B2(n58), .C1(n49), .C2(n736), .A(n52), .ZN(n148)
         );
  OAI21_X2 U31 ( .B1(B[7]), .B2(n57), .A(n52), .ZN(n157) );
  OAI221_X2 U33 ( .B1(A[7]), .B2(n58), .C1(n49), .C2(n737), .A(n52), .ZN(n159)
         );
  OAI21_X2 U38 ( .B1(B[6]), .B2(n57), .A(n52), .ZN(n170) );
  OAI221_X2 U40 ( .B1(A[6]), .B2(n58), .C1(n49), .C2(n738), .A(n52), .ZN(n172)
         );
  OAI21_X2 U45 ( .B1(B[5]), .B2(n57), .A(n52), .ZN(n183) );
  OAI221_X2 U47 ( .B1(A[5]), .B2(n58), .C1(n49), .C2(n739), .A(n52), .ZN(n184)
         );
  OAI21_X2 U52 ( .B1(B[4]), .B2(n57), .A(n53), .ZN(n192) );
  OAI221_X2 U54 ( .B1(A[4]), .B2(n58), .C1(n49), .C2(n740), .A(n52), .ZN(n195)
         );
  AOI221_X2 U60 ( .B1(A[3]), .B2(n51), .C1(n62), .C2(n741), .A(n56), .ZN(n202)
         );
  AOI22_X2 U61 ( .A1(n703), .A2(n723), .B1(A[3]), .B2(n203), .ZN(n198) );
  OAI21_X2 U62 ( .B1(B[3]), .B2(n57), .A(n53), .ZN(n203) );
  AOI22_X2 U63 ( .A1(n205), .A2(n206), .B1(n207), .B2(n208), .ZN(n204) );
  OAI221_X2 U64 ( .B1(n209), .B2(n730), .C1(n208), .C2(n206), .A(n210), .ZN(
        n197) );
  AOI22_X2 U65 ( .A1(n163), .A2(n701), .B1(n162), .B2(n213), .ZN(n211) );
  OAI221_X2 U66 ( .B1(n48), .B2(n734), .C1(n735), .C2(n40), .A(n214), .ZN(n163) );
  AOI22_X2 U67 ( .A1(A[8]), .A2(n24), .B1(A[7]), .B2(n30), .ZN(n214) );
  OAI22_X2 U68 ( .A1(n726), .A2(n744), .B1(n217), .B2(n10), .ZN(n209) );
  AOI221_X2 U69 ( .B1(A[6]), .B2(n46), .C1(A[5]), .C2(n36), .A(n220), .ZN(n217) );
  OAI22_X2 U70 ( .A1(n28), .A2(n741), .B1(n20), .B2(n740), .ZN(n220) );
  OAI22_X2 U77 ( .A1(n20), .A2(n706), .B1(n707), .B2(n40), .ZN(n235) );
  AOI211_X2 U87 ( .C1(A[27]), .C2(n45), .A(n253), .B(n254), .ZN(n247) );
  OAI22_X2 U88 ( .A1(n20), .A2(n707), .B1(n708), .B2(n40), .ZN(n253) );
  AOI221_X2 U95 ( .B1(A[2]), .B2(n51), .C1(n62), .C2(n742), .A(n56), .ZN(n263)
         );
  AOI22_X2 U96 ( .A1(n703), .A2(n724), .B1(A[2]), .B2(n264), .ZN(n259) );
  OAI21_X2 U97 ( .B1(B[2]), .B2(n57), .A(n53), .ZN(n264) );
  AOI22_X2 U98 ( .A1(n266), .A2(n206), .B1(n267), .B2(n208), .ZN(n265) );
  OAI221_X2 U99 ( .B1(n268), .B2(n731), .C1(n208), .C2(n206), .A(n210), .ZN(
        n258) );
  AOI22_X2 U100 ( .A1(n176), .A2(n701), .B1(n175), .B2(n213), .ZN(n269) );
  OAI221_X2 U101 ( .B1(n735), .B2(n48), .C1(n41), .C2(n736), .A(n270), .ZN(
        n176) );
  AOI22_X2 U102 ( .A1(A[7]), .A2(n24), .B1(A[6]), .B2(n30), .ZN(n270) );
  OAI22_X2 U103 ( .A1(n727), .A2(n744), .B1(n271), .B2(n10), .ZN(n268) );
  AOI221_X2 U104 ( .B1(A[5]), .B2(n46), .C1(A[4]), .C2(n36), .A(n272), .ZN(
        n271) );
  OAI22_X2 U105 ( .A1(n28), .A2(n742), .B1(n20), .B2(n741), .ZN(n272) );
  AOI221_X2 U112 ( .B1(A[26]), .B2(n46), .C1(A[27]), .C2(n36), .A(n285), .ZN(
        n279) );
  OAI22_X2 U113 ( .A1(n28), .A2(n707), .B1(n20), .B2(n708), .ZN(n285) );
  AOI221_X2 U124 ( .B1(A[25]), .B2(n45), .C1(A[26]), .C2(n36), .A(n302), .ZN(
        n295) );
  OAI22_X2 U125 ( .A1(n28), .A2(n708), .B1(n20), .B2(n709), .ZN(n302) );
  AOI221_X2 U227 ( .B1(A[1]), .B2(n51), .C1(n61), .C2(n743), .A(n56), .ZN(n405) );
  AOI22_X2 U228 ( .A1(n703), .A2(n725), .B1(A[1]), .B2(n406), .ZN(n402) );
  OAI21_X2 U229 ( .B1(B[1]), .B2(n57), .A(n53), .ZN(n406) );
  AOI22_X2 U230 ( .A1(n408), .A2(n206), .B1(n409), .B2(n208), .ZN(n407) );
  OAI221_X2 U231 ( .B1(n410), .B2(n732), .C1(n208), .C2(n206), .A(n210), .ZN(
        n401) );
  NOR2_X2 U232 ( .A1(n411), .A2(N19), .ZN(n206) );
  NOR2_X2 U233 ( .A1(n239), .A2(N19), .ZN(n208) );
  AOI22_X2 U234 ( .A1(n186), .A2(n701), .B1(n136), .B2(n213), .ZN(n412) );
  OAI221_X2 U235 ( .B1(n20), .B2(n734), .C1(n735), .C2(n28), .A(n413), .ZN(
        n136) );
  AOI22_X2 U236 ( .A1(A[12]), .A2(n43), .B1(A[11]), .B2(n37), .ZN(n413) );
  OAI221_X2 U237 ( .B1(n20), .B2(n738), .C1(n28), .C2(n739), .A(n414), .ZN(
        n186) );
  AOI22_X2 U238 ( .A1(A[8]), .A2(n43), .B1(A[7]), .B2(n36), .ZN(n414) );
  OAI22_X2 U239 ( .A1(n728), .A2(n744), .B1(n415), .B2(n10), .ZN(n410) );
  AOI221_X2 U240 ( .B1(A[4]), .B2(n45), .C1(A[3]), .C2(n36), .A(n416), .ZN(
        n415) );
  OAI22_X2 U241 ( .A1(n28), .A2(n743), .B1(n20), .B2(n742), .ZN(n416) );
  NAND2_X2 U249 ( .A1(n232), .A2(A[31]), .ZN(n378) );
  AOI22_X2 U292 ( .A1(A[13]), .A2(n43), .B1(A[14]), .B2(n36), .ZN(n454) );
  AOI22_X2 U305 ( .A1(A[12]), .A2(n43), .B1(A[13]), .B2(n36), .ZN(n465) );
  AOI22_X2 U318 ( .A1(A[11]), .A2(n43), .B1(A[12]), .B2(n36), .ZN(n474) );
  AOI21_X2 U326 ( .B1(A[31]), .B2(B[1]), .A(n480), .ZN(n338) );
  AOI22_X2 U329 ( .A1(A[28]), .A2(n43), .B1(A[27]), .B2(n36), .ZN(n482) );
  AOI22_X2 U332 ( .A1(A[20]), .A2(n43), .B1(A[19]), .B2(n36), .ZN(n483) );
  AOI22_X2 U334 ( .A1(A[24]), .A2(n43), .B1(A[23]), .B2(n36), .ZN(n484) );
  AOI22_X2 U336 ( .A1(A[16]), .A2(n43), .B1(A[15]), .B2(n37), .ZN(n485) );
  AOI22_X2 U341 ( .A1(A[2]), .A2(n43), .B1(A[3]), .B2(n37), .ZN(n487) );
  AOI22_X2 U344 ( .A1(A[10]), .A2(n44), .B1(A[11]), .B2(n38), .ZN(n488) );
  AOI22_X2 U346 ( .A1(A[6]), .A2(n43), .B1(A[7]), .B2(n37), .ZN(n489) );
  AOI22_X2 U359 ( .A1(A[1]), .A2(n44), .B1(A[2]), .B2(n37), .ZN(n496) );
  AOI22_X2 U361 ( .A1(A[5]), .A2(n45), .B1(A[6]), .B2(n37), .ZN(n497) );
  OAI21_X2 U369 ( .B1(B[11]), .B2(n57), .A(n53), .ZN(n503) );
  OAI221_X2 U371 ( .B1(A[11]), .B2(n58), .C1(n49), .C2(n733), .A(n52), .ZN(
        n504) );
  AOI22_X2 U377 ( .A1(A[26]), .A2(n45), .B1(A[25]), .B2(n37), .ZN(n506) );
  AOI22_X2 U380 ( .A1(A[18]), .A2(n45), .B1(A[17]), .B2(n37), .ZN(n507) );
  AOI22_X2 U382 ( .A1(A[22]), .A2(n45), .B1(A[21]), .B2(n37), .ZN(n508) );
  OAI221_X2 U383 ( .B1(n20), .B2(n710), .C1(n28), .C2(n733), .A(n509), .ZN(
        n162) );
  AOI22_X2 U384 ( .A1(A[14]), .A2(n45), .B1(A[13]), .B2(n37), .ZN(n509) );
  AOI22_X2 U390 ( .A1(A[0]), .A2(n45), .B1(A[1]), .B2(n37), .ZN(n512) );
  AOI22_X2 U392 ( .A1(A[4]), .A2(n43), .B1(A[5]), .B2(n37), .ZN(n513) );
  OAI21_X2 U395 ( .B1(B[10]), .B2(n57), .A(n53), .ZN(n518) );
  NAND2_X2 U397 ( .A1(B[3]), .A2(A[31]), .ZN(n339) );
  AOI22_X2 U402 ( .A1(A[25]), .A2(n45), .B1(A[24]), .B2(n38), .ZN(n520) );
  OAI221_X2 U404 ( .B1(A[10]), .B2(n58), .C1(n49), .C2(n734), .A(n52), .ZN(
        n519) );
  AOI22_X2 U406 ( .A1(A[21]), .A2(n44), .B1(A[20]), .B2(n38), .ZN(n521) );
  OAI221_X2 U409 ( .B1(n20), .B2(n733), .C1(n28), .C2(n734), .A(n522), .ZN(
        n175) );
  AOI22_X2 U410 ( .A1(A[13]), .A2(n45), .B1(A[12]), .B2(n38), .ZN(n522) );
  AOI22_X2 U413 ( .A1(A[17]), .A2(n44), .B1(A[16]), .B2(n38), .ZN(n523) );
  NOR2_X2 U421 ( .A1(n411), .A2(n210), .ZN(n131) );
  AOI22_X2 U425 ( .A1(A[7]), .A2(n44), .B1(A[8]), .B2(n38), .ZN(n527) );
  AOI22_X2 U428 ( .A1(A[3]), .A2(n44), .B1(A[4]), .B2(n38), .ZN(n528) );
  AOI22_X2 U433 ( .A1(n61), .A2(n713), .B1(n51), .B2(B[0]), .ZN(n534) );
  AOI22_X2 U439 ( .A1(n536), .A2(n537), .B1(B[0]), .B2(n538), .ZN(n530) );
  OAI21_X2 U440 ( .B1(A[0]), .B2(n57), .A(n53), .ZN(n538) );
  OAI22_X2 U441 ( .A1(n455), .A2(n210), .B1(n703), .B2(n539), .ZN(n537) );
  AOI221_X2 U442 ( .B1(n213), .B2(n151), .C1(n701), .C2(n196), .A(n540), .ZN(
        n539) );
  OAI22_X2 U443 ( .A1(n729), .A2(n744), .B1(n541), .B2(n10), .ZN(n540) );
  AOI211_X2 U444 ( .C1(A[3]), .C2(n45), .A(n542), .B(n702), .ZN(n541) );
  OAI22_X2 U446 ( .A1(n22), .A2(n743), .B1(n41), .B2(n742), .ZN(n542) );
  AOI22_X2 U448 ( .A1(A[15]), .A2(n44), .B1(A[14]), .B2(n38), .ZN(n543) );
  OAI221_X2 U449 ( .B1(n20), .B2(n739), .C1(n28), .C2(n740), .A(n544), .ZN(
        n196) );
  AOI22_X2 U450 ( .A1(A[7]), .A2(n44), .B1(A[6]), .B2(n38), .ZN(n544) );
  OAI221_X2 U451 ( .B1(n735), .B2(n22), .C1(n28), .C2(n736), .A(n545), .ZN(
        n151) );
  AOI22_X2 U452 ( .A1(A[11]), .A2(n44), .B1(A[10]), .B2(n38), .ZN(n545) );
  NAND2_X2 U453 ( .A1(B[4]), .A2(n714), .ZN(n210) );
  AOI22_X2 U457 ( .A1(A[27]), .A2(n44), .B1(A[26]), .B2(n38), .ZN(n547) );
  NOR2_X2 U458 ( .A1(n711), .A2(B[2]), .ZN(n213) );
  NOR2_X2 U461 ( .A1(n712), .A2(n711), .ZN(n232) );
  AOI22_X2 U464 ( .A1(A[19]), .A2(n44), .B1(A[18]), .B2(n38), .ZN(n549) );
  AOI22_X2 U467 ( .A1(A[23]), .A2(n44), .B1(A[22]), .B2(n39), .ZN(n550) );
  NOR2_X2 U468 ( .A1(n746), .A2(B[0]), .ZN(n219) );
  NOR2_X2 U469 ( .A1(n713), .A2(n746), .ZN(n218) );
  NOR2_X2 U472 ( .A1(N19), .A2(n524), .ZN(n536) );
  AND2_X2 U473 ( .A1(n411), .A2(n239), .ZN(n524) );
  OAI21_X2 U477 ( .B1(FUNC[1]), .B2(n552), .A(n553), .ZN(n551) );
  AOI22_X2 U478 ( .A1(N794), .A2(n705), .B1(N795), .B2(FUNC[0]), .ZN(n552) );
  NAND3_X1 U577 ( .A1(n551), .A2(n704), .A3(FUNC[3]), .ZN(n529) );
  NAND3_X1 U578 ( .A1(FUNC[1]), .A2(n705), .A3(N796), .ZN(n553) );
  ALU_DATA_W32_DW01_cmp6_0 r80 ( .A(B), .B(A), .TC(1'b0), .LE(N794), .GE(N795), 
        .NE(N796) );
  ALU_DATA_W32_DW01_sub_2 sub_128 ( .A(A), .B(B), .CI(1'b0), .DIFF({N122, N121, 
        N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91}) );
  ALU_DATA_W32_DW01_add_2 add_125 ( .A(A), .B(B), .CI(1'b0), .SUM({N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, 
        N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60, N59}) );
  INV_X2 U3 ( .A(n12), .ZN(n10) );
  INV_X2 U4 ( .A(n12), .ZN(n11) );
  INV_X2 U6 ( .A(n25), .ZN(n20) );
  INV_X2 U7 ( .A(n24), .ZN(n22) );
  INV_X2 U8 ( .A(n30), .ZN(n28) );
  INV_X2 U9 ( .A(n30), .ZN(n29) );
  INV_X2 U10 ( .A(n42), .ZN(n36) );
  INV_X2 U12 ( .A(n42), .ZN(n37) );
  INV_X2 U13 ( .A(n41), .ZN(n38) );
  INV_X2 U15 ( .A(n41), .ZN(n39) );
  INV_X2 U16 ( .A(n48), .ZN(n45) );
  INV_X2 U18 ( .A(n48), .ZN(n46) );
  INV_X2 U20 ( .A(n64), .ZN(n57) );
  INV_X2 U21 ( .A(n63), .ZN(n58) );
  INV_X2 U22 ( .A(n63), .ZN(n59) );
  INV_X2 U23 ( .A(n185), .ZN(n308) );
  INV_X2 U25 ( .A(n229), .ZN(n241) );
  INV_X2 U27 ( .A(n99), .ZN(n310) );
  INV_X2 U28 ( .A(n305), .ZN(n212) );
  INV_X2 U29 ( .A(n281), .ZN(n595) );
  INV_X2 U30 ( .A(n331), .ZN(n596) );
  INV_X2 U32 ( .A(n248), .ZN(n598) );
  INV_X2 U34 ( .A(n348), .ZN(n641) );
  INV_X2 U35 ( .A(n351), .ZN(n637) );
  CLKBUF_X3 U36 ( .A(n594), .Z(n1) );
  CLKBUF_X3 U37 ( .A(n594), .Z(n2) );
  CLKBUF_X3 U39 ( .A(n594), .Z(n3) );
  CLKBUF_X3 U41 ( .A(n693), .Z(n4) );
  CLKBUF_X3 U42 ( .A(n693), .Z(n5) );
  CLKBUF_X3 U43 ( .A(n693), .Z(n6) );
  CLKBUF_X3 U44 ( .A(n695), .Z(n7) );
  CLKBUF_X3 U46 ( .A(n695), .Z(n8) );
  CLKBUF_X3 U48 ( .A(n695), .Z(n9) );
  INV_X1 U49 ( .A(n745), .ZN(n12) );
  INV_X1 U50 ( .A(n745), .ZN(n13) );
  INV_X1 U51 ( .A(n745), .ZN(n14) );
  INV_X1 U53 ( .A(n745), .ZN(n15) );
  INV_X1 U55 ( .A(n745), .ZN(n16) );
  CLKBUF_X3 U56 ( .A(n747), .Z(n19) );
  INV_X1 U57 ( .A(n24), .ZN(n23) );
  INV_X2 U58 ( .A(n19), .ZN(n24) );
  INV_X2 U59 ( .A(n19), .ZN(n25) );
  INV_X2 U71 ( .A(n19), .ZN(n26) );
  INV_X2 U72 ( .A(n19), .ZN(n27) );
  CLKBUF_X3 U73 ( .A(n35), .Z(n30) );
  CLKBUF_X3 U74 ( .A(n35), .Z(n31) );
  CLKBUF_X3 U75 ( .A(n34), .Z(n32) );
  CLKBUF_X3 U76 ( .A(n34), .Z(n33) );
  INV_X2 U78 ( .A(n748), .ZN(n34) );
  INV_X2 U79 ( .A(n748), .ZN(n35) );
  INV_X2 U80 ( .A(n219), .ZN(n40) );
  INV_X2 U81 ( .A(n219), .ZN(n41) );
  INV_X2 U82 ( .A(n219), .ZN(n42) );
  INV_X1 U83 ( .A(n48), .ZN(n43) );
  INV_X1 U84 ( .A(n48), .ZN(n44) );
  INV_X1 U85 ( .A(n48), .ZN(n47) );
  INV_X4 U86 ( .A(n218), .ZN(n48) );
  INV_X1 U89 ( .A(n51), .ZN(n49) );
  INV_X1 U90 ( .A(n51), .ZN(n50) );
  INV_X8 U91 ( .A(n130), .ZN(n51) );
  INV_X1 U92 ( .A(n56), .ZN(n52) );
  INV_X1 U93 ( .A(n56), .ZN(n53) );
  INV_X1 U94 ( .A(n56), .ZN(n54) );
  INV_X1 U106 ( .A(n56), .ZN(n55) );
  INV_X8 U107 ( .A(n124), .ZN(n56) );
  INV_X1 U108 ( .A(n63), .ZN(n60) );
  INV_X1 U109 ( .A(n123), .ZN(n61) );
  INV_X1 U110 ( .A(n123), .ZN(n62) );
  INV_X1 U111 ( .A(n123), .ZN(n63) );
  INV_X1 U114 ( .A(n123), .ZN(n64) );
  INV_X1 U115 ( .A(n123), .ZN(n65) );
  INV_X1 U116 ( .A(B[1]), .ZN(n66) );
  NAND2_X1 U117 ( .A1(B[0]), .A2(n66), .ZN(n747) );
  INV_X1 U118 ( .A(B[0]), .ZN(n713) );
  NAND2_X1 U119 ( .A1(n66), .A2(n713), .ZN(n748) );
  NAND2_X1 U120 ( .A1(A[13]), .A2(n25), .ZN(n286) );
  NAND2_X1 U121 ( .A1(n33), .A2(A[12]), .ZN(n216) );
  NAND3_X1 U122 ( .A1(n543), .A2(n286), .A3(n216), .ZN(n150) );
  INV_X1 U123 ( .A(FUNC[2]), .ZN(n704) );
  NAND2_X1 U126 ( .A1(FUNC[0]), .A2(n704), .ZN(n67) );
  INV_X1 U127 ( .A(n67), .ZN(n77) );
  INV_X1 U128 ( .A(FUNC[3]), .ZN(n74) );
  NAND2_X1 U129 ( .A1(FUNC[1]), .A2(n74), .ZN(n68) );
  INV_X1 U130 ( .A(n68), .ZN(n344) );
  NAND2_X1 U131 ( .A1(n77), .A2(n344), .ZN(n124) );
  NAND2_X1 U132 ( .A1(FUNC[2]), .A2(FUNC[0]), .ZN(n69) );
  INV_X1 U133 ( .A(n69), .ZN(n79) );
  NAND2_X1 U134 ( .A1(n79), .A2(n344), .ZN(n239) );
  INV_X1 U135 ( .A(B[3]), .ZN(n711) );
  INV_X1 U136 ( .A(B[2]), .ZN(n712) );
  NAND2_X1 U137 ( .A1(n711), .A2(n712), .ZN(n745) );
  NAND2_X1 U138 ( .A1(n534), .A2(n55), .ZN(n71) );
  INV_X1 U139 ( .A(n239), .ZN(n349) );
  NAND3_X1 U140 ( .A1(A[31]), .A2(N19), .A3(n349), .ZN(n178) );
  NAND2_X1 U141 ( .A1(n530), .A2(n178), .ZN(n70) );
  AOI21_X1 U142 ( .B1(A[0]), .B2(n71), .A(n70), .ZN(n82) );
  INV_X1 U143 ( .A(FUNC[0]), .ZN(n705) );
  NAND2_X1 U144 ( .A1(n704), .A2(n705), .ZN(n72) );
  INV_X1 U145 ( .A(n72), .ZN(n199) );
  INV_X1 U146 ( .A(FUNC[1]), .ZN(n73) );
  NAND2_X1 U147 ( .A1(n74), .A2(n73), .ZN(n75) );
  INV_X1 U148 ( .A(n75), .ZN(n194) );
  NAND2_X1 U149 ( .A1(n199), .A2(n194), .ZN(n76) );
  INV_X1 U150 ( .A(n76), .ZN(n695) );
  NAND2_X1 U151 ( .A1(n77), .A2(n194), .ZN(n78) );
  INV_X1 U152 ( .A(n78), .ZN(n693) );
  NAND2_X1 U153 ( .A1(A[0]), .A2(n33), .ZN(n491) );
  INV_X1 U154 ( .A(n491), .ZN(n702) );
  INV_X1 U155 ( .A(N19), .ZN(n714) );
  NAND2_X1 U156 ( .A1(n210), .A2(n714), .ZN(n296) );
  INV_X1 U157 ( .A(n296), .ZN(n350) );
  NAND2_X1 U158 ( .A1(n79), .A2(n194), .ZN(n80) );
  INV_X1 U159 ( .A(n80), .ZN(n606) );
  NAND2_X1 U160 ( .A1(n350), .A2(n606), .ZN(n95) );
  INV_X1 U161 ( .A(n95), .ZN(n246) );
  NAND2_X1 U162 ( .A1(n246), .A2(n12), .ZN(n330) );
  INV_X1 U163 ( .A(n330), .ZN(n594) );
  AOI222_X1 U164 ( .A1(N59), .A2(n7), .B1(N91), .B2(n5), .C1(n702), .C2(n2), 
        .ZN(n81) );
  NAND3_X1 U165 ( .A1(n82), .A2(n81), .A3(n529), .ZN(RES[0]) );
  AOI22_X1 U166 ( .A1(N92), .A2(n5), .B1(N60), .B2(n8), .ZN(n85) );
  INV_X1 U167 ( .A(A[1]), .ZN(n86) );
  INV_X1 U168 ( .A(A[0]), .ZN(n87) );
  OAI22_X1 U169 ( .A1(n28), .A2(n86), .B1(n22), .B2(n87), .ZN(n625) );
  NAND2_X1 U170 ( .A1(n401), .A2(n402), .ZN(n83) );
  INV_X1 U171 ( .A(n178), .ZN(n153) );
  AOI211_X1 U172 ( .C1(n1), .C2(n625), .A(n83), .B(n153), .ZN(n84) );
  OAI211_X1 U173 ( .C1(n405), .C2(n746), .A(n85), .B(n84), .ZN(RES[1]) );
  AOI22_X1 U174 ( .A1(N93), .A2(n4), .B1(N61), .B2(n9), .ZN(n90) );
  INV_X1 U175 ( .A(A[2]), .ZN(n742) );
  OAI222_X1 U176 ( .A1(n742), .A2(n29), .B1(n42), .B2(n87), .C1(n22), .C2(n86), 
        .ZN(n649) );
  NAND2_X1 U177 ( .A1(n258), .A2(n259), .ZN(n88) );
  AOI211_X1 U178 ( .C1(n1), .C2(n649), .A(n88), .B(n153), .ZN(n89) );
  OAI211_X1 U179 ( .C1(n263), .C2(n712), .A(n90), .B(n89), .ZN(RES[2]) );
  AOI22_X1 U180 ( .A1(N94), .A2(n4), .B1(N62), .B2(n9), .ZN(n93) );
  INV_X1 U181 ( .A(A[3]), .ZN(n741) );
  OAI221_X1 U182 ( .B1(n742), .B2(n22), .C1(n741), .C2(n29), .A(n512), .ZN(
        n674) );
  NAND2_X1 U183 ( .A1(n197), .A2(n198), .ZN(n91) );
  AOI211_X1 U184 ( .C1(n1), .C2(n674), .A(n91), .B(n153), .ZN(n92) );
  OAI211_X1 U185 ( .C1(n202), .C2(n711), .A(n93), .B(n92), .ZN(RES[3]) );
  INV_X1 U186 ( .A(A[29]), .ZN(n707) );
  INV_X1 U187 ( .A(A[28]), .ZN(n708) );
  AOI22_X1 U188 ( .A1(A[30]), .A2(n39), .B1(A[31]), .B2(n47), .ZN(n94) );
  OAI221_X1 U189 ( .B1(n707), .B2(n22), .C1(n708), .C2(n29), .A(n94), .ZN(n227) );
  INV_X1 U190 ( .A(n227), .ZN(n327) );
  INV_X1 U191 ( .A(n213), .ZN(n579) );
  NAND2_X1 U192 ( .A1(A[21]), .A2(n27), .ZN(n450) );
  NAND2_X1 U193 ( .A1(A[20]), .A2(n32), .ZN(n417) );
  NAND3_X1 U194 ( .A1(n550), .A2(n450), .A3(n417), .ZN(n324) );
  INV_X1 U195 ( .A(n324), .ZN(n140) );
  NAND2_X1 U196 ( .A1(A[25]), .A2(n27), .ZN(n567) );
  NAND2_X1 U197 ( .A1(A[24]), .A2(n32), .ZN(n498) );
  NAND3_X1 U198 ( .A1(n547), .A2(n567), .A3(n498), .ZN(n200) );
  INV_X1 U199 ( .A(n200), .ZN(n326) );
  NAND2_X1 U200 ( .A1(B[2]), .A2(n711), .ZN(n684) );
  OAI222_X1 U201 ( .A1(n327), .A2(n579), .B1(n11), .B2(n140), .C1(n326), .C2(
        n684), .ZN(n422) );
  NOR2_X1 U202 ( .A1(B[3]), .A2(n95), .ZN(n96) );
  INV_X1 U203 ( .A(A[4]), .ZN(n740) );
  OAI221_X1 U204 ( .B1(n741), .B2(n22), .C1(n740), .C2(n29), .A(n496), .ZN(
        n320) );
  INV_X1 U205 ( .A(n320), .ZN(n492) );
  MUX2_X1 U206 ( .A(n492), .B(n491), .S(B[2]), .Z(n608) );
  INV_X1 U207 ( .A(n608), .ZN(n399) );
  AOI221_X1 U208 ( .B1(n131), .B2(n422), .C1(n96), .C2(n399), .A(n153), .ZN(
        n104) );
  INV_X1 U209 ( .A(n524), .ZN(n97) );
  NAND2_X1 U210 ( .A1(n350), .A2(n97), .ZN(n329) );
  INV_X1 U211 ( .A(n329), .ZN(n100) );
  INV_X1 U212 ( .A(n684), .ZN(n701) );
  NAND2_X1 U213 ( .A1(n100), .A2(n701), .ZN(n185) );
  INV_X1 U214 ( .A(n210), .ZN(n703) );
  NAND2_X1 U215 ( .A1(n349), .A2(n703), .ZN(n229) );
  INV_X1 U216 ( .A(n422), .ZN(n98) );
  NAND2_X1 U217 ( .A1(n98), .A2(n378), .ZN(n424) );
  NAND2_X1 U218 ( .A1(n100), .A2(n232), .ZN(n306) );
  INV_X1 U219 ( .A(n306), .ZN(n201) );
  NAND2_X1 U220 ( .A1(A[17]), .A2(n27), .ZN(n370) );
  NAND2_X1 U221 ( .A1(A[16]), .A2(n32), .ZN(n321) );
  NAND3_X1 U222 ( .A1(n549), .A2(n370), .A3(n321), .ZN(n323) );
  AOI222_X1 U223 ( .A1(n151), .A2(n308), .B1(n241), .B2(n424), .C1(n201), .C2(
        n323), .ZN(n103) );
  NAND2_X1 U224 ( .A1(n100), .A2(n213), .ZN(n99) );
  NAND2_X1 U225 ( .A1(n100), .A2(n15), .ZN(n305) );
  AOI222_X1 U226 ( .A1(N95), .A2(n4), .B1(n310), .B2(n150), .C1(n196), .C2(
        n212), .ZN(n102) );
  AOI222_X1 U242 ( .A1(n192), .A2(A[4]), .B1(N63), .B2(n9), .C1(B[4]), .C2(
        n195), .ZN(n101) );
  NAND4_X1 U243 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .ZN(RES[4]) );
  INV_X1 U244 ( .A(A[30]), .ZN(n706) );
  OAI22_X1 U245 ( .A1(n707), .A2(n29), .B1(n706), .B2(n22), .ZN(n480) );
  NAND2_X1 U246 ( .A1(A[22]), .A2(n27), .ZN(n471) );
  NAND2_X1 U247 ( .A1(A[21]), .A2(n32), .ZN(n434) );
  NAND3_X1 U248 ( .A1(n484), .A2(n471), .A3(n434), .ZN(n257) );
  INV_X1 U250 ( .A(n257), .ZN(n337) );
  NAND2_X1 U251 ( .A1(A[26]), .A2(n27), .ZN(n588) );
  NAND2_X1 U252 ( .A1(A[25]), .A2(n32), .ZN(n533) );
  NAND3_X1 U253 ( .A1(n482), .A2(n588), .A3(n533), .ZN(n149) );
  INV_X1 U254 ( .A(n149), .ZN(n341) );
  OAI22_X1 U255 ( .A1(n10), .A2(n337), .B1(n341), .B2(n684), .ZN(n105) );
  INV_X1 U256 ( .A(n105), .ZN(n108) );
  OAI211_X1 U257 ( .C1(n338), .C2(n579), .A(n108), .B(n378), .ZN(n439) );
  NAND2_X1 U258 ( .A1(A[18]), .A2(n26), .ZN(n389) );
  NAND2_X1 U259 ( .A1(A[17]), .A2(n32), .ZN(n357) );
  NAND3_X1 U260 ( .A1(n483), .A2(n389), .A3(n357), .ZN(n336) );
  INV_X1 U261 ( .A(n625), .ZN(n154) );
  NAND2_X1 U262 ( .A1(n246), .A2(n701), .ZN(n331) );
  OAI21_X1 U263 ( .B1(n154), .B2(n331), .A(n178), .ZN(n106) );
  AOI221_X1 U264 ( .B1(n241), .B2(n439), .C1(n201), .C2(n336), .A(n106), .ZN(
        n112) );
  INV_X1 U265 ( .A(A[5]), .ZN(n739) );
  OAI221_X1 U266 ( .B1(n740), .B2(n22), .C1(n739), .C2(n29), .A(n487), .ZN(
        n626) );
  NAND2_X1 U267 ( .A1(A[14]), .A2(n26), .ZN(n304) );
  NAND2_X1 U268 ( .A1(A[13]), .A2(n32), .ZN(n252) );
  NAND3_X1 U269 ( .A1(n485), .A2(n304), .A3(n252), .ZN(n255) );
  INV_X1 U270 ( .A(A[31]), .ZN(n117) );
  INV_X1 U271 ( .A(n480), .ZN(n107) );
  OAI21_X1 U272 ( .B1(n42), .B2(n117), .A(n107), .ZN(n243) );
  INV_X1 U273 ( .A(n243), .ZN(n644) );
  OAI21_X1 U274 ( .B1(n644), .B2(n579), .A(n108), .ZN(n440) );
  AOI222_X1 U275 ( .A1(n1), .A2(n626), .B1(n310), .B2(n255), .C1(n131), .C2(
        n440), .ZN(n111) );
  AOI222_X1 U276 ( .A1(N96), .A2(n4), .B1(n136), .B2(n308), .C1(n186), .C2(
        n212), .ZN(n110) );
  AOI222_X1 U277 ( .A1(n183), .A2(A[5]), .B1(N64), .B2(n9), .C1(B[5]), .C2(
        n184), .ZN(n109) );
  NAND4_X1 U278 ( .A1(n112), .A2(n111), .A3(n110), .A4(n109), .ZN(RES[5]) );
  NAND2_X1 U279 ( .A1(n33), .A2(A[30]), .ZN(n700) );
  OAI21_X1 U280 ( .B1(n33), .B2(n117), .A(n700), .ZN(n113) );
  INV_X1 U281 ( .A(n113), .ZN(n663) );
  NAND2_X1 U282 ( .A1(A[23]), .A2(n26), .ZN(n499) );
  NAND2_X1 U283 ( .A1(A[22]), .A2(n31), .ZN(n451) );
  NAND3_X1 U284 ( .A1(n520), .A2(n499), .A3(n451), .ZN(n288) );
  INV_X1 U285 ( .A(n288), .ZN(n363) );
  INV_X1 U286 ( .A(A[27]), .ZN(n709) );
  NAND2_X1 U287 ( .A1(A[26]), .A2(n31), .ZN(n568) );
  AOI22_X1 U288 ( .A1(A[28]), .A2(n39), .B1(A[29]), .B2(n47), .ZN(n114) );
  OAI211_X1 U289 ( .C1(n709), .C2(n22), .A(n568), .B(n114), .ZN(n161) );
  INV_X1 U290 ( .A(n161), .ZN(n365) );
  OAI22_X1 U291 ( .A1(n10), .A2(n363), .B1(n365), .B2(n684), .ZN(n115) );
  INV_X1 U293 ( .A(n115), .ZN(n118) );
  OAI211_X1 U294 ( .C1(n663), .C2(n579), .A(n378), .B(n118), .ZN(n458) );
  NAND2_X1 U295 ( .A1(A[19]), .A2(n26), .ZN(n418) );
  NAND2_X1 U296 ( .A1(A[18]), .A2(n31), .ZN(n371) );
  NAND3_X1 U297 ( .A1(n521), .A2(n418), .A3(n371), .ZN(n362) );
  INV_X1 U298 ( .A(n649), .ZN(n561) );
  OAI21_X1 U299 ( .B1(n561), .B2(n331), .A(n178), .ZN(n116) );
  AOI221_X1 U300 ( .B1(n241), .B2(n458), .C1(n201), .C2(n362), .A(n116), .ZN(
        n125) );
  INV_X1 U301 ( .A(A[6]), .ZN(n738) );
  OAI221_X1 U302 ( .B1(n739), .B2(n22), .C1(n738), .C2(n29), .A(n528), .ZN(
        n650) );
  NAND2_X1 U303 ( .A1(A[15]), .A2(n25), .ZN(n322) );
  NAND2_X1 U304 ( .A1(A[14]), .A2(n31), .ZN(n284) );
  NAND3_X1 U306 ( .A1(n523), .A2(n322), .A3(n284), .ZN(n167) );
  OAI21_X1 U307 ( .B1(n22), .B2(n117), .A(n700), .ZN(n277) );
  INV_X1 U308 ( .A(n277), .ZN(n669) );
  OAI21_X1 U309 ( .B1(n669), .B2(n579), .A(n118), .ZN(n457) );
  AOI222_X1 U310 ( .A1(n1), .A2(n650), .B1(n310), .B2(n167), .C1(n131), .C2(
        n457), .ZN(n122) );
  AOI222_X1 U311 ( .A1(N97), .A2(n4), .B1(n175), .B2(n308), .C1(n176), .C2(
        n212), .ZN(n120) );
  AOI222_X1 U312 ( .A1(n170), .A2(A[6]), .B1(N65), .B2(n9), .C1(B[6]), .C2(
        n172), .ZN(n119) );
  NAND4_X1 U313 ( .A1(n125), .A2(n122), .A3(n120), .A4(n119), .ZN(RES[6]) );
  NAND2_X1 U314 ( .A1(A[24]), .A2(n26), .ZN(n535) );
  NAND2_X1 U315 ( .A1(A[23]), .A2(n31), .ZN(n472) );
  NAND3_X1 U316 ( .A1(n506), .A2(n535), .A3(n472), .ZN(n309) );
  INV_X1 U317 ( .A(n309), .ZN(n382) );
  NAND2_X1 U319 ( .A1(n33), .A2(A[27]), .ZN(n589) );
  AOI22_X1 U320 ( .A1(A[29]), .A2(n39), .B1(A[30]), .B2(n46), .ZN(n126) );
  OAI211_X1 U321 ( .C1(n708), .C2(n23), .A(n589), .B(n126), .ZN(n177) );
  INV_X1 U322 ( .A(n177), .ZN(n384) );
  OAI22_X1 U323 ( .A1(n10), .A2(n382), .B1(n384), .B2(n684), .ZN(n128) );
  INV_X1 U324 ( .A(n128), .ZN(n132) );
  NAND2_X1 U325 ( .A1(n132), .A2(n339), .ZN(n478) );
  NAND2_X1 U327 ( .A1(A[20]), .A2(n25), .ZN(n435) );
  NAND2_X1 U328 ( .A1(A[19]), .A2(n31), .ZN(n390) );
  NAND3_X1 U330 ( .A1(n508), .A2(n435), .A3(n390), .ZN(n380) );
  INV_X1 U331 ( .A(n674), .ZN(n580) );
  OAI21_X1 U333 ( .B1(n580), .B2(n331), .A(n178), .ZN(n129) );
  AOI221_X1 U335 ( .B1(n241), .B2(n478), .C1(n201), .C2(n380), .A(n129), .ZN(
        n137) );
  INV_X1 U337 ( .A(A[7]), .ZN(n737) );
  OAI221_X1 U338 ( .B1(n738), .B2(n22), .C1(n737), .C2(n29), .A(n513), .ZN(
        n675) );
  NAND2_X1 U339 ( .A1(A[16]), .A2(n25), .ZN(n356) );
  NAND2_X1 U340 ( .A1(A[15]), .A2(n31), .ZN(n303) );
  NAND3_X1 U342 ( .A1(n507), .A2(n356), .A3(n303), .ZN(n182) );
  NAND2_X1 U343 ( .A1(A[31]), .A2(n30), .ZN(n699) );
  OAI21_X1 U345 ( .B1(n699), .B2(n579), .A(n132), .ZN(n477) );
  AOI222_X1 U347 ( .A1(n1), .A2(n675), .B1(n310), .B2(n182), .C1(n131), .C2(
        n477), .ZN(n135) );
  AOI222_X1 U348 ( .A1(N98), .A2(n4), .B1(n162), .B2(n308), .C1(n163), .C2(
        n212), .ZN(n134) );
  AOI222_X1 U349 ( .A1(n157), .A2(A[7]), .B1(N66), .B2(n9), .C1(B[7]), .C2(
        n159), .ZN(n133) );
  NAND4_X1 U350 ( .A1(n137), .A2(n135), .A3(n134), .A4(n133), .ZN(RES[7]) );
  NAND2_X1 U351 ( .A1(n246), .A2(n213), .ZN(n281) );
  OAI22_X1 U352 ( .A1(n10), .A2(n326), .B1(n327), .B2(n684), .ZN(n505) );
  INV_X1 U353 ( .A(n505), .ZN(n139) );
  INV_X1 U354 ( .A(n131), .ZN(n228) );
  OAI21_X1 U355 ( .B1(n139), .B2(n228), .A(n178), .ZN(n138) );
  AOI221_X1 U356 ( .B1(n702), .B2(n595), .C1(n596), .C2(n320), .A(n138), .ZN(
        n147) );
  NAND2_X1 U357 ( .A1(n139), .A2(n339), .ZN(n510) );
  INV_X1 U358 ( .A(A[8]), .ZN(n736) );
  OAI221_X1 U360 ( .B1(n737), .B2(n22), .C1(n736), .C2(n29), .A(n497), .ZN(
        n423) );
  AOI222_X1 U362 ( .A1(n310), .A2(n323), .B1(n241), .B2(n510), .C1(n2), .C2(
        n423), .ZN(n145) );
  INV_X1 U363 ( .A(n150), .ZN(n141) );
  OAI22_X1 U364 ( .A1(n141), .A2(n185), .B1(n140), .B2(n306), .ZN(n142) );
  AOI221_X1 U365 ( .B1(n151), .B2(n212), .C1(N99), .C2(n4), .A(n142), .ZN(n144) );
  AOI222_X1 U366 ( .A1(n146), .A2(A[8]), .B1(N67), .B2(n9), .C1(B[8]), .C2(
        n148), .ZN(n143) );
  NAND4_X1 U367 ( .A1(n147), .A2(n145), .A3(n144), .A4(n143), .ZN(RES[8]) );
  NAND2_X1 U368 ( .A1(n149), .A2(n16), .ZN(n152) );
  OAI211_X1 U370 ( .C1(n338), .C2(n684), .A(n339), .B(n152), .ZN(n555) );
  OAI21_X1 U372 ( .B1(n644), .B2(n684), .A(n152), .ZN(n531) );
  AOI221_X1 U373 ( .B1(n241), .B2(n555), .C1(n131), .C2(n531), .A(n153), .ZN(
        n160) );
  INV_X1 U374 ( .A(n626), .ZN(n249) );
  INV_X1 U375 ( .A(A[9]), .ZN(n735) );
  OAI221_X1 U376 ( .B1(n736), .B2(n22), .C1(n735), .C2(n29), .A(n489), .ZN(
        n441) );
  INV_X1 U378 ( .A(n441), .ZN(n628) );
  OAI222_X1 U379 ( .A1(n249), .A2(n684), .B1(n11), .B2(n628), .C1(n154), .C2(
        n579), .ZN(n556) );
  AOI222_X1 U381 ( .A1(n308), .A2(n255), .B1(n246), .B2(n556), .C1(n310), .C2(
        n336), .ZN(n158) );
  AOI222_X1 U385 ( .A1(N100), .A2(n4), .B1(n201), .B2(n257), .C1(n136), .C2(
        n212), .ZN(n156) );
  AOI222_X1 U386 ( .A1(n121), .A2(A[9]), .B1(N68), .B2(n9), .C1(B[9]), .C2(
        n127), .ZN(n155) );
  NAND4_X1 U387 ( .A1(n160), .A2(n158), .A3(n156), .A4(n155), .ZN(RES[9]) );
  NAND2_X1 U388 ( .A1(n161), .A2(n15), .ZN(n166) );
  OAI21_X1 U389 ( .B1(n669), .B2(n684), .A(n166), .ZN(n572) );
  INV_X1 U391 ( .A(n572), .ZN(n164) );
  OAI21_X1 U393 ( .B1(n164), .B2(n228), .A(n178), .ZN(n165) );
  AOI221_X1 U394 ( .B1(n595), .B2(n649), .C1(n596), .C2(n650), .A(n165), .ZN(
        n174) );
  OAI211_X1 U396 ( .C1(n663), .C2(n684), .A(n339), .B(n166), .ZN(n573) );
  INV_X1 U398 ( .A(A[10]), .ZN(n734) );
  OAI221_X1 U399 ( .B1(n735), .B2(n22), .C1(n734), .C2(n29), .A(n527), .ZN(
        n459) );
  AOI222_X1 U400 ( .A1(n310), .A2(n362), .B1(n241), .B2(n573), .C1(n3), .C2(
        n459), .ZN(n173) );
  INV_X1 U401 ( .A(n167), .ZN(n727) );
  OAI22_X1 U403 ( .A1(n363), .A2(n306), .B1(n727), .B2(n185), .ZN(n168) );
  AOI221_X1 U405 ( .B1(n175), .B2(n212), .C1(N101), .C2(n4), .A(n168), .ZN(
        n171) );
  AOI222_X1 U407 ( .A1(n518), .A2(A[10]), .B1(N69), .B2(n9), .C1(B[10]), .C2(
        n519), .ZN(n169) );
  NAND4_X1 U408 ( .A1(n174), .A2(n173), .A3(n171), .A4(n169), .ZN(RES[10]) );
  NAND2_X1 U411 ( .A1(n177), .A2(n15), .ZN(n590) );
  NAND3_X1 U412 ( .A1(n241), .A2(A[31]), .A3(n10), .ZN(n179) );
  NAND2_X1 U414 ( .A1(n179), .A2(n178), .ZN(n230) );
  INV_X1 U415 ( .A(n230), .ZN(n274) );
  OAI21_X1 U416 ( .B1(n590), .B2(n229), .A(n274), .ZN(n180) );
  AOI221_X1 U417 ( .B1(n595), .B2(n674), .C1(n596), .C2(n675), .A(n180), .ZN(
        n191) );
  OAI21_X1 U418 ( .B1(n699), .B2(n684), .A(n590), .ZN(n597) );
  INV_X1 U419 ( .A(A[11]), .ZN(n221) );
  AOI22_X1 U420 ( .A1(n46), .A2(A[8]), .B1(n39), .B2(A[9]), .ZN(n181) );
  OAI221_X1 U422 ( .B1(n734), .B2(n22), .C1(n29), .C2(n221), .A(n181), .ZN(
        n578) );
  AOI222_X1 U423 ( .A1(n310), .A2(n380), .B1(n131), .B2(n597), .C1(n3), .C2(
        n578), .ZN(n190) );
  INV_X1 U424 ( .A(n182), .ZN(n726) );
  OAI22_X1 U426 ( .A1(n382), .A2(n306), .B1(n726), .B2(n185), .ZN(n187) );
  AOI221_X1 U427 ( .B1(n162), .B2(n212), .C1(N102), .C2(n4), .A(n187), .ZN(
        n189) );
  AOI222_X1 U429 ( .A1(n503), .A2(A[11]), .B1(N70), .B2(n9), .C1(B[11]), .C2(
        n504), .ZN(n188) );
  NAND4_X1 U430 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(RES[11]) );
  NAND2_X1 U431 ( .A1(FUNC[2]), .A2(n705), .ZN(n193) );
  INV_X1 U432 ( .A(n193), .ZN(n343) );
  NAND2_X1 U434 ( .A1(n343), .A2(n194), .ZN(n123) );
  NAND2_X1 U435 ( .A1(n199), .A2(n344), .ZN(n130) );
  AOI222_X1 U436 ( .A1(n310), .A2(n324), .B1(n308), .B2(n323), .C1(n201), .C2(
        n200), .ZN(n238) );
  AOI222_X1 U437 ( .A1(N71), .A2(n8), .B1(n212), .B2(n150), .C1(N103), .C2(n5), 
        .ZN(n237) );
  INV_X1 U438 ( .A(n423), .ZN(n610) );
  AOI22_X1 U445 ( .A1(n46), .A2(A[9]), .B1(A[10]), .B2(n39), .ZN(n215) );
  OAI211_X1 U447 ( .C1(n22), .C2(n221), .A(n216), .B(n215), .ZN(n511) );
  INV_X1 U454 ( .A(n511), .ZN(n609) );
  MUX2_X1 U455 ( .A(n64), .B(n51), .S(B[12]), .Z(n222) );
  OAI21_X1 U456 ( .B1(n56), .B2(n222), .A(A[12]), .ZN(n223) );
  OAI221_X1 U459 ( .B1(n610), .B2(n331), .C1(n609), .C2(n330), .A(n223), .ZN(
        n234) );
  INV_X1 U460 ( .A(A[12]), .ZN(n710) );
  AOI21_X1 U462 ( .B1(n65), .B2(n710), .A(n56), .ZN(n226) );
  INV_X1 U463 ( .A(B[12]), .ZN(n225) );
  NAND3_X1 U465 ( .A1(n246), .A2(B[3]), .A3(n399), .ZN(n224) );
  OAI21_X1 U466 ( .B1(n226), .B2(n225), .A(n224), .ZN(n233) );
  NAND2_X1 U470 ( .A1(n227), .A2(n14), .ZN(n604) );
  AOI21_X1 U471 ( .B1(n229), .B2(n228), .A(n604), .ZN(n231) );
  NOR4_X1 U474 ( .A1(n234), .A2(n233), .A3(n231), .A4(n230), .ZN(n236) );
  NAND3_X1 U475 ( .A1(n238), .A2(n237), .A3(n236), .ZN(RES[12]) );
  OAI21_X1 U476 ( .B1(A[13]), .B2(n58), .A(n55), .ZN(n244) );
  NAND2_X1 U479 ( .A1(n131), .A2(n14), .ZN(n240) );
  INV_X1 U480 ( .A(n240), .ZN(n301) );
  NAND2_X1 U481 ( .A1(n241), .A2(n13), .ZN(n275) );
  OAI21_X1 U482 ( .B1(n338), .B2(n275), .A(n274), .ZN(n242) );
  AOI221_X1 U483 ( .B1(B[13]), .B2(n244), .C1(n301), .C2(n243), .A(n242), .ZN(
        n273) );
  MUX2_X1 U484 ( .A(n59), .B(n50), .S(B[13]), .Z(n245) );
  NAND2_X1 U485 ( .A1(n245), .A2(n55), .ZN(n251) );
  NAND2_X1 U486 ( .A1(n246), .A2(n232), .ZN(n248) );
  OAI22_X1 U487 ( .A1(n628), .A2(n331), .B1(n249), .B2(n281), .ZN(n250) );
  AOI221_X1 U488 ( .B1(A[13]), .B2(n251), .C1(n598), .C2(n625), .A(n250), .ZN(
        n262) );
  OAI211_X1 U489 ( .C1(n710), .C2(n22), .A(n488), .B(n252), .ZN(n624) );
  INV_X1 U490 ( .A(n255), .ZN(n728) );
  OAI22_X1 U491 ( .A1(n341), .A2(n306), .B1(n728), .B2(n305), .ZN(n256) );
  AOI221_X1 U492 ( .B1(n2), .B2(n624), .C1(n308), .C2(n336), .A(n256), .ZN(
        n261) );
  AOI222_X1 U493 ( .A1(N72), .A2(n8), .B1(n310), .B2(n257), .C1(N104), .C2(n6), 
        .ZN(n260) );
  NAND4_X1 U494 ( .A1(n273), .A2(n262), .A3(n261), .A4(n260), .ZN(RES[13]) );
  OAI21_X1 U495 ( .B1(A[14]), .B2(n58), .A(n54), .ZN(n278) );
  OAI21_X1 U496 ( .B1(n663), .B2(n275), .A(n274), .ZN(n276) );
  AOI221_X1 U497 ( .B1(B[14]), .B2(n278), .C1(n301), .C2(n277), .A(n276), .ZN(
        n292) );
  MUX2_X1 U498 ( .A(n60), .B(n50), .S(B[14]), .Z(n280) );
  NAND2_X1 U499 ( .A1(n280), .A2(n55), .ZN(n283) );
  INV_X1 U500 ( .A(n459), .ZN(n652) );
  INV_X1 U501 ( .A(n650), .ZN(n562) );
  OAI22_X1 U502 ( .A1(n652), .A2(n331), .B1(n562), .B2(n281), .ZN(n282) );
  AOI221_X1 U503 ( .B1(A[14]), .B2(n283), .C1(n598), .C2(n649), .A(n282), .ZN(
        n291) );
  NAND3_X1 U504 ( .A1(n474), .A2(n286), .A3(n284), .ZN(n648) );
  OAI22_X1 U505 ( .A1(n365), .A2(n306), .B1(n727), .B2(n305), .ZN(n287) );
  AOI221_X1 U506 ( .B1(n2), .B2(n648), .C1(n308), .C2(n362), .A(n287), .ZN(
        n290) );
  AOI222_X1 U507 ( .A1(N73), .A2(n8), .B1(n310), .B2(n288), .C1(N105), .C2(n6), 
        .ZN(n289) );
  NAND4_X1 U508 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(RES[14]) );
  INV_X1 U509 ( .A(n699), .ZN(n679) );
  MUX2_X1 U510 ( .A(n60), .B(n50), .S(B[15]), .Z(n293) );
  NAND2_X1 U511 ( .A1(n293), .A2(n55), .ZN(n300) );
  INV_X1 U512 ( .A(A[15]), .ZN(n294) );
  AOI21_X1 U513 ( .B1(n64), .B2(n294), .A(n56), .ZN(n298) );
  INV_X1 U514 ( .A(B[15]), .ZN(n297) );
  NAND3_X1 U515 ( .A1(A[31]), .A2(n349), .A3(n296), .ZN(n582) );
  OAI21_X1 U516 ( .B1(n298), .B2(n297), .A(n582), .ZN(n299) );
  AOI221_X1 U517 ( .B1(n301), .B2(n679), .C1(A[15]), .C2(n300), .A(n299), .ZN(
        n314) );
  AOI222_X1 U518 ( .A1(n596), .A2(n578), .B1(n598), .B2(n674), .C1(n595), .C2(
        n675), .ZN(n313) );
  NAND3_X1 U519 ( .A1(n465), .A2(n304), .A3(n303), .ZN(n673) );
  OAI22_X1 U520 ( .A1(n384), .A2(n306), .B1(n726), .B2(n305), .ZN(n307) );
  AOI221_X1 U521 ( .B1(n2), .B2(n673), .C1(n308), .C2(n380), .A(n307), .ZN(
        n312) );
  AOI222_X1 U522 ( .A1(N74), .A2(n8), .B1(n310), .B2(n309), .C1(N106), .C2(n6), 
        .ZN(n311) );
  NAND4_X1 U523 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(RES[15]) );
  NAND2_X1 U524 ( .A1(n606), .A2(n703), .ZN(n398) );
  INV_X1 U525 ( .A(n398), .ZN(n586) );
  NAND2_X1 U526 ( .A1(n586), .A2(n13), .ZN(n315) );
  INV_X1 U527 ( .A(n315), .ZN(n468) );
  OAI21_X1 U528 ( .B1(A[16]), .B2(n58), .A(n54), .ZN(n316) );
  INV_X1 U529 ( .A(n582), .ZN(n563) );
  AOI221_X1 U530 ( .B1(n468), .B2(n702), .C1(B[16]), .C2(n316), .A(n563), .ZN(
        n335) );
  MUX2_X1 U531 ( .A(n60), .B(n50), .S(B[16]), .Z(n318) );
  INV_X1 U532 ( .A(A[16]), .ZN(n317) );
  AOI21_X1 U533 ( .B1(n318), .B2(n54), .A(n317), .ZN(n319) );
  AOI221_X1 U534 ( .B1(n595), .B2(n423), .C1(n598), .C2(n320), .A(n319), .ZN(
        n334) );
  NAND3_X1 U535 ( .A1(n454), .A2(n322), .A3(n321), .ZN(n514) );
  INV_X1 U536 ( .A(n514), .ZN(n614) );
  INV_X1 U537 ( .A(n232), .ZN(n744) );
  AOI22_X1 U538 ( .A1(n701), .A2(n324), .B1(n323), .B2(n16), .ZN(n325) );
  OAI221_X1 U539 ( .B1(n744), .B2(n327), .C1(n326), .C2(n579), .A(n325), .ZN(
        n328) );
  INV_X1 U540 ( .A(n328), .ZN(n455) );
  OAI222_X1 U541 ( .A1(n609), .A2(n331), .B1(n614), .B2(n330), .C1(n455), .C2(
        n329), .ZN(n332) );
  AOI221_X1 U542 ( .B1(N107), .B2(n5), .C1(N75), .C2(n7), .A(n332), .ZN(n333)
         );
  NAND3_X1 U543 ( .A1(n335), .A2(n334), .A3(n333), .ZN(RES[16]) );
  INV_X1 U544 ( .A(n336), .ZN(n340) );
  OAI222_X1 U545 ( .A1(n341), .A2(n579), .B1(n11), .B2(n340), .C1(n337), .C2(
        n684), .ZN(n342) );
  INV_X1 U546 ( .A(n342), .ZN(n345) );
  OAI21_X1 U547 ( .B1(n338), .B2(n744), .A(n345), .ZN(n409) );
  NAND2_X1 U548 ( .A1(n344), .A2(n343), .ZN(n411) );
  OAI21_X1 U549 ( .B1(n744), .B2(n644), .A(n345), .ZN(n408) );
  OAI21_X1 U550 ( .B1(A[17]), .B2(n58), .A(n54), .ZN(n346) );
  AOI221_X1 U551 ( .B1(n468), .B2(n625), .C1(B[17]), .C2(n346), .A(n563), .ZN(
        n361) );
  INV_X1 U552 ( .A(n411), .ZN(n347) );
  NAND2_X1 U553 ( .A1(n350), .A2(n347), .ZN(n348) );
  NAND2_X1 U554 ( .A1(n350), .A2(n349), .ZN(n351) );
  MUX2_X1 U555 ( .A(n59), .B(n50), .S(B[17]), .Z(n353) );
  INV_X1 U556 ( .A(A[17]), .ZN(n352) );
  AOI21_X1 U557 ( .B1(n353), .B2(n54), .A(n352), .ZN(n354) );
  AOI221_X1 U558 ( .B1(n641), .B2(n408), .C1(n637), .C2(n409), .A(n354), .ZN(
        n360) );
  AOI22_X1 U559 ( .A1(A[14]), .A2(n46), .B1(A[15]), .B2(n39), .ZN(n355) );
  NAND3_X1 U560 ( .A1(n357), .A2(n356), .A3(n355), .ZN(n630) );
  AOI222_X1 U561 ( .A1(n595), .A2(n441), .B1(n2), .B2(n630), .C1(n598), .C2(
        n626), .ZN(n359) );
  AOI222_X1 U562 ( .A1(N76), .A2(n8), .B1(n596), .B2(n624), .C1(N108), .C2(n6), 
        .ZN(n358) );
  NAND4_X1 U563 ( .A1(n361), .A2(n360), .A3(n359), .A4(n358), .ZN(RES[17]) );
  INV_X1 U564 ( .A(n362), .ZN(n364) );
  OAI222_X1 U565 ( .A1(n365), .A2(n579), .B1(n11), .B2(n364), .C1(n363), .C2(
        n684), .ZN(n366) );
  INV_X1 U566 ( .A(n366), .ZN(n367) );
  OAI21_X1 U567 ( .B1(n744), .B2(n663), .A(n367), .ZN(n267) );
  OAI21_X1 U568 ( .B1(n744), .B2(n669), .A(n367), .ZN(n266) );
  OAI21_X1 U569 ( .B1(A[18]), .B2(n59), .A(n54), .ZN(n368) );
  AOI221_X1 U570 ( .B1(n468), .B2(n649), .C1(B[18]), .C2(n368), .A(n563), .ZN(
        n379) );
  AOI22_X1 U571 ( .A1(A[15]), .A2(n46), .B1(A[16]), .B2(n39), .ZN(n369) );
  NAND3_X1 U572 ( .A1(n371), .A2(n370), .A3(n369), .ZN(n654) );
  MUX2_X1 U573 ( .A(n59), .B(n50), .S(B[18]), .Z(n373) );
  INV_X1 U574 ( .A(A[18]), .ZN(n372) );
  AOI21_X1 U575 ( .B1(n373), .B2(n54), .A(n372), .ZN(n374) );
  AOI221_X1 U576 ( .B1(n637), .B2(n267), .C1(n1), .C2(n654), .A(n374), .ZN(
        n377) );
  AOI222_X1 U579 ( .A1(n595), .A2(n459), .B1(n641), .B2(n266), .C1(n598), .C2(
        n650), .ZN(n376) );
  AOI222_X1 U580 ( .A1(N77), .A2(n8), .B1(n596), .B2(n648), .C1(N109), .C2(n6), 
        .ZN(n375) );
  NAND4_X1 U581 ( .A1(n379), .A2(n377), .A3(n376), .A4(n375), .ZN(RES[18]) );
  INV_X1 U582 ( .A(n380), .ZN(n381) );
  OAI22_X1 U583 ( .A1(n382), .A2(n684), .B1(n10), .B2(n381), .ZN(n383) );
  INV_X1 U584 ( .A(n383), .ZN(n385) );
  OAI211_X1 U585 ( .C1(n384), .C2(n579), .A(n385), .B(n378), .ZN(n207) );
  MUX2_X1 U586 ( .A(n384), .B(n699), .S(B[2]), .Z(n386) );
  OAI21_X1 U587 ( .B1(n711), .B2(n386), .A(n385), .ZN(n205) );
  OAI21_X1 U588 ( .B1(A[19]), .B2(n59), .A(n54), .ZN(n387) );
  AOI221_X1 U589 ( .B1(n468), .B2(n674), .C1(B[19]), .C2(n387), .A(n563), .ZN(
        n397) );
  AOI22_X1 U590 ( .A1(A[16]), .A2(n46), .B1(A[17]), .B2(n39), .ZN(n388) );
  NAND3_X1 U591 ( .A1(n390), .A2(n389), .A3(n388), .ZN(n681) );
  MUX2_X1 U592 ( .A(n59), .B(n50), .S(B[19]), .Z(n392) );
  INV_X1 U593 ( .A(A[19]), .ZN(n391) );
  AOI21_X1 U594 ( .B1(n392), .B2(n54), .A(n391), .ZN(n393) );
  AOI221_X1 U595 ( .B1(n637), .B2(n207), .C1(n2), .C2(n681), .A(n393), .ZN(
        n396) );
  AOI222_X1 U596 ( .A1(n595), .A2(n578), .B1(n641), .B2(n205), .C1(n598), .C2(
        n675), .ZN(n395) );
  AOI222_X1 U597 ( .A1(N78), .A2(n8), .B1(n596), .B2(n673), .C1(N110), .C2(n6), 
        .ZN(n394) );
  NAND4_X1 U598 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(RES[19]) );
  OAI21_X1 U599 ( .B1(A[20]), .B2(n59), .A(n54), .ZN(n403) );
  NOR2_X1 U600 ( .A1(B[3]), .A2(n398), .ZN(n400) );
  AOI221_X1 U601 ( .B1(B[20]), .B2(n403), .C1(n400), .C2(n399), .A(n563), .ZN(
        n428) );
  AOI22_X1 U602 ( .A1(A[17]), .A2(n46), .B1(A[18]), .B2(n39), .ZN(n404) );
  NAND3_X1 U603 ( .A1(n418), .A2(n417), .A3(n404), .ZN(n611) );
  MUX2_X1 U604 ( .A(n59), .B(n50), .S(B[20]), .Z(n420) );
  INV_X1 U605 ( .A(A[20]), .ZN(n419) );
  AOI21_X1 U606 ( .B1(n420), .B2(n53), .A(n419), .ZN(n421) );
  AOI221_X1 U607 ( .B1(n2), .B2(n611), .C1(n641), .C2(n422), .A(n421), .ZN(
        n427) );
  AOI222_X1 U608 ( .A1(n595), .A2(n511), .B1(n637), .B2(n424), .C1(n598), .C2(
        n423), .ZN(n426) );
  AOI222_X1 U609 ( .A1(N79), .A2(n7), .B1(n596), .B2(n514), .C1(N111), .C2(n6), 
        .ZN(n425) );
  NAND4_X1 U610 ( .A1(n428), .A2(n427), .A3(n426), .A4(n425), .ZN(RES[20]) );
  NAND2_X1 U611 ( .A1(n586), .A2(n701), .ZN(n429) );
  INV_X1 U612 ( .A(n429), .ZN(n469) );
  INV_X1 U613 ( .A(A[21]), .ZN(n436) );
  AOI21_X1 U614 ( .B1(n65), .B2(n436), .A(n56), .ZN(n431) );
  INV_X1 U615 ( .A(B[21]), .ZN(n430) );
  OAI21_X1 U616 ( .B1(n431), .B2(n430), .A(n582), .ZN(n432) );
  AOI221_X1 U617 ( .B1(n469), .B2(n625), .C1(n468), .C2(n626), .A(n432), .ZN(
        n445) );
  AOI22_X1 U618 ( .A1(A[18]), .A2(n46), .B1(A[19]), .B2(n39), .ZN(n433) );
  NAND3_X1 U619 ( .A1(n435), .A2(n434), .A3(n433), .ZN(n631) );
  MUX2_X1 U620 ( .A(n59), .B(n50), .S(B[21]), .Z(n437) );
  AOI21_X1 U621 ( .B1(n437), .B2(n54), .A(n436), .ZN(n438) );
  AOI221_X1 U622 ( .B1(n637), .B2(n439), .C1(n1), .C2(n631), .A(n438), .ZN(
        n444) );
  AOI222_X1 U623 ( .A1(n598), .A2(n441), .B1(n641), .B2(n440), .C1(n596), .C2(
        n630), .ZN(n443) );
  AOI222_X1 U624 ( .A1(N80), .A2(n7), .B1(n595), .B2(n624), .C1(N112), .C2(n6), 
        .ZN(n442) );
  NAND4_X1 U625 ( .A1(n445), .A2(n444), .A3(n443), .A4(n442), .ZN(RES[21]) );
  INV_X1 U626 ( .A(A[22]), .ZN(n452) );
  AOI21_X1 U627 ( .B1(n64), .B2(n452), .A(n56), .ZN(n447) );
  INV_X1 U628 ( .A(B[22]), .ZN(n446) );
  OAI21_X1 U629 ( .B1(n447), .B2(n446), .A(n582), .ZN(n448) );
  AOI221_X1 U630 ( .B1(n469), .B2(n649), .C1(n468), .C2(n650), .A(n448), .ZN(
        n463) );
  AOI22_X1 U631 ( .A1(A[19]), .A2(n46), .B1(A[20]), .B2(n39), .ZN(n449) );
  NAND3_X1 U632 ( .A1(n451), .A2(n450), .A3(n449), .ZN(n655) );
  MUX2_X1 U633 ( .A(n59), .B(n49), .S(B[22]), .Z(n453) );
  AOI21_X1 U634 ( .B1(n453), .B2(n54), .A(n452), .ZN(n456) );
  AOI221_X1 U635 ( .B1(n596), .B2(n654), .C1(n1), .C2(n655), .A(n456), .ZN(
        n462) );
  AOI222_X1 U636 ( .A1(n598), .A2(n459), .B1(n637), .B2(n458), .C1(n641), .C2(
        n457), .ZN(n461) );
  AOI222_X1 U637 ( .A1(N81), .A2(n8), .B1(n595), .B2(n648), .C1(N113), .C2(n6), 
        .ZN(n460) );
  NAND4_X1 U638 ( .A1(n463), .A2(n462), .A3(n461), .A4(n460), .ZN(RES[22]) );
  INV_X1 U639 ( .A(A[23]), .ZN(n473) );
  AOI21_X1 U640 ( .B1(n65), .B2(n473), .A(n56), .ZN(n466) );
  INV_X1 U641 ( .A(B[23]), .ZN(n464) );
  OAI21_X1 U642 ( .B1(n466), .B2(n464), .A(n582), .ZN(n467) );
  AOI221_X1 U643 ( .B1(n469), .B2(n674), .C1(n468), .C2(n675), .A(n467), .ZN(
        n490) );
  AOI22_X1 U644 ( .A1(A[20]), .A2(n46), .B1(A[21]), .B2(n39), .ZN(n470) );
  NAND3_X1 U645 ( .A1(n472), .A2(n471), .A3(n470), .ZN(n682) );
  MUX2_X1 U646 ( .A(n59), .B(n49), .S(B[23]), .Z(n475) );
  AOI21_X1 U647 ( .B1(n475), .B2(n53), .A(n473), .ZN(n476) );
  AOI221_X1 U648 ( .B1(n596), .B2(n681), .C1(n1), .C2(n682), .A(n476), .ZN(
        n486) );
  AOI222_X1 U649 ( .A1(n598), .A2(n578), .B1(n637), .B2(n478), .C1(n641), .C2(
        n477), .ZN(n481) );
  AOI222_X1 U650 ( .A1(N82), .A2(n7), .B1(n595), .B2(n673), .C1(N114), .C2(n5), 
        .ZN(n479) );
  NAND4_X1 U651 ( .A1(n490), .A2(n486), .A3(n481), .A4(n479), .ZN(RES[23]) );
  OAI222_X1 U652 ( .A1(n492), .A2(n684), .B1(n11), .B2(n610), .C1(n579), .C2(
        n491), .ZN(n494) );
  OAI21_X1 U653 ( .B1(A[24]), .B2(n58), .A(n54), .ZN(n493) );
  AOI221_X1 U654 ( .B1(n586), .B2(n494), .C1(B[24]), .C2(n493), .A(n563), .ZN(
        n525) );
  AOI22_X1 U655 ( .A1(A[21]), .A2(n46), .B1(A[22]), .B2(n39), .ZN(n495) );
  NAND3_X1 U656 ( .A1(n499), .A2(n498), .A3(n495), .ZN(n612) );
  MUX2_X1 U657 ( .A(n59), .B(n49), .S(B[24]), .Z(n501) );
  INV_X1 U658 ( .A(A[24]), .ZN(n500) );
  AOI21_X1 U659 ( .B1(n501), .B2(n53), .A(n500), .ZN(n502) );
  AOI221_X1 U660 ( .B1(n2), .B2(n612), .C1(n641), .C2(n505), .A(n502), .ZN(
        n517) );
  AOI222_X1 U661 ( .A1(n598), .A2(n511), .B1(n596), .B2(n611), .C1(n637), .C2(
        n510), .ZN(n516) );
  AOI222_X1 U662 ( .A1(N83), .A2(n7), .B1(n595), .B2(n514), .C1(N115), .C2(n5), 
        .ZN(n515) );
  NAND4_X1 U663 ( .A1(n525), .A2(n517), .A3(n516), .A4(n515), .ZN(RES[24]) );
  OAI21_X1 U664 ( .B1(A[25]), .B2(n59), .A(n54), .ZN(n526) );
  AOI221_X1 U665 ( .B1(n641), .B2(n531), .C1(B[25]), .C2(n526), .A(n563), .ZN(
        n560) );
  AOI22_X1 U666 ( .A1(A[22]), .A2(n46), .B1(A[23]), .B2(n39), .ZN(n532) );
  NAND3_X1 U667 ( .A1(n535), .A2(n533), .A3(n532), .ZN(n632) );
  MUX2_X1 U668 ( .A(n59), .B(n49), .S(B[25]), .Z(n548) );
  INV_X1 U669 ( .A(A[25]), .ZN(n546) );
  AOI21_X1 U670 ( .B1(n548), .B2(n53), .A(n546), .ZN(n554) );
  AOI221_X1 U671 ( .B1(n596), .B2(n631), .C1(n1), .C2(n632), .A(n554), .ZN(
        n559) );
  AOI222_X1 U672 ( .A1(n586), .A2(n556), .B1(n637), .B2(n555), .C1(n595), .C2(
        n630), .ZN(n558) );
  AOI222_X1 U673 ( .A1(N84), .A2(n7), .B1(n598), .B2(n624), .C1(N116), .C2(n5), 
        .ZN(n557) );
  NAND4_X1 U674 ( .A1(n560), .A2(n559), .A3(n558), .A4(n557), .ZN(RES[25]) );
  OAI222_X1 U675 ( .A1(n562), .A2(n684), .B1(n11), .B2(n652), .C1(n561), .C2(
        n579), .ZN(n565) );
  OAI21_X1 U676 ( .B1(A[26]), .B2(n58), .A(n54), .ZN(n564) );
  AOI221_X1 U677 ( .B1(n586), .B2(n565), .C1(B[26]), .C2(n564), .A(n563), .ZN(
        n577) );
  AOI22_X1 U678 ( .A1(A[23]), .A2(n46), .B1(A[24]), .B2(n39), .ZN(n566) );
  NAND3_X1 U679 ( .A1(n568), .A2(n567), .A3(n566), .ZN(n656) );
  MUX2_X1 U680 ( .A(n59), .B(n49), .S(B[26]), .Z(n570) );
  INV_X1 U681 ( .A(A[26]), .ZN(n569) );
  AOI21_X1 U682 ( .B1(n570), .B2(n53), .A(n569), .ZN(n571) );
  AOI221_X1 U683 ( .B1(n2), .B2(n656), .C1(n641), .C2(n572), .A(n571), .ZN(
        n576) );
  AOI222_X1 U684 ( .A1(n637), .A2(n573), .B1(n596), .B2(n655), .C1(n595), .C2(
        n654), .ZN(n575) );
  AOI222_X1 U685 ( .A1(N85), .A2(n7), .B1(n598), .B2(n648), .C1(N117), .C2(n5), 
        .ZN(n574) );
  NAND4_X1 U686 ( .A1(n577), .A2(n576), .A3(n575), .A4(n574), .ZN(RES[26]) );
  INV_X1 U687 ( .A(n675), .ZN(n581) );
  INV_X1 U688 ( .A(n578), .ZN(n677) );
  OAI222_X1 U689 ( .A1(n581), .A2(n684), .B1(n11), .B2(n677), .C1(n580), .C2(
        n579), .ZN(n585) );
  OAI21_X1 U690 ( .B1(A[27]), .B2(n59), .A(n54), .ZN(n584) );
  NAND3_X1 U691 ( .A1(n637), .A2(A[31]), .A3(n10), .ZN(n583) );
  NAND2_X1 U692 ( .A1(n583), .A2(n582), .ZN(n603) );
  AOI221_X1 U693 ( .B1(n586), .B2(n585), .C1(B[27]), .C2(n584), .A(n603), .ZN(
        n602) );
  AOI22_X1 U694 ( .A1(A[24]), .A2(n46), .B1(A[25]), .B2(n39), .ZN(n587) );
  NAND3_X1 U695 ( .A1(n589), .A2(n588), .A3(n587), .ZN(n680) );
  INV_X1 U696 ( .A(n590), .ZN(n593) );
  MUX2_X1 U697 ( .A(n59), .B(n49), .S(B[27]), .Z(n591) );
  AOI21_X1 U698 ( .B1(n591), .B2(n53), .A(n709), .ZN(n592) );
  AOI221_X1 U699 ( .B1(n2), .B2(n680), .C1(n593), .C2(n637), .A(n592), .ZN(
        n601) );
  AOI222_X1 U700 ( .A1(n641), .A2(n597), .B1(n596), .B2(n682), .C1(n595), .C2(
        n681), .ZN(n600) );
  AOI222_X1 U701 ( .A1(N86), .A2(n7), .B1(n598), .B2(n673), .C1(N118), .C2(n5), 
        .ZN(n599) );
  NAND4_X1 U702 ( .A1(n602), .A2(n601), .A3(n600), .A4(n599), .ZN(RES[27]) );
  INV_X1 U703 ( .A(n603), .ZN(n661) );
  INV_X1 U704 ( .A(n604), .ZN(n605) );
  OAI21_X1 U705 ( .B1(n641), .B2(n637), .A(n605), .ZN(n623) );
  OAI21_X1 U706 ( .B1(A[28]), .B2(n59), .A(n54), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n606), .A2(n714), .ZN(n607) );
  INV_X1 U708 ( .A(n607), .ZN(n690) );
  OAI222_X1 U709 ( .A1(n610), .A2(n684), .B1(n10), .B2(n609), .C1(n711), .C2(
        n608), .ZN(n616) );
  AOI22_X1 U710 ( .A1(n701), .A2(n612), .B1(n213), .B2(n611), .ZN(n613) );
  OAI221_X1 U711 ( .B1(n744), .B2(n614), .C1(n295), .C2(n11), .A(n613), .ZN(
        n615) );
  MUX2_X1 U712 ( .A(n616), .B(n615), .S(n210), .Z(n617) );
  AOI22_X1 U713 ( .A1(B[28]), .A2(n618), .B1(n690), .B2(n617), .ZN(n622) );
  MUX2_X1 U714 ( .A(n59), .B(n49), .S(B[28]), .Z(n619) );
  AOI21_X1 U715 ( .B1(n619), .B2(n53), .A(n708), .ZN(n620) );
  AOI221_X1 U716 ( .B1(N87), .B2(n8), .C1(N119), .C2(n4), .A(n620), .ZN(n621)
         );
  NAND4_X1 U717 ( .A1(n661), .A2(n623), .A3(n622), .A4(n621), .ZN(RES[28]) );
  OAI21_X1 U718 ( .B1(A[29]), .B2(n59), .A(n54), .ZN(n640) );
  INV_X1 U719 ( .A(n624), .ZN(n629) );
  AOI22_X1 U720 ( .A1(n213), .A2(n626), .B1(n625), .B2(n232), .ZN(n627) );
  OAI221_X1 U721 ( .B1(n10), .B2(n629), .C1(n628), .C2(n684), .A(n627), .ZN(
        n636) );
  INV_X1 U722 ( .A(n630), .ZN(n634) );
  AOI22_X1 U723 ( .A1(n701), .A2(n632), .B1(n213), .B2(n631), .ZN(n633) );
  OAI221_X1 U724 ( .B1(n744), .B2(n634), .C1(n279), .C2(n11), .A(n633), .ZN(
        n635) );
  MUX2_X1 U725 ( .A(n636), .B(n635), .S(n210), .Z(n639) );
  NAND2_X1 U726 ( .A1(n637), .A2(n14), .ZN(n662) );
  OAI21_X1 U727 ( .B1(n338), .B2(n662), .A(n661), .ZN(n638) );
  AOI221_X1 U728 ( .B1(B[29]), .B2(n640), .C1(n690), .C2(n639), .A(n638), .ZN(
        n647) );
  NAND2_X1 U729 ( .A1(n641), .A2(n13), .ZN(n698) );
  MUX2_X1 U730 ( .A(n63), .B(n51), .S(B[29]), .Z(n642) );
  OAI21_X1 U731 ( .B1(n56), .B2(n642), .A(A[29]), .ZN(n643) );
  OAI21_X1 U732 ( .B1(n644), .B2(n698), .A(n643), .ZN(n645) );
  AOI221_X1 U733 ( .B1(N120), .B2(n5), .C1(N88), .C2(n7), .A(n645), .ZN(n646)
         );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(RES[29]) );
  OAI21_X1 U735 ( .B1(A[30]), .B2(n59), .A(n54), .ZN(n666) );
  INV_X1 U736 ( .A(n648), .ZN(n653) );
  AOI22_X1 U737 ( .A1(n213), .A2(n650), .B1(n649), .B2(n232), .ZN(n651) );
  OAI221_X1 U738 ( .B1(n10), .B2(n653), .C1(n652), .C2(n684), .A(n651), .ZN(
        n660) );
  INV_X1 U739 ( .A(n654), .ZN(n658) );
  AOI22_X1 U740 ( .A1(n701), .A2(n656), .B1(n213), .B2(n655), .ZN(n657) );
  OAI221_X1 U741 ( .B1(n744), .B2(n658), .C1(n247), .C2(n11), .A(n657), .ZN(
        n659) );
  MUX2_X1 U742 ( .A(n660), .B(n659), .S(n210), .Z(n665) );
  OAI21_X1 U743 ( .B1(n663), .B2(n662), .A(n661), .ZN(n664) );
  AOI221_X1 U744 ( .B1(B[30]), .B2(n666), .C1(n690), .C2(n665), .A(n664), .ZN(
        n672) );
  MUX2_X1 U745 ( .A(n65), .B(n51), .S(B[30]), .Z(n667) );
  OAI21_X1 U746 ( .B1(n56), .B2(n667), .A(A[30]), .ZN(n668) );
  OAI21_X1 U747 ( .B1(n669), .B2(n698), .A(n668), .ZN(n670) );
  AOI221_X1 U748 ( .B1(N121), .B2(n5), .C1(N89), .C2(n7), .A(n670), .ZN(n671)
         );
  NAND2_X1 U749 ( .A1(n672), .A2(n671), .ZN(RES[30]) );
  OAI21_X1 U750 ( .B1(A[31]), .B2(n59), .A(n54), .ZN(n691) );
  INV_X1 U751 ( .A(n673), .ZN(n678) );
  AOI22_X1 U752 ( .A1(n213), .A2(n675), .B1(n674), .B2(n232), .ZN(n676) );
  OAI221_X1 U753 ( .B1(n10), .B2(n678), .C1(n677), .C2(n684), .A(n676), .ZN(
        n688) );
  AOI211_X1 U754 ( .C1(A[28]), .C2(n46), .A(n235), .B(n679), .ZN(n686) );
  INV_X1 U755 ( .A(n680), .ZN(n685) );
  AOI22_X1 U756 ( .A1(n213), .A2(n682), .B1(n681), .B2(n232), .ZN(n683) );
  OAI221_X1 U757 ( .B1(n10), .B2(n686), .C1(n685), .C2(n684), .A(n683), .ZN(
        n687) );
  MUX2_X1 U758 ( .A(n688), .B(n687), .S(n210), .Z(n689) );
  AOI22_X1 U759 ( .A1(B[31]), .A2(n691), .B1(n690), .B2(n689), .ZN(n697) );
  MUX2_X1 U760 ( .A(n59), .B(n49), .S(B[31]), .Z(n692) );
  NAND3_X1 U761 ( .A1(n239), .A2(n55), .A3(n692), .ZN(n694) );
  AOI222_X1 U762 ( .A1(N90), .A2(n8), .B1(A[31]), .B2(n694), .C1(N122), .C2(n6), .ZN(n696) );
  OAI211_X1 U763 ( .C1(n699), .C2(n698), .A(n697), .B(n696), .ZN(RES[31]) );
  INV_X1 U764 ( .A(n412), .ZN(n732) );
  INV_X1 U765 ( .A(n407), .ZN(n725) );
  INV_X1 U766 ( .A(n269), .ZN(n731) );
  INV_X1 U767 ( .A(n265), .ZN(n724) );
  INV_X1 U768 ( .A(n700), .ZN(n254) );
  INV_X1 U769 ( .A(n211), .ZN(n730) );
  INV_X1 U770 ( .A(n204), .ZN(n723) );
  OR3_X1 U771 ( .A1(B[15]), .A2(B[14]), .A3(B[13]), .ZN(n715) );
  NOR4_X1 U772 ( .A1(n715), .A2(B[10]), .A3(B[12]), .A4(B[11]), .ZN(n722) );
  OR4_X1 U773 ( .A1(B[20]), .A2(B[19]), .A3(B[22]), .A4(B[21]), .ZN(n716) );
  NOR4_X1 U774 ( .A1(n716), .A2(B[16]), .A3(B[18]), .A4(B[17]), .ZN(n721) );
  OR4_X1 U775 ( .A1(B[27]), .A2(B[26]), .A3(B[29]), .A4(B[28]), .ZN(n717) );
  NOR4_X1 U776 ( .A1(n717), .A2(B[23]), .A3(B[25]), .A4(B[24]), .ZN(n720) );
  OR4_X1 U777 ( .A1(B[7]), .A2(B[6]), .A3(B[9]), .A4(B[8]), .ZN(n718) );
  NOR4_X1 U778 ( .A1(n718), .A2(B[30]), .A3(B[5]), .A4(B[31]), .ZN(n719) );
  NAND4_X1 U779 ( .A1(n722), .A2(n721), .A3(n720), .A4(n719), .ZN(N19) );
  INV_X2 U780 ( .A(n150), .ZN(n729) );
  INV_X2 U781 ( .A(A[11]), .ZN(n733) );
  INV_X2 U782 ( .A(A[1]), .ZN(n743) );
  INV_X2 U783 ( .A(B[1]), .ZN(n746) );
endmodule


module REG_PIPO_6_00_00_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  AOI22_X2 U3 ( .A1(DIN[0]), .A2(n20), .B1(n14), .B2(DOUT[0]), .ZN(n21) );
  AOI22_X2 U5 ( .A1(DIN[1]), .A2(n20), .B1(n14), .B2(DOUT[1]), .ZN(n19) );
  AOI22_X2 U7 ( .A1(DIN[2]), .A2(n20), .B1(n14), .B2(DOUT[2]), .ZN(n18) );
  AOI22_X2 U9 ( .A1(DIN[3]), .A2(n20), .B1(n14), .B2(DOUT[3]), .ZN(n17) );
  AOI22_X2 U11 ( .A1(DIN[4]), .A2(n20), .B1(n14), .B2(DOUT[4]), .ZN(n16) );
  AOI22_X2 U13 ( .A1(DIN[5]), .A2(n20), .B1(n14), .B2(DOUT[5]), .ZN(n15) );
  NOR2_X2 U14 ( .A1(INIT), .A2(n14), .ZN(n20) );
  INV_X2 U2 ( .A(n15), .ZN(n3) );
  INV_X2 U4 ( .A(n16), .ZN(n9) );
  INV_X2 U6 ( .A(n17), .ZN(n10) );
  INV_X2 U8 ( .A(n18), .ZN(n11) );
  INV_X2 U10 ( .A(n19), .ZN(n12) );
  INV_X2 U12 ( .A(n21), .ZN(n13) );
  INV_X2 U15 ( .A(EN), .ZN(n14) );
endmodule


module REG_PIPO_32_00000000_00000000_6 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_5 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n103), .CK(CLK), .RN(n4), .Q(DOUT[31]), .QN(
        n135) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n104), .CK(CLK), .RN(n4), .Q(DOUT[30]), .QN(
        n136) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n105), .CK(CLK), .RN(n4), .Q(DOUT[29]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n106), .CK(CLK), .RN(n4), .Q(DOUT[28]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n107), .CK(CLK), .RN(n4), .Q(DOUT[27]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n108), .CK(CLK), .RN(n4), .Q(DOUT[26]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n109), .CK(CLK), .RN(n4), .Q(DOUT[25]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n110), .CK(CLK), .RN(n4), .Q(DOUT[24]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n111), .CK(CLK), .RN(n4), .Q(DOUT[23]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n112), .CK(CLK), .RN(n4), .Q(DOUT[22]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n113), .CK(CLK), .RN(n3), .Q(DOUT[21]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n114), .CK(CLK), .RN(n3), .Q(DOUT[20]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n115), .CK(CLK), .RN(n3), .Q(DOUT[19]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n116), .CK(CLK), .RN(n3), .Q(DOUT[18]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n117), .CK(CLK), .RN(n3), .Q(DOUT[17]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n118), .CK(CLK), .RN(n3), .Q(DOUT[16]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n119), .CK(CLK), .RN(n3), .Q(DOUT[15]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n120), .CK(CLK), .RN(n3), .Q(DOUT[14]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n121), .CK(CLK), .RN(n3), .Q(DOUT[13]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n122), .CK(CLK), .RN(n3), .Q(DOUT[12]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n123), .CK(CLK), .RN(n3), .Q(DOUT[11]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n124), .CK(CLK), .RN(n2), .Q(DOUT[10]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n125), .CK(CLK), .RN(n2), .Q(DOUT[9]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n126), .CK(CLK), .RN(n2), .Q(DOUT[8]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n127), .CK(CLK), .RN(n2), .Q(DOUT[7]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n128), .CK(CLK), .RN(n2), .Q(DOUT[6]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n129), .CK(CLK), .RN(n2), .Q(DOUT[5]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n130), .CK(CLK), .RN(n2), .Q(DOUT[4]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n131), .CK(CLK), .RN(n2), .Q(DOUT[3]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n132), .CK(CLK), .RN(n2), .Q(DOUT[2]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n133), .CK(CLK), .RN(n2), .Q(DOUT[1]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n134), .CK(CLK), .RN(n2), .Q(DOUT[0]), .QN(
        n166) );
  OAI22_X2 U2 ( .A1(n166), .A2(EN), .B1(n167), .B2(n102), .ZN(n134) );
  OAI22_X2 U4 ( .A1(n165), .A2(EN), .B1(n167), .B2(n101), .ZN(n133) );
  OAI22_X2 U6 ( .A1(n164), .A2(EN), .B1(n167), .B2(n100), .ZN(n132) );
  OAI22_X2 U8 ( .A1(n163), .A2(EN), .B1(n167), .B2(n99), .ZN(n131) );
  OAI22_X2 U10 ( .A1(n162), .A2(EN), .B1(n167), .B2(n34), .ZN(n130) );
  OAI22_X2 U12 ( .A1(n161), .A2(EN), .B1(n167), .B2(n33), .ZN(n129) );
  OAI22_X2 U14 ( .A1(n160), .A2(EN), .B1(n167), .B2(n32), .ZN(n128) );
  OAI22_X2 U16 ( .A1(n159), .A2(EN), .B1(n167), .B2(n31), .ZN(n127) );
  OAI22_X2 U18 ( .A1(n158), .A2(EN), .B1(n167), .B2(n30), .ZN(n126) );
  OAI22_X2 U20 ( .A1(n157), .A2(EN), .B1(n167), .B2(n29), .ZN(n125) );
  OAI22_X2 U22 ( .A1(n156), .A2(EN), .B1(n167), .B2(n28), .ZN(n124) );
  OAI22_X2 U24 ( .A1(n155), .A2(EN), .B1(n167), .B2(n27), .ZN(n123) );
  CLKBUF_X3 U3 ( .A(RST_AN), .Z(n2) );
  CLKBUF_X3 U5 ( .A(RST_AN), .Z(n3) );
  CLKBUF_X3 U7 ( .A(RST_AN), .Z(n4) );
  INV_X1 U9 ( .A(EN), .ZN(n5) );
  OR2_X1 U11 ( .A1(INIT), .A2(n5), .ZN(n167) );
  INV_X1 U13 ( .A(n167), .ZN(n25) );
  NAND2_X1 U15 ( .A1(DIN[12]), .A2(n25), .ZN(n6) );
  OAI21_X1 U17 ( .B1(n154), .B2(EN), .A(n6), .ZN(n122) );
  NAND2_X1 U19 ( .A1(DIN[13]), .A2(n25), .ZN(n7) );
  OAI21_X1 U21 ( .B1(n153), .B2(EN), .A(n7), .ZN(n121) );
  NAND2_X1 U23 ( .A1(DIN[14]), .A2(n25), .ZN(n8) );
  OAI21_X1 U25 ( .B1(n152), .B2(EN), .A(n8), .ZN(n120) );
  NAND2_X1 U26 ( .A1(DIN[15]), .A2(n25), .ZN(n9) );
  OAI21_X1 U27 ( .B1(n151), .B2(EN), .A(n9), .ZN(n119) );
  NAND2_X1 U28 ( .A1(DIN[16]), .A2(n25), .ZN(n10) );
  OAI21_X1 U29 ( .B1(n150), .B2(EN), .A(n10), .ZN(n118) );
  NAND2_X1 U30 ( .A1(DIN[17]), .A2(n25), .ZN(n11) );
  OAI21_X1 U31 ( .B1(n149), .B2(EN), .A(n11), .ZN(n117) );
  NAND2_X1 U32 ( .A1(DIN[18]), .A2(n25), .ZN(n12) );
  OAI21_X1 U33 ( .B1(n148), .B2(EN), .A(n12), .ZN(n116) );
  NAND2_X1 U34 ( .A1(DIN[19]), .A2(n25), .ZN(n13) );
  OAI21_X1 U35 ( .B1(n147), .B2(EN), .A(n13), .ZN(n115) );
  NAND2_X1 U36 ( .A1(DIN[20]), .A2(n25), .ZN(n14) );
  OAI21_X1 U37 ( .B1(n146), .B2(EN), .A(n14), .ZN(n114) );
  NAND2_X1 U38 ( .A1(DIN[21]), .A2(n25), .ZN(n15) );
  OAI21_X1 U39 ( .B1(n145), .B2(EN), .A(n15), .ZN(n113) );
  NAND2_X1 U40 ( .A1(DIN[22]), .A2(n25), .ZN(n16) );
  OAI21_X1 U41 ( .B1(n144), .B2(EN), .A(n16), .ZN(n112) );
  NAND2_X1 U42 ( .A1(DIN[23]), .A2(n25), .ZN(n17) );
  OAI21_X1 U43 ( .B1(n143), .B2(EN), .A(n17), .ZN(n111) );
  NAND2_X1 U44 ( .A1(DIN[24]), .A2(n25), .ZN(n18) );
  OAI21_X1 U45 ( .B1(n142), .B2(EN), .A(n18), .ZN(n110) );
  NAND2_X1 U46 ( .A1(DIN[25]), .A2(n25), .ZN(n19) );
  OAI21_X1 U47 ( .B1(n141), .B2(EN), .A(n19), .ZN(n109) );
  NAND2_X1 U48 ( .A1(DIN[26]), .A2(n25), .ZN(n20) );
  OAI21_X1 U49 ( .B1(n140), .B2(EN), .A(n20), .ZN(n108) );
  NAND2_X1 U50 ( .A1(DIN[27]), .A2(n25), .ZN(n21) );
  OAI21_X1 U51 ( .B1(n139), .B2(EN), .A(n21), .ZN(n107) );
  NAND2_X1 U52 ( .A1(DIN[28]), .A2(n25), .ZN(n22) );
  OAI21_X1 U53 ( .B1(n138), .B2(EN), .A(n22), .ZN(n106) );
  NAND2_X1 U54 ( .A1(DIN[29]), .A2(n25), .ZN(n23) );
  OAI21_X1 U55 ( .B1(n137), .B2(EN), .A(n23), .ZN(n105) );
  NAND2_X1 U56 ( .A1(DIN[30]), .A2(n25), .ZN(n24) );
  OAI21_X1 U57 ( .B1(n136), .B2(EN), .A(n24), .ZN(n104) );
  NAND2_X1 U58 ( .A1(DIN[31]), .A2(n25), .ZN(n26) );
  OAI21_X1 U59 ( .B1(n135), .B2(EN), .A(n26), .ZN(n103) );
  INV_X2 U60 ( .A(DIN[11]), .ZN(n27) );
  INV_X2 U61 ( .A(DIN[10]), .ZN(n28) );
  INV_X2 U62 ( .A(DIN[9]), .ZN(n29) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n30) );
  INV_X2 U64 ( .A(DIN[7]), .ZN(n31) );
  INV_X2 U65 ( .A(DIN[6]), .ZN(n32) );
  INV_X2 U66 ( .A(DIN[5]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[4]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[3]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[2]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[1]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[0]), .ZN(n102) );
endmodule


module REG_PIPO_32_00000000_00000000_4 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_5_00_00_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  AOI22_X2 U3 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  AOI22_X2 U5 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  AOI22_X2 U7 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  AOI22_X2 U9 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  AOI22_X2 U11 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  NOR2_X2 U12 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X2 U2 ( .A(n13), .ZN(n3) );
  INV_X2 U4 ( .A(n14), .ZN(n8) );
  INV_X2 U6 ( .A(n15), .ZN(n9) );
  INV_X2 U8 ( .A(n16), .ZN(n10) );
  INV_X2 U10 ( .A(n18), .ZN(n11) );
  INV_X2 U13 ( .A(EN), .ZN(n12) );
endmodule


module REG_PIPO_1_0_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [0:0] DIN;
  output [0:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n3, n4, n2;

  DFFR_X1 \reg_mem_reg[0]  ( .D(n4), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]), .QN(
        n3) );
  NAND3_X1 U3 ( .A1(DIN[0]), .A2(n2), .A3(EN), .ZN(n1) );
  OAI21_X2 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n4) );
  INV_X2 U4 ( .A(INIT), .ZN(n2) );
endmodule


module REG_PIPO_32_00000000_00000000_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n103), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n102), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n101), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n100), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n99), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n34), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n33), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n32), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n31), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n30), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n29), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n28), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n27), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n26), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n25), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n24), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n23), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n22), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n21), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n20), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n19), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n18), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n17), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n16), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n15), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n14), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n13), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n12), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n11), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n10), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n9), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n8), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n104), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(DIN[31]), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[30]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[29]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[28]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[27]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[26]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[25]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[24]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[23]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[22]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[21]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[20]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[19]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[18]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[17]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[16]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[15]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[14]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[13]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[12]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[11]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[10]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[9]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[8]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[7]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[6]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[5]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[4]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[3]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[2]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[1]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[0]), .ZN(n103) );
  INV_X2 U73 ( .A(INIT), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n103), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n102), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n101), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n100), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n99), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n34), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n33), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n32), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n31), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n30), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n29), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n28), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n27), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n26), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n25), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n24), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n23), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n22), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n21), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n20), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n19), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n18), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n17), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n16), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n15), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n14), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n13), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n12), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n11), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n10), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n9), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n8), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n104), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(DIN[31]), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[30]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[29]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[28]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[27]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[26]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[25]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[24]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[23]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[22]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[21]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[20]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[19]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[18]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[17]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[16]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[15]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[14]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[13]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[12]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[11]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[10]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[9]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[8]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[7]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[6]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[5]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[4]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[3]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[2]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[1]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[0]), .ZN(n103) );
  INV_X2 U73 ( .A(INIT), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  OAI22_X2 U2 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  OAI22_X2 U4 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  OAI22_X2 U6 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  OAI22_X2 U8 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  OAI22_X2 U10 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  OAI22_X2 U12 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  OAI22_X2 U14 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  OAI22_X2 U16 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  OAI22_X2 U18 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  OAI22_X2 U20 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  OAI22_X2 U22 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  OAI22_X2 U24 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  OAI22_X2 U26 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  OAI22_X2 U28 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  OAI22_X2 U30 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  OAI22_X2 U32 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  OAI22_X2 U34 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  OAI22_X2 U36 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  OAI22_X2 U38 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  OAI22_X2 U40 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  OAI22_X2 U42 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  OAI22_X2 U44 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  OAI22_X2 U46 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  OAI22_X2 U48 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  OAI22_X2 U50 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  OAI22_X2 U52 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  OAI22_X2 U54 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  OAI22_X2 U56 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  OAI22_X2 U58 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  OAI22_X2 U60 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  OAI22_X2 U62 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  OAI22_X2 U64 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  NAND2_X2 U66 ( .A1(n8), .A2(EN), .ZN(n169) );
  BUF_X4 U3 ( .A(n169), .Z(n2) );
  BUF_X4 U5 ( .A(n169), .Z(n3) );
  CLKBUF_X3 U7 ( .A(n169), .Z(n4) );
  CLKBUF_X3 U9 ( .A(RST_AN), .Z(n5) );
  CLKBUF_X3 U11 ( .A(RST_AN), .Z(n6) );
  CLKBUF_X3 U13 ( .A(RST_AN), .Z(n7) );
  INV_X2 U15 ( .A(INIT), .ZN(n8) );
  INV_X2 U17 ( .A(DIN[31]), .ZN(n9) );
  INV_X2 U19 ( .A(DIN[30]), .ZN(n10) );
  INV_X2 U21 ( .A(DIN[29]), .ZN(n11) );
  INV_X2 U23 ( .A(DIN[28]), .ZN(n12) );
  INV_X2 U25 ( .A(DIN[27]), .ZN(n13) );
  INV_X2 U27 ( .A(DIN[26]), .ZN(n14) );
  INV_X2 U29 ( .A(DIN[25]), .ZN(n15) );
  INV_X2 U31 ( .A(DIN[24]), .ZN(n16) );
  INV_X2 U33 ( .A(DIN[23]), .ZN(n17) );
  INV_X2 U35 ( .A(DIN[22]), .ZN(n18) );
  INV_X2 U37 ( .A(DIN[21]), .ZN(n19) );
  INV_X2 U39 ( .A(DIN[20]), .ZN(n20) );
  INV_X2 U41 ( .A(DIN[19]), .ZN(n21) );
  INV_X2 U43 ( .A(DIN[18]), .ZN(n22) );
  INV_X2 U45 ( .A(DIN[17]), .ZN(n23) );
  INV_X2 U47 ( .A(DIN[16]), .ZN(n24) );
  INV_X2 U49 ( .A(DIN[15]), .ZN(n25) );
  INV_X2 U51 ( .A(DIN[14]), .ZN(n26) );
  INV_X2 U53 ( .A(DIN[13]), .ZN(n27) );
  INV_X2 U55 ( .A(DIN[12]), .ZN(n28) );
  INV_X2 U57 ( .A(DIN[11]), .ZN(n29) );
  INV_X2 U59 ( .A(DIN[10]), .ZN(n30) );
  INV_X2 U61 ( .A(DIN[9]), .ZN(n31) );
  INV_X2 U63 ( .A(DIN[8]), .ZN(n32) );
  INV_X2 U65 ( .A(DIN[7]), .ZN(n33) );
  INV_X2 U67 ( .A(DIN[6]), .ZN(n34) );
  INV_X2 U68 ( .A(DIN[5]), .ZN(n99) );
  INV_X2 U69 ( .A(DIN[4]), .ZN(n100) );
  INV_X2 U70 ( .A(DIN[3]), .ZN(n101) );
  INV_X2 U71 ( .A(DIN[2]), .ZN(n102) );
  INV_X2 U72 ( .A(DIN[1]), .ZN(n103) );
  INV_X2 U73 ( .A(DIN[0]), .ZN(n104) );
endmodule


module REG_PIPO_5_00_00_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  AOI22_X2 U3 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  AOI22_X2 U5 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  AOI22_X2 U7 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  AOI22_X2 U9 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  AOI22_X2 U11 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  NOR2_X2 U12 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X2 U2 ( .A(n13), .ZN(n3) );
  INV_X2 U4 ( .A(n14), .ZN(n8) );
  INV_X2 U6 ( .A(n15), .ZN(n9) );
  INV_X2 U8 ( .A(n16), .ZN(n10) );
  INV_X2 U10 ( .A(n18), .ZN(n11) );
  INV_X2 U13 ( .A(EN), .ZN(n12) );
endmodule


module DATAPATH_DW01_add_2 ( A, B, CI, SUM, CO );
  input [30:0] A;
  input [30:0] B;
  output [30:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_X2 U2 ( .A(n26), .ZN(n25) );
  INV_X2 U3 ( .A(n32), .ZN(n34) );
  INV_X2 U4 ( .A(n36), .ZN(n31) );
  INV_X2 U5 ( .A(n38), .ZN(n41) );
  NOR2_X2 U6 ( .A1(n43), .A2(n44), .ZN(n37) );
  INV_X2 U7 ( .A(n46), .ZN(n50) );
  INV_X2 U8 ( .A(n57), .ZN(n52) );
  INV_X2 U9 ( .A(n47), .ZN(n59) );
  INV_X2 U10 ( .A(n43), .ZN(n58) );
  INV_X2 U11 ( .A(n62), .ZN(n65) );
  NOR2_X2 U12 ( .A1(n67), .A2(n68), .ZN(n61) );
  INV_X2 U13 ( .A(n70), .ZN(n74) );
  INV_X2 U14 ( .A(n69), .ZN(n77) );
  INV_X2 U15 ( .A(n79), .ZN(n76) );
  INV_X2 U16 ( .A(n71), .ZN(n81) );
  INV_X2 U17 ( .A(n67), .ZN(n80) );
  INV_X2 U18 ( .A(n83), .ZN(n85) );
  NOR2_X2 U19 ( .A1(n86), .A2(n87), .ZN(n82) );
  INV_X2 U20 ( .A(n89), .ZN(n93) );
  INV_X2 U21 ( .A(n95), .ZN(n92) );
  INV_X2 U22 ( .A(n88), .ZN(n97) );
  INV_X2 U23 ( .A(n98), .ZN(n96) );
  INV_X2 U24 ( .A(n90), .ZN(n101) );
  INV_X2 U25 ( .A(n86), .ZN(n99) );
  INV_X2 U26 ( .A(n103), .ZN(n105) );
  INV_X2 U27 ( .A(n107), .ZN(n102) );
  INV_X2 U28 ( .A(n115), .ZN(n122) );
  INV_X2 U29 ( .A(n124), .ZN(n121) );
  INV_X2 U30 ( .A(n114), .ZN(n126) );
  NOR2_X2 U31 ( .A1(n127), .A2(n128), .ZN(n125) );
  INV_X2 U32 ( .A(n113), .ZN(n131) );
  NOR2_X2 U33 ( .A1(n132), .A2(n133), .ZN(n129) );
  INV_X2 U34 ( .A(n112), .ZN(n136) );
  NOR2_X2 U35 ( .A1(n137), .A2(n117), .ZN(n134) );
  INV_X2 U36 ( .A(n138), .ZN(n142) );
  NOR2_X2 U37 ( .A1(n144), .A2(n145), .ZN(n143) );
  NOR2_X2 U38 ( .A1(n3), .A2(n1), .ZN(n149) );
  INV_X2 U39 ( .A(n6), .ZN(n4) );
  NOR2_X2 U40 ( .A1(n20), .A2(n120), .ZN(n5) );
  NOR2_X2 U41 ( .A1(n19), .A2(n20), .ZN(n17) );
  INV_X2 U42 ( .A(n21), .ZN(n22) );
  NOR2_X2 U43 ( .A1(n14), .A2(n15), .ZN(n11) );
  INV_X2 U44 ( .A(n16), .ZN(n18) );
  INV_X2 U45 ( .A(n10), .ZN(n7) );
  INV_X2 U46 ( .A(n12), .ZN(n13) );
  INV_X2 U47 ( .A(n9), .ZN(n8) );
  INV_X2 U48 ( .A(n155), .ZN(n23) );
  INV_X2 U49 ( .A(n26), .ZN(n33) );
  INV_X2 U50 ( .A(n27), .ZN(n24) );
  NOR2_X2 U51 ( .A1(n26), .A2(n156), .ZN(n119) );
  INV_X2 U52 ( .A(A[2]), .ZN(n26) );
  INV_X2 U53 ( .A(n35), .ZN(n32) );
  INV_X2 U54 ( .A(n157), .ZN(n27) );
  INV_X2 U55 ( .A(n154), .ZN(n21) );
  INV_X2 U56 ( .A(n153), .ZN(n16) );
  INV_X2 U57 ( .A(n152), .ZN(n12) );
  INV_X2 U58 ( .A(n151), .ZN(n9) );
  INV_X2 U59 ( .A(n150), .ZN(n6) );
  INV_X2 U60 ( .A(n148), .ZN(n139) );
  INV_X2 U61 ( .A(n146), .ZN(n138) );
  INV_X2 U62 ( .A(n141), .ZN(n112) );
  INV_X2 U63 ( .A(n135), .ZN(n113) );
  INV_X2 U64 ( .A(n130), .ZN(n114) );
  INV_X2 U65 ( .A(n123), .ZN(n115) );
  INV_X2 U66 ( .A(n158), .ZN(n140) );
  INV_X2 U67 ( .A(n106), .ZN(n103) );
  INV_X2 U68 ( .A(n104), .ZN(n90) );
  INV_X2 U69 ( .A(n100), .ZN(n88) );
  INV_X2 U70 ( .A(n94), .ZN(n89) );
  INV_X2 U71 ( .A(n91), .ZN(n83) );
  INV_X2 U72 ( .A(n84), .ZN(n71) );
  INV_X2 U73 ( .A(n78), .ZN(n69) );
  INV_X2 U74 ( .A(n75), .ZN(n70) );
  INV_X2 U75 ( .A(n66), .ZN(n62) );
  INV_X2 U76 ( .A(n60), .ZN(n47) );
  INV_X2 U77 ( .A(n56), .ZN(n45) );
  INV_X2 U78 ( .A(n51), .ZN(n46) );
  INV_X2 U79 ( .A(n42), .ZN(n38) );
  NAND2_X2 U80 ( .A1(n31), .A2(n32), .ZN(n28) );
  NAND2_X2 U81 ( .A1(n45), .A2(n52), .ZN(n48) );
  INV_X2 U82 ( .A(n55), .ZN(n54) );
  NAND2_X2 U83 ( .A1(n69), .A2(n76), .ZN(n72) );
  NAND2_X2 U84 ( .A1(n108), .A2(n109), .ZN(n107) );
  INV_X2 U85 ( .A(n145), .ZN(n147) );
  INV_X2 U86 ( .A(n3), .ZN(n2) );
  NAND2_X2 U87 ( .A1(n118), .A2(n119), .ZN(n116) );
  INV_X2 U88 ( .A(n33), .ZN(SUM[2]) );
  INV_X2 U89 ( .A(A[30]), .ZN(n30) );
  XNOR2_X1 U90 ( .A(n1), .B(n2), .ZN(SUM[9]) );
  XNOR2_X1 U91 ( .A(n4), .B(n5), .ZN(SUM[8]) );
  XNOR2_X2 U92 ( .A(n7), .B(n8), .ZN(SUM[7]) );
  NAND2_X2 U93 ( .A1(n11), .A2(n12), .ZN(n10) );
  XNOR2_X2 U94 ( .A(n13), .B(n11), .ZN(SUM[6]) );
  INV_X1 U95 ( .A(n16), .ZN(n15) );
  INV_X1 U96 ( .A(n17), .ZN(n14) );
  XNOR2_X1 U97 ( .A(n18), .B(n17), .ZN(SUM[5]) );
  INV_X1 U98 ( .A(n21), .ZN(n19) );
  XNOR2_X2 U99 ( .A(n22), .B(n23), .ZN(SUM[4]) );
  XNOR2_X2 U100 ( .A(n24), .B(n25), .ZN(SUM[3]) );
  XNOR2_X2 U101 ( .A(n28), .B(n29), .ZN(SUM[30]) );
  INV_X2 U102 ( .A(n30), .ZN(n29) );
  XNOR2_X2 U103 ( .A(n31), .B(n34), .ZN(SUM[29]) );
  INV_X2 U104 ( .A(A[29]), .ZN(n35) );
  NAND2_X1 U105 ( .A1(n37), .A2(n38), .ZN(n36) );
  XNOR2_X2 U106 ( .A(n39), .B(n40), .ZN(SUM[28]) );
  INV_X1 U107 ( .A(n41), .ZN(n40) );
  INV_X2 U108 ( .A(A[28]), .ZN(n42) );
  INV_X1 U109 ( .A(n37), .ZN(n39) );
  NAND3_X1 U110 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n44) );
  XNOR2_X2 U111 ( .A(n48), .B(n49), .ZN(SUM[27]) );
  INV_X1 U112 ( .A(n50), .ZN(n49) );
  INV_X2 U113 ( .A(A[27]), .ZN(n51) );
  XNOR2_X2 U114 ( .A(n53), .B(n54), .ZN(SUM[26]) );
  INV_X1 U115 ( .A(n45), .ZN(n55) );
  INV_X2 U116 ( .A(A[26]), .ZN(n56) );
  INV_X1 U117 ( .A(n52), .ZN(n53) );
  NAND2_X2 U118 ( .A1(n47), .A2(n58), .ZN(n57) );
  XNOR2_X2 U119 ( .A(n58), .B(n59), .ZN(SUM[25]) );
  INV_X2 U120 ( .A(A[25]), .ZN(n60) );
  NAND2_X2 U121 ( .A1(n61), .A2(n62), .ZN(n43) );
  XNOR2_X2 U122 ( .A(n63), .B(n64), .ZN(SUM[24]) );
  INV_X1 U123 ( .A(n65), .ZN(n64) );
  INV_X2 U124 ( .A(A[24]), .ZN(n66) );
  INV_X1 U125 ( .A(n61), .ZN(n63) );
  NAND3_X1 U126 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n68) );
  XNOR2_X2 U127 ( .A(n72), .B(n73), .ZN(SUM[23]) );
  INV_X1 U128 ( .A(n74), .ZN(n73) );
  INV_X2 U129 ( .A(A[23]), .ZN(n75) );
  XNOR2_X2 U130 ( .A(n76), .B(n77), .ZN(SUM[22]) );
  INV_X2 U131 ( .A(A[22]), .ZN(n78) );
  NAND2_X2 U132 ( .A1(n71), .A2(n80), .ZN(n79) );
  XNOR2_X2 U133 ( .A(n81), .B(n80), .ZN(SUM[21]) );
  NAND2_X2 U134 ( .A1(n82), .A2(n83), .ZN(n67) );
  INV_X2 U135 ( .A(A[21]), .ZN(n84) );
  XNOR2_X1 U136 ( .A(n85), .B(n82), .ZN(SUM[20]) );
  NAND3_X1 U137 ( .A1(n88), .A2(n89), .A3(n90), .ZN(n87) );
  INV_X2 U138 ( .A(A[20]), .ZN(n91) );
  XNOR2_X2 U139 ( .A(n92), .B(n93), .ZN(SUM[19]) );
  INV_X2 U140 ( .A(A[19]), .ZN(n94) );
  NAND2_X2 U141 ( .A1(n96), .A2(n88), .ZN(n95) );
  XNOR2_X2 U142 ( .A(n97), .B(n96), .ZN(SUM[18]) );
  NAND2_X2 U143 ( .A1(n90), .A2(n99), .ZN(n98) );
  INV_X2 U144 ( .A(A[18]), .ZN(n100) );
  XNOR2_X2 U145 ( .A(n101), .B(n99), .ZN(SUM[17]) );
  NAND2_X2 U146 ( .A1(n102), .A2(n103), .ZN(n86) );
  INV_X2 U147 ( .A(A[17]), .ZN(n104) );
  XNOR2_X2 U148 ( .A(n102), .B(n105), .ZN(SUM[16]) );
  INV_X2 U149 ( .A(A[16]), .ZN(n106) );
  NOR2_X2 U150 ( .A1(n110), .A2(n111), .ZN(n109) );
  NAND2_X2 U151 ( .A1(n112), .A2(n113), .ZN(n111) );
  NAND2_X2 U152 ( .A1(n114), .A2(n115), .ZN(n110) );
  NOR2_X2 U153 ( .A1(n116), .A2(n117), .ZN(n108) );
  INV_X1 U154 ( .A(n120), .ZN(n118) );
  XNOR2_X2 U155 ( .A(n121), .B(n122), .ZN(SUM[15]) );
  INV_X2 U156 ( .A(A[15]), .ZN(n123) );
  NAND2_X2 U157 ( .A1(n125), .A2(n114), .ZN(n124) );
  XNOR2_X2 U158 ( .A(n126), .B(n125), .ZN(SUM[14]) );
  INV_X1 U159 ( .A(n113), .ZN(n128) );
  INV_X1 U160 ( .A(n129), .ZN(n127) );
  INV_X2 U161 ( .A(A[14]), .ZN(n130) );
  XNOR2_X1 U162 ( .A(n131), .B(n129), .ZN(SUM[13]) );
  INV_X1 U163 ( .A(n134), .ZN(n133) );
  INV_X1 U164 ( .A(n112), .ZN(n132) );
  INV_X2 U165 ( .A(A[13]), .ZN(n135) );
  XNOR2_X2 U166 ( .A(n136), .B(n134), .ZN(SUM[12]) );
  NAND4_X2 U167 ( .A1(n138), .A2(n139), .A3(n140), .A4(n6), .ZN(n117) );
  INV_X1 U168 ( .A(n5), .ZN(n137) );
  INV_X2 U169 ( .A(A[12]), .ZN(n141) );
  XNOR2_X1 U170 ( .A(n142), .B(n143), .ZN(SUM[11]) );
  INV_X2 U171 ( .A(A[11]), .ZN(n146) );
  XNOR2_X1 U172 ( .A(n144), .B(n147), .ZN(SUM[10]) );
  INV_X1 U173 ( .A(n139), .ZN(n145) );
  INV_X2 U174 ( .A(A[10]), .ZN(n148) );
  INV_X1 U175 ( .A(n149), .ZN(n144) );
  NAND2_X2 U176 ( .A1(n5), .A2(n6), .ZN(n1) );
  INV_X2 U177 ( .A(A[8]), .ZN(n150) );
  NAND4_X2 U178 ( .A1(n21), .A2(n16), .A3(n12), .A4(n9), .ZN(n120) );
  INV_X2 U179 ( .A(A[7]), .ZN(n151) );
  INV_X2 U180 ( .A(A[6]), .ZN(n152) );
  INV_X2 U181 ( .A(A[5]), .ZN(n153) );
  INV_X2 U182 ( .A(A[4]), .ZN(n154) );
  INV_X1 U183 ( .A(n23), .ZN(n20) );
  INV_X1 U184 ( .A(n119), .ZN(n155) );
  INV_X1 U185 ( .A(n27), .ZN(n156) );
  INV_X2 U186 ( .A(A[3]), .ZN(n157) );
  INV_X1 U187 ( .A(n140), .ZN(n3) );
  INV_X2 U188 ( .A(A[9]), .ZN(n158) );
endmodule


module DATAPATH ( CLK, RST_AN, .CTRL_WORD({\CTRL_WORD[J_TYPE_IMM_SEL] , 
        \CTRL_WORD[R_TYPE_SEL] , \CTRL_WORD[IMM_SEL] , 
        \CTRL_WORD[PC_PLS_4_SEL] , \CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] , \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }), INSTR_CU, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .DP_SIG({
        \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] , 
        \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] , 
        \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] , 
        \DP_SIG[INSTR_OPCODE_M][0] }), IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] INSTR_CU;
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN, \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] , \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  wire   \npc_f[31] , n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n184, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n277, n278, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n291, n302, n1,
         n2, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n183;
  wire   [30:0] pc_pls_4_f;
  wire   [31:0] pc_pls_4_d;
  wire   [31:0] instr_d;
  wire   [4:0] rf_waddr_d;
  wire   [31:0] rf_dout1_d;
  wire   [31:0] rf_dout2_d;
  wire   [4:0] rf_waddr_wb;
  wire   [31:16] imm_d;
  wire   [5:0] instr_opcode_e;
  wire   [31:0] pc_pls_4_e;
  wire   [31:0] rf_dout1_e;
  wire   [31:0] rf_dout2_e;
  wire   [31:0] imm_e;
  wire   [4:0] rs2_e;
  wire   [4:0] rs3_e;
  wire   [31:0] alu_a_e;
  wire   [31:0] alu_out_e;
  wire   [31:0] pc_pls_4_m;
  wire   [4:0] rf_waddr_m;
  wire   [31:0] pc_pls_4_wb;
  wire   [31:0] alu_out_wb;
  wire   [31:0] dmem_dout_wb;
  assign INSTR_CU[31] = IMEM_DOUT[31];
  assign INSTR_CU[30] = IMEM_DOUT[30];
  assign INSTR_CU[29] = IMEM_DOUT[29];
  assign INSTR_CU[28] = IMEM_DOUT[28];
  assign INSTR_CU[27] = IMEM_DOUT[27];
  assign INSTR_CU[26] = IMEM_DOUT[26];
  assign INSTR_CU[25] = IMEM_DOUT[25];
  assign INSTR_CU[24] = IMEM_DOUT[24];
  assign INSTR_CU[23] = IMEM_DOUT[23];
  assign INSTR_CU[22] = IMEM_DOUT[22];
  assign INSTR_CU[21] = IMEM_DOUT[21];
  assign INSTR_CU[20] = IMEM_DOUT[20];
  assign INSTR_CU[19] = IMEM_DOUT[19];
  assign INSTR_CU[18] = IMEM_DOUT[18];
  assign INSTR_CU[17] = IMEM_DOUT[17];
  assign INSTR_CU[16] = IMEM_DOUT[16];
  assign INSTR_CU[15] = IMEM_DOUT[15];
  assign INSTR_CU[14] = IMEM_DOUT[14];
  assign INSTR_CU[13] = IMEM_DOUT[13];
  assign INSTR_CU[12] = IMEM_DOUT[12];
  assign INSTR_CU[11] = IMEM_DOUT[11];
  assign INSTR_CU[10] = IMEM_DOUT[10];
  assign INSTR_CU[9] = IMEM_DOUT[9];
  assign INSTR_CU[8] = IMEM_DOUT[8];
  assign INSTR_CU[7] = IMEM_DOUT[7];
  assign INSTR_CU[6] = IMEM_DOUT[6];
  assign INSTR_CU[5] = IMEM_DOUT[5];
  assign INSTR_CU[4] = IMEM_DOUT[4];
  assign INSTR_CU[3] = IMEM_DOUT[3];
  assign INSTR_CU[2] = IMEM_DOUT[2];
  assign INSTR_CU[1] = IMEM_DOUT[1];
  assign INSTR_CU[0] = IMEM_DOUT[0];

  AOI22_X2 U7 ( .A1(rs2_e[4]), .A2(n143), .B1(rs3_e[4]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n144) );
  AOI22_X2 U8 ( .A1(rs2_e[3]), .A2(n143), .B1(rs3_e[3]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n145) );
  AOI22_X2 U9 ( .A1(rs2_e[2]), .A2(n143), .B1(rs3_e[2]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n146) );
  AOI22_X2 U10 ( .A1(rs2_e[1]), .A2(n143), .B1(rs3_e[1]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n147) );
  AOI22_X2 U11 ( .A1(rs2_e[0]), .A2(n143), .B1(rs3_e[0]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n148) );
  OR2_X2 U12 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[4]), .ZN(
        rf_waddr_d[4]) );
  OR2_X2 U13 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[3]), .ZN(
        rf_waddr_d[3]) );
  OR2_X2 U14 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[2]), .ZN(
        rf_waddr_d[2]) );
  OR2_X2 U15 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[1]), .ZN(
        rf_waddr_d[1]) );
  OR2_X2 U16 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[0]), .ZN(
        rf_waddr_d[0]) );
  AOI222_X2 U17 ( .A1(dmem_dout_wb[9]), .A2(n15), .B1(alu_out_wb[9]), .B2(n12), 
        .C1(pc_pls_4_wb[9]), .C2(n9), .ZN(n149) );
  AOI222_X2 U18 ( .A1(dmem_dout_wb[8]), .A2(n15), .B1(alu_out_wb[8]), .B2(n12), 
        .C1(pc_pls_4_wb[8]), .C2(n9), .ZN(n152) );
  AOI222_X2 U19 ( .A1(dmem_dout_wb[7]), .A2(n15), .B1(alu_out_wb[7]), .B2(n12), 
        .C1(pc_pls_4_wb[7]), .C2(n9), .ZN(n153) );
  AOI222_X2 U20 ( .A1(dmem_dout_wb[6]), .A2(n15), .B1(alu_out_wb[6]), .B2(n12), 
        .C1(pc_pls_4_wb[6]), .C2(n9), .ZN(n154) );
  AOI222_X2 U21 ( .A1(dmem_dout_wb[5]), .A2(n15), .B1(alu_out_wb[5]), .B2(n12), 
        .C1(pc_pls_4_wb[5]), .C2(n9), .ZN(n155) );
  AOI222_X2 U22 ( .A1(dmem_dout_wb[4]), .A2(n15), .B1(alu_out_wb[4]), .B2(n12), 
        .C1(pc_pls_4_wb[4]), .C2(n9), .ZN(n156) );
  AOI222_X2 U23 ( .A1(dmem_dout_wb[3]), .A2(n15), .B1(alu_out_wb[3]), .B2(n12), 
        .C1(pc_pls_4_wb[3]), .C2(n9), .ZN(n157) );
  AOI222_X2 U24 ( .A1(dmem_dout_wb[31]), .A2(n15), .B1(alu_out_wb[31]), .B2(
        n12), .C1(pc_pls_4_wb[31]), .C2(n9), .ZN(n158) );
  AOI222_X2 U25 ( .A1(dmem_dout_wb[30]), .A2(n15), .B1(alu_out_wb[30]), .B2(
        n11), .C1(pc_pls_4_wb[30]), .C2(n8), .ZN(n159) );
  AOI222_X2 U26 ( .A1(dmem_dout_wb[2]), .A2(n15), .B1(alu_out_wb[2]), .B2(n11), 
        .C1(pc_pls_4_wb[2]), .C2(n8), .ZN(n160) );
  AOI222_X2 U27 ( .A1(dmem_dout_wb[29]), .A2(n14), .B1(alu_out_wb[29]), .B2(
        n11), .C1(pc_pls_4_wb[29]), .C2(n8), .ZN(n161) );
  AOI222_X2 U28 ( .A1(dmem_dout_wb[28]), .A2(n14), .B1(alu_out_wb[28]), .B2(
        n11), .C1(pc_pls_4_wb[28]), .C2(n8), .ZN(n162) );
  AOI222_X2 U29 ( .A1(dmem_dout_wb[27]), .A2(n14), .B1(alu_out_wb[27]), .B2(
        n11), .C1(pc_pls_4_wb[27]), .C2(n8), .ZN(n163) );
  AOI222_X2 U30 ( .A1(dmem_dout_wb[26]), .A2(n14), .B1(alu_out_wb[26]), .B2(
        n11), .C1(pc_pls_4_wb[26]), .C2(n8), .ZN(n164) );
  AOI222_X2 U31 ( .A1(dmem_dout_wb[25]), .A2(n14), .B1(alu_out_wb[25]), .B2(
        n11), .C1(pc_pls_4_wb[25]), .C2(n8), .ZN(n165) );
  AOI222_X2 U32 ( .A1(dmem_dout_wb[24]), .A2(n14), .B1(alu_out_wb[24]), .B2(
        n11), .C1(pc_pls_4_wb[24]), .C2(n8), .ZN(n166) );
  AOI222_X2 U33 ( .A1(dmem_dout_wb[23]), .A2(n14), .B1(alu_out_wb[23]), .B2(
        n11), .C1(pc_pls_4_wb[23]), .C2(n8), .ZN(n167) );
  AOI222_X2 U34 ( .A1(dmem_dout_wb[22]), .A2(n14), .B1(alu_out_wb[22]), .B2(
        n11), .C1(pc_pls_4_wb[22]), .C2(n8), .ZN(n168) );
  AOI222_X2 U35 ( .A1(dmem_dout_wb[21]), .A2(n14), .B1(alu_out_wb[21]), .B2(
        n11), .C1(pc_pls_4_wb[21]), .C2(n8), .ZN(n169) );
  AOI222_X2 U36 ( .A1(dmem_dout_wb[20]), .A2(n14), .B1(alu_out_wb[20]), .B2(
        n11), .C1(pc_pls_4_wb[20]), .C2(n8), .ZN(n170) );
  AOI222_X2 U37 ( .A1(dmem_dout_wb[1]), .A2(n14), .B1(alu_out_wb[1]), .B2(n10), 
        .C1(pc_pls_4_wb[1]), .C2(n7), .ZN(n171) );
  AOI222_X2 U38 ( .A1(dmem_dout_wb[19]), .A2(n14), .B1(alu_out_wb[19]), .B2(
        n10), .C1(pc_pls_4_wb[19]), .C2(n7), .ZN(n172) );
  AOI222_X2 U39 ( .A1(dmem_dout_wb[18]), .A2(n13), .B1(alu_out_wb[18]), .B2(
        n10), .C1(pc_pls_4_wb[18]), .C2(n7), .ZN(n173) );
  AOI222_X2 U40 ( .A1(dmem_dout_wb[17]), .A2(n13), .B1(alu_out_wb[17]), .B2(
        n10), .C1(pc_pls_4_wb[17]), .C2(n7), .ZN(n174) );
  AOI222_X2 U41 ( .A1(dmem_dout_wb[16]), .A2(n13), .B1(alu_out_wb[16]), .B2(
        n10), .C1(pc_pls_4_wb[16]), .C2(n7), .ZN(n175) );
  AOI222_X2 U42 ( .A1(dmem_dout_wb[15]), .A2(n13), .B1(alu_out_wb[15]), .B2(
        n10), .C1(pc_pls_4_wb[15]), .C2(n7), .ZN(n176) );
  AOI222_X2 U43 ( .A1(dmem_dout_wb[14]), .A2(n13), .B1(alu_out_wb[14]), .B2(
        n10), .C1(pc_pls_4_wb[14]), .C2(n7), .ZN(n177) );
  AOI222_X2 U44 ( .A1(dmem_dout_wb[13]), .A2(n13), .B1(alu_out_wb[13]), .B2(
        n10), .C1(pc_pls_4_wb[13]), .C2(n7), .ZN(n178) );
  AOI222_X2 U45 ( .A1(dmem_dout_wb[12]), .A2(n13), .B1(alu_out_wb[12]), .B2(
        n10), .C1(pc_pls_4_wb[12]), .C2(n7), .ZN(n179) );
  AOI222_X2 U46 ( .A1(dmem_dout_wb[11]), .A2(n13), .B1(alu_out_wb[11]), .B2(
        n10), .C1(pc_pls_4_wb[11]), .C2(n7), .ZN(n180) );
  AOI222_X2 U47 ( .A1(dmem_dout_wb[10]), .A2(n13), .B1(alu_out_wb[10]), .B2(
        n10), .C1(pc_pls_4_wb[10]), .C2(n7), .ZN(n181) );
  AOI222_X2 U48 ( .A1(dmem_dout_wb[0]), .A2(n13), .B1(alu_out_wb[0]), .B2(n10), 
        .C1(pc_pls_4_wb[0]), .C2(n7), .ZN(n182) );
  NOR2_X2 U49 ( .A1(n183), .A2(n13), .ZN(n151) );
  NOR2_X2 U50 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(n13), .ZN(n150) );
  AND2_X2 U58 ( .A1(DMEM_RWADDR[31]), .A2(n184), .ZN(\npc_f[31] ) );
  NOR2_X2 U86 ( .A1(n217), .A2(n218), .ZN(n302) );
  NAND4_X2 U87 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(n218) );
  NOR4_X2 U88 ( .A1(rf_dout1_e[23]), .A2(rf_dout1_e[22]), .A3(rf_dout1_e[21]), 
        .A4(rf_dout1_e[20]), .ZN(n222) );
  NOR4_X2 U89 ( .A1(rf_dout1_e[1]), .A2(rf_dout1_e[19]), .A3(rf_dout1_e[18]), 
        .A4(rf_dout1_e[17]), .ZN(n221) );
  NOR4_X2 U90 ( .A1(rf_dout1_e[16]), .A2(rf_dout1_e[15]), .A3(rf_dout1_e[14]), 
        .A4(rf_dout1_e[13]), .ZN(n220) );
  NOR4_X2 U91 ( .A1(rf_dout1_e[12]), .A2(rf_dout1_e[11]), .A3(rf_dout1_e[10]), 
        .A4(rf_dout1_e[0]), .ZN(n219) );
  NAND4_X2 U92 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(n217) );
  NOR4_X2 U93 ( .A1(rf_dout1_e[9]), .A2(rf_dout1_e[8]), .A3(rf_dout1_e[7]), 
        .A4(rf_dout1_e[6]), .ZN(n226) );
  NOR4_X2 U94 ( .A1(rf_dout1_e[5]), .A2(rf_dout1_e[4]), .A3(rf_dout1_e[3]), 
        .A4(rf_dout1_e[31]), .ZN(n225) );
  NOR4_X2 U95 ( .A1(rf_dout1_e[30]), .A2(rf_dout1_e[2]), .A3(rf_dout1_e[29]), 
        .A4(rf_dout1_e[28]), .ZN(n224) );
  NOR4_X2 U96 ( .A1(rf_dout1_e[27]), .A2(rf_dout1_e[26]), .A3(rf_dout1_e[25]), 
        .A4(rf_dout1_e[24]), .ZN(n223) );
  NAND2_X2 U97 ( .A1(n227), .A2(n228), .ZN(imm_d[31]) );
  NAND2_X2 U98 ( .A1(instr_d[25]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n228)
         );
  NAND2_X2 U99 ( .A1(n227), .A2(n229), .ZN(imm_d[24]) );
  NAND2_X2 U100 ( .A1(instr_d[24]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n229) );
  NAND2_X2 U101 ( .A1(n227), .A2(n230), .ZN(imm_d[23]) );
  NAND2_X2 U102 ( .A1(instr_d[23]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n230) );
  NAND2_X2 U103 ( .A1(n227), .A2(n231), .ZN(imm_d[22]) );
  NAND2_X2 U104 ( .A1(instr_d[22]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n231) );
  NAND2_X2 U105 ( .A1(n227), .A2(n232), .ZN(imm_d[21]) );
  NAND2_X2 U106 ( .A1(instr_d[21]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n232) );
  NAND2_X2 U107 ( .A1(n227), .A2(n233), .ZN(imm_d[20]) );
  NAND2_X2 U108 ( .A1(instr_d[20]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n233) );
  NAND2_X2 U109 ( .A1(n227), .A2(n234), .ZN(imm_d[19]) );
  NAND2_X2 U110 ( .A1(instr_d[19]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n234) );
  NAND2_X2 U111 ( .A1(n227), .A2(n235), .ZN(imm_d[18]) );
  NAND2_X2 U112 ( .A1(instr_d[18]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n235) );
  NAND2_X2 U113 ( .A1(n227), .A2(n236), .ZN(imm_d[17]) );
  NAND2_X2 U114 ( .A1(instr_d[17]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n236) );
  NAND2_X2 U115 ( .A1(n227), .A2(n237), .ZN(imm_d[16]) );
  NAND2_X2 U116 ( .A1(instr_d[16]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n237) );
  NAND2_X2 U117 ( .A1(instr_d[15]), .A2(n142), .ZN(n227) );
  OAI21_X2 U164 ( .B1(n20), .B2(n64), .A(n277), .ZN(alu_a_e[31]) );
  NAND2_X2 U165 ( .A1(pc_pls_4_e[31]), .A2(n18), .ZN(n277) );
  OAI21_X2 U166 ( .B1(n19), .B2(n65), .A(n278), .ZN(alu_a_e[30]) );
  NAND2_X2 U167 ( .A1(pc_pls_4_e[30]), .A2(n18), .ZN(n278) );
  OAI21_X2 U170 ( .B1(n19), .B2(n66), .A(n280), .ZN(alu_a_e[29]) );
  NAND2_X2 U171 ( .A1(pc_pls_4_e[29]), .A2(n18), .ZN(n280) );
  OAI21_X2 U172 ( .B1(n19), .B2(n67), .A(n281), .ZN(alu_a_e[28]) );
  NAND2_X2 U173 ( .A1(pc_pls_4_e[28]), .A2(n18), .ZN(n281) );
  OAI21_X2 U174 ( .B1(n19), .B2(n68), .A(n282), .ZN(alu_a_e[27]) );
  NAND2_X2 U175 ( .A1(pc_pls_4_e[27]), .A2(n18), .ZN(n282) );
  OAI21_X2 U176 ( .B1(n19), .B2(n69), .A(n283), .ZN(alu_a_e[26]) );
  NAND2_X2 U177 ( .A1(pc_pls_4_e[26]), .A2(n18), .ZN(n283) );
  OAI21_X2 U178 ( .B1(n19), .B2(n70), .A(n284), .ZN(alu_a_e[25]) );
  NAND2_X2 U179 ( .A1(pc_pls_4_e[25]), .A2(n18), .ZN(n284) );
  OAI21_X2 U180 ( .B1(n19), .B2(n71), .A(n285), .ZN(alu_a_e[24]) );
  NAND2_X2 U181 ( .A1(pc_pls_4_e[24]), .A2(n18), .ZN(n285) );
  OAI21_X2 U182 ( .B1(n19), .B2(n72), .A(n286), .ZN(alu_a_e[23]) );
  NAND2_X2 U183 ( .A1(pc_pls_4_e[23]), .A2(n18), .ZN(n286) );
  OAI21_X2 U184 ( .B1(n19), .B2(n73), .A(n287), .ZN(alu_a_e[22]) );
  NAND2_X2 U185 ( .A1(pc_pls_4_e[22]), .A2(n18), .ZN(n287) );
  OAI21_X2 U186 ( .B1(n19), .B2(n74), .A(n288), .ZN(alu_a_e[21]) );
  NAND2_X2 U187 ( .A1(pc_pls_4_e[21]), .A2(n19), .ZN(n288) );
  OAI21_X2 U188 ( .B1(n19), .B2(n75), .A(n289), .ZN(alu_a_e[20]) );
  NAND2_X2 U189 ( .A1(pc_pls_4_e[20]), .A2(n18), .ZN(n289) );
  OAI21_X2 U192 ( .B1(n20), .B2(n76), .A(n291), .ZN(alu_a_e[19]) );
  NAND2_X2 U193 ( .A1(pc_pls_4_e[19]), .A2(n18), .ZN(n291) );
  REG_PIPO_32_fffffffc_fffffffc U_PC_REG ( .CLK(CLK), .RST_AN(n26), .EN(1'b1), 
        .INIT(1'b0), .DIN({\npc_f[31] , n29, n30, n31, n32, n33, n34, n35, n36, 
        n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
        n51, n52, n53, n54, n55, n56, n57, n58, n109}), .DOUT(IMEM_ADDR) );
  REG_PIPO_32_00000000_00000000_0 U_PC_PLS_4_REG_FD ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN({1'b0, pc_pls_4_f}), 
        .DOUT(pc_pls_4_d) );
  REG_PIPO_32_00000000_00000000_11 U_INSTR_REG_FD ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN(IMEM_DOUT), .DOUT(instr_d) );
  RF_ADDR_W5_DATA_W32 U_RF ( .CLK(CLK), .RST_AN(n25), .ENABLE(1'b1), .RD1(1'b1), .RD2(1'b1), .WR(\CTRL_WORD[RF_WEN] ), .ADD_WR(rf_waddr_d), .ADD_RD1(
        instr_d[25:21]), .ADD_RD2(instr_d[20:16]), .DATAIN({n110, n111, n112, 
        n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
        n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
        n137, n138, n139, n140, n141}), .OUT1(rf_dout1_d), .OUT2(rf_dout2_d)
         );
  REG_PIPO_6_00_00_0 U_INSTR_OPCODE_REG_DE ( .CLK(CLK), .RST_AN(n25), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[31:26]), .DOUT(instr_opcode_e) );
  REG_PIPO_32_00000000_00000000_10 U_PC_PLS_4_REG_DE ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(pc_pls_4_d), .DOUT(
        pc_pls_4_e) );
  REG_PIPO_32_00000000_00000000_9 U_RF_DOUT1_REG_DE ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout1_d), .DOUT(
        rf_dout1_e) );
  REG_PIPO_32_00000000_00000000_8 U_RF_DOUT2_REG_DE ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout2_d), .DOUT(
        rf_dout2_e) );
  REG_PIPO_32_00000000_00000000_7 U_IMM_REG_DE ( .CLK(CLK), .RST_AN(n26), .EN(
        1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN({imm_d[31], imm_d[31], 
        imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[24:16], 
        instr_d[15:0]}), .DOUT(imm_e) );
  REG_PIPO_5_00_00_0 U_RS2_REG_DE ( .CLK(CLK), .RST_AN(n25), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[20:16]), .DOUT(rs2_e) );
  REG_PIPO_5_00_00_3 U_RS3_REG_DE ( .CLK(CLK), .RST_AN(n25), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[15:11]), .DOUT(rs3_e) );
  ALU_DATA_W32 U_ALU ( .FUNC({\CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] }), .A(alu_a_e), .B({n77, n78, n79, n80, n81, 
        n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
        n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
        n108}), .RES(alu_out_e) );
  REG_PIPO_6_00_00_1 U_INSTR_OPCODE_REG_EM ( .CLK(CLK), .RST_AN(n25), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(instr_opcode_e), .DOUT({
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }) );
  REG_PIPO_32_00000000_00000000_6 U_PC_PLS_4_REG_EM ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(pc_pls_4_e), .DOUT(
        pc_pls_4_m) );
  REG_PIPO_32_00000000_00000000_5 U_ALU_OUT_REG_EM ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(alu_out_e), .DOUT(
        DMEM_RWADDR) );
  REG_PIPO_32_00000000_00000000_4 U_DMEM_DOUT_REG_EM ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(rf_dout2_e), .DOUT(
        DMEM_DIN) );
  REG_PIPO_5_00_00_2 U_RF_WADDR_REG_EM ( .CLK(CLK), .RST_AN(n25), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN({n59, n60, n61, n62, n63}), .DOUT(
        rf_waddr_m) );
  REG_PIPO_1_0_0 U_IS_0_REG_EM ( .CLK(CLK), .RST_AN(n26), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_EM] ), .DIN(n302), .DOUT(\DP_SIG[CMPR_0_IS_0_M] ) );
  REG_PIPO_32_00000000_00000000_3 U_PC_PLS_4_REG_MWB ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(pc_pls_4_m), .DOUT(
        pc_pls_4_wb) );
  REG_PIPO_32_00000000_00000000_2 U_ALU_OUT_REG_MWB ( .CLK(CLK), .RST_AN(n26), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_RWADDR), .DOUT(
        alu_out_wb) );
  REG_PIPO_32_00000000_00000000_1 U_DMEM_DOUT_REG_MWB ( .CLK(CLK), .RST_AN(n26), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_DOUT), .DOUT(dmem_dout_wb) );
  REG_PIPO_5_00_00_1 U_RF_WADDR_REG_MWB ( .CLK(CLK), .RST_AN(n25), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(rf_waddr_m), .DOUT(rf_waddr_wb) );
  DATAPATH_DW01_add_2 add_242 ( .A(IMEM_ADDR[30:0]), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_pls_4_f) );
  BUF_X4 U5 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n13) );
  BUF_X4 U51 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n14) );
  BUF_X4 U52 ( .A(n16), .Z(n18) );
  BUF_X4 U53 ( .A(n16), .Z(n19) );
  BUF_X4 U54 ( .A(n17), .Z(n20) );
  BUF_X4 U55 ( .A(RST_AN), .Z(n26) );
  CLKBUF_X3 U56 ( .A(n28), .Z(n1) );
  CLKBUF_X3 U57 ( .A(n28), .Z(n2) );
  CLKBUF_X3 U59 ( .A(n28), .Z(n6) );
  CLKBUF_X3 U60 ( .A(n151), .Z(n7) );
  CLKBUF_X3 U61 ( .A(n151), .Z(n8) );
  CLKBUF_X3 U62 ( .A(n151), .Z(n9) );
  CLKBUF_X3 U63 ( .A(n150), .Z(n10) );
  CLKBUF_X3 U64 ( .A(n150), .Z(n11) );
  CLKBUF_X3 U65 ( .A(n150), .Z(n12) );
  CLKBUF_X3 U66 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n15) );
  CLKBUF_X2 U67 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n16) );
  CLKBUF_X2 U68 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n17) );
  CLKBUF_X3 U69 ( .A(n17), .Z(n21) );
  CLKBUF_X3 U70 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n22) );
  CLKBUF_X3 U71 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n23) );
  CLKBUF_X3 U72 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n24) );
  CLKBUF_X3 U73 ( .A(RST_AN), .Z(n25) );
  MUX2_X1 U74 ( .A(rf_dout2_e[0]), .B(imm_e[0]), .S(n22), .Z(n108) );
  MUX2_X1 U75 ( .A(rf_dout2_e[1]), .B(imm_e[1]), .S(n22), .Z(n107) );
  MUX2_X1 U76 ( .A(rf_dout2_e[2]), .B(imm_e[2]), .S(n22), .Z(n106) );
  MUX2_X1 U77 ( .A(rf_dout2_e[3]), .B(imm_e[3]), .S(n22), .Z(n105) );
  MUX2_X1 U78 ( .A(rf_dout2_e[4]), .B(imm_e[4]), .S(n22), .Z(n104) );
  MUX2_X1 U79 ( .A(rf_dout2_e[5]), .B(imm_e[5]), .S(n22), .Z(n103) );
  MUX2_X1 U80 ( .A(rf_dout2_e[6]), .B(imm_e[6]), .S(n22), .Z(n102) );
  MUX2_X1 U81 ( .A(rf_dout2_e[7]), .B(imm_e[7]), .S(n22), .Z(n101) );
  MUX2_X1 U82 ( .A(rf_dout2_e[8]), .B(imm_e[8]), .S(n22), .Z(n100) );
  MUX2_X1 U83 ( .A(rf_dout2_e[9]), .B(imm_e[9]), .S(n22), .Z(n99) );
  MUX2_X1 U84 ( .A(rf_dout2_e[10]), .B(imm_e[10]), .S(n22), .Z(n98) );
  MUX2_X1 U85 ( .A(rf_dout2_e[11]), .B(imm_e[11]), .S(n23), .Z(n97) );
  MUX2_X1 U118 ( .A(rf_dout2_e[12]), .B(imm_e[12]), .S(n23), .Z(n96) );
  MUX2_X1 U119 ( .A(rf_dout2_e[13]), .B(imm_e[13]), .S(n23), .Z(n95) );
  MUX2_X1 U120 ( .A(rf_dout2_e[14]), .B(imm_e[14]), .S(n23), .Z(n94) );
  MUX2_X1 U121 ( .A(rf_dout2_e[15]), .B(imm_e[15]), .S(n23), .Z(n93) );
  MUX2_X1 U122 ( .A(rf_dout2_e[16]), .B(imm_e[16]), .S(n23), .Z(n92) );
  MUX2_X1 U123 ( .A(rf_dout2_e[17]), .B(imm_e[17]), .S(n23), .Z(n91) );
  MUX2_X1 U124 ( .A(rf_dout2_e[18]), .B(imm_e[18]), .S(n23), .Z(n90) );
  MUX2_X1 U125 ( .A(rf_dout2_e[19]), .B(imm_e[19]), .S(n23), .Z(n89) );
  MUX2_X1 U126 ( .A(rf_dout2_e[20]), .B(imm_e[20]), .S(n23), .Z(n88) );
  MUX2_X1 U127 ( .A(rf_dout2_e[21]), .B(imm_e[21]), .S(n23), .Z(n87) );
  MUX2_X1 U128 ( .A(rf_dout2_e[22]), .B(imm_e[22]), .S(n24), .Z(n86) );
  MUX2_X1 U129 ( .A(rf_dout2_e[23]), .B(imm_e[23]), .S(n24), .Z(n85) );
  MUX2_X1 U130 ( .A(rf_dout2_e[24]), .B(imm_e[24]), .S(n24), .Z(n84) );
  MUX2_X1 U131 ( .A(rf_dout2_e[25]), .B(imm_e[25]), .S(n24), .Z(n83) );
  MUX2_X1 U132 ( .A(rf_dout2_e[26]), .B(imm_e[26]), .S(n24), .Z(n82) );
  MUX2_X1 U133 ( .A(rf_dout2_e[27]), .B(imm_e[27]), .S(n24), .Z(n81) );
  MUX2_X1 U134 ( .A(rf_dout2_e[28]), .B(imm_e[28]), .S(n24), .Z(n80) );
  MUX2_X1 U135 ( .A(rf_dout2_e[29]), .B(imm_e[29]), .S(n24), .Z(n79) );
  MUX2_X1 U136 ( .A(rf_dout2_e[30]), .B(imm_e[30]), .S(n24), .Z(n78) );
  MUX2_X1 U137 ( .A(rf_dout2_e[31]), .B(imm_e[31]), .S(n24), .Z(n77) );
  MUX2_X1 U138 ( .A(rf_dout1_e[0]), .B(pc_pls_4_e[0]), .S(n21), .Z(alu_a_e[0])
         );
  MUX2_X1 U139 ( .A(rf_dout1_e[1]), .B(pc_pls_4_e[1]), .S(n21), .Z(alu_a_e[1])
         );
  MUX2_X1 U140 ( .A(rf_dout1_e[2]), .B(pc_pls_4_e[2]), .S(n21), .Z(alu_a_e[2])
         );
  MUX2_X1 U141 ( .A(rf_dout1_e[3]), .B(pc_pls_4_e[3]), .S(n21), .Z(alu_a_e[3])
         );
  MUX2_X1 U142 ( .A(rf_dout1_e[4]), .B(pc_pls_4_e[4]), .S(n20), .Z(alu_a_e[4])
         );
  MUX2_X1 U143 ( .A(rf_dout1_e[5]), .B(pc_pls_4_e[5]), .S(n20), .Z(alu_a_e[5])
         );
  MUX2_X1 U144 ( .A(rf_dout1_e[6]), .B(pc_pls_4_e[6]), .S(n20), .Z(alu_a_e[6])
         );
  MUX2_X1 U145 ( .A(rf_dout1_e[7]), .B(pc_pls_4_e[7]), .S(n20), .Z(alu_a_e[7])
         );
  MUX2_X1 U146 ( .A(rf_dout1_e[8]), .B(pc_pls_4_e[8]), .S(n20), .Z(alu_a_e[8])
         );
  MUX2_X1 U147 ( .A(rf_dout1_e[9]), .B(pc_pls_4_e[9]), .S(n20), .Z(alu_a_e[9])
         );
  MUX2_X1 U148 ( .A(rf_dout1_e[10]), .B(pc_pls_4_e[10]), .S(n20), .Z(
        alu_a_e[10]) );
  MUX2_X1 U149 ( .A(rf_dout1_e[11]), .B(pc_pls_4_e[11]), .S(n20), .Z(
        alu_a_e[11]) );
  MUX2_X1 U150 ( .A(rf_dout1_e[12]), .B(pc_pls_4_e[12]), .S(n20), .Z(
        alu_a_e[12]) );
  MUX2_X1 U151 ( .A(rf_dout1_e[13]), .B(pc_pls_4_e[13]), .S(n20), .Z(
        alu_a_e[13]) );
  MUX2_X1 U152 ( .A(rf_dout1_e[14]), .B(pc_pls_4_e[14]), .S(n20), .Z(
        alu_a_e[14]) );
  MUX2_X1 U153 ( .A(rf_dout1_e[15]), .B(pc_pls_4_e[15]), .S(n20), .Z(
        alu_a_e[15]) );
  MUX2_X1 U154 ( .A(rf_dout1_e[16]), .B(pc_pls_4_e[16]), .S(n20), .Z(
        alu_a_e[16]) );
  MUX2_X1 U155 ( .A(rf_dout1_e[17]), .B(pc_pls_4_e[17]), .S(n20), .Z(
        alu_a_e[17]) );
  MUX2_X1 U156 ( .A(rf_dout1_e[18]), .B(pc_pls_4_e[18]), .S(n20), .Z(
        alu_a_e[18]) );
  XOR2_X1 U157 ( .A(\DP_SIG[CMPR_0_IS_0_M] ), .B(\CTRL_WORD[COMP_0_INVERT] ), 
        .Z(n27) );
  MUX2_X1 U158 ( .A(\CTRL_WORD[JUMP_EN] ), .B(n27), .S(\CTRL_WORD[BRANCH_EN] ), 
        .Z(n184) );
  INV_X1 U159 ( .A(n184), .ZN(n28) );
  MUX2_X1 U160 ( .A(DMEM_RWADDR[0]), .B(pc_pls_4_f[0]), .S(n1), .Z(n109) );
  MUX2_X1 U161 ( .A(DMEM_RWADDR[1]), .B(pc_pls_4_f[1]), .S(n1), .Z(n58) );
  MUX2_X1 U162 ( .A(DMEM_RWADDR[2]), .B(pc_pls_4_f[2]), .S(n1), .Z(n57) );
  MUX2_X1 U163 ( .A(DMEM_RWADDR[3]), .B(pc_pls_4_f[3]), .S(n1), .Z(n56) );
  MUX2_X1 U168 ( .A(DMEM_RWADDR[4]), .B(pc_pls_4_f[4]), .S(n1), .Z(n55) );
  MUX2_X1 U169 ( .A(DMEM_RWADDR[5]), .B(pc_pls_4_f[5]), .S(n1), .Z(n54) );
  MUX2_X1 U190 ( .A(DMEM_RWADDR[6]), .B(pc_pls_4_f[6]), .S(n1), .Z(n53) );
  MUX2_X1 U191 ( .A(DMEM_RWADDR[7]), .B(pc_pls_4_f[7]), .S(n1), .Z(n52) );
  MUX2_X1 U194 ( .A(DMEM_RWADDR[8]), .B(pc_pls_4_f[8]), .S(n1), .Z(n51) );
  MUX2_X1 U195 ( .A(DMEM_RWADDR[9]), .B(pc_pls_4_f[9]), .S(n1), .Z(n50) );
  MUX2_X1 U196 ( .A(DMEM_RWADDR[10]), .B(pc_pls_4_f[10]), .S(n1), .Z(n49) );
  MUX2_X1 U197 ( .A(DMEM_RWADDR[11]), .B(pc_pls_4_f[11]), .S(n2), .Z(n48) );
  MUX2_X1 U198 ( .A(DMEM_RWADDR[12]), .B(pc_pls_4_f[12]), .S(n2), .Z(n47) );
  MUX2_X1 U199 ( .A(DMEM_RWADDR[13]), .B(pc_pls_4_f[13]), .S(n2), .Z(n46) );
  MUX2_X1 U200 ( .A(DMEM_RWADDR[14]), .B(pc_pls_4_f[14]), .S(n2), .Z(n45) );
  MUX2_X1 U201 ( .A(DMEM_RWADDR[15]), .B(pc_pls_4_f[15]), .S(n2), .Z(n44) );
  MUX2_X1 U202 ( .A(DMEM_RWADDR[16]), .B(pc_pls_4_f[16]), .S(n2), .Z(n43) );
  MUX2_X1 U203 ( .A(DMEM_RWADDR[17]), .B(pc_pls_4_f[17]), .S(n2), .Z(n42) );
  MUX2_X1 U204 ( .A(DMEM_RWADDR[18]), .B(pc_pls_4_f[18]), .S(n2), .Z(n41) );
  MUX2_X1 U205 ( .A(DMEM_RWADDR[19]), .B(pc_pls_4_f[19]), .S(n2), .Z(n40) );
  MUX2_X1 U206 ( .A(DMEM_RWADDR[20]), .B(pc_pls_4_f[20]), .S(n2), .Z(n39) );
  MUX2_X1 U207 ( .A(DMEM_RWADDR[21]), .B(pc_pls_4_f[21]), .S(n2), .Z(n38) );
  MUX2_X1 U208 ( .A(DMEM_RWADDR[22]), .B(pc_pls_4_f[22]), .S(n6), .Z(n37) );
  MUX2_X1 U209 ( .A(DMEM_RWADDR[23]), .B(pc_pls_4_f[23]), .S(n6), .Z(n36) );
  MUX2_X1 U210 ( .A(DMEM_RWADDR[24]), .B(pc_pls_4_f[24]), .S(n6), .Z(n35) );
  MUX2_X1 U211 ( .A(DMEM_RWADDR[25]), .B(pc_pls_4_f[25]), .S(n6), .Z(n34) );
  MUX2_X1 U212 ( .A(DMEM_RWADDR[26]), .B(pc_pls_4_f[26]), .S(n6), .Z(n33) );
  MUX2_X1 U213 ( .A(DMEM_RWADDR[27]), .B(pc_pls_4_f[27]), .S(n6), .Z(n32) );
  MUX2_X1 U214 ( .A(DMEM_RWADDR[28]), .B(pc_pls_4_f[28]), .S(n6), .Z(n31) );
  MUX2_X1 U215 ( .A(DMEM_RWADDR[29]), .B(pc_pls_4_f[29]), .S(n6), .Z(n30) );
  MUX2_X1 U216 ( .A(DMEM_RWADDR[30]), .B(pc_pls_4_f[30]), .S(n6), .Z(n29) );
  INV_X2 U217 ( .A(n144), .ZN(n59) );
  INV_X2 U218 ( .A(n145), .ZN(n60) );
  INV_X2 U219 ( .A(n146), .ZN(n61) );
  INV_X2 U220 ( .A(n147), .ZN(n62) );
  INV_X2 U221 ( .A(n148), .ZN(n63) );
  INV_X2 U222 ( .A(rf_dout1_e[31]), .ZN(n64) );
  INV_X2 U223 ( .A(rf_dout1_e[30]), .ZN(n65) );
  INV_X2 U224 ( .A(rf_dout1_e[29]), .ZN(n66) );
  INV_X2 U225 ( .A(rf_dout1_e[28]), .ZN(n67) );
  INV_X2 U226 ( .A(rf_dout1_e[27]), .ZN(n68) );
  INV_X2 U227 ( .A(rf_dout1_e[26]), .ZN(n69) );
  INV_X2 U228 ( .A(rf_dout1_e[25]), .ZN(n70) );
  INV_X2 U229 ( .A(rf_dout1_e[24]), .ZN(n71) );
  INV_X2 U230 ( .A(rf_dout1_e[23]), .ZN(n72) );
  INV_X2 U231 ( .A(rf_dout1_e[22]), .ZN(n73) );
  INV_X2 U232 ( .A(rf_dout1_e[21]), .ZN(n74) );
  INV_X2 U233 ( .A(rf_dout1_e[20]), .ZN(n75) );
  INV_X2 U234 ( .A(rf_dout1_e[19]), .ZN(n76) );
  INV_X2 U235 ( .A(n158), .ZN(n110) );
  INV_X2 U236 ( .A(n159), .ZN(n111) );
  INV_X2 U237 ( .A(n161), .ZN(n112) );
  INV_X2 U238 ( .A(n162), .ZN(n113) );
  INV_X2 U239 ( .A(n163), .ZN(n114) );
  INV_X2 U240 ( .A(n164), .ZN(n115) );
  INV_X2 U241 ( .A(n165), .ZN(n116) );
  INV_X2 U242 ( .A(n166), .ZN(n117) );
  INV_X2 U243 ( .A(n167), .ZN(n118) );
  INV_X2 U244 ( .A(n168), .ZN(n119) );
  INV_X2 U245 ( .A(n169), .ZN(n120) );
  INV_X2 U246 ( .A(n170), .ZN(n121) );
  INV_X2 U247 ( .A(n172), .ZN(n122) );
  INV_X2 U248 ( .A(n173), .ZN(n123) );
  INV_X2 U249 ( .A(n174), .ZN(n124) );
  INV_X2 U250 ( .A(n175), .ZN(n125) );
  INV_X2 U251 ( .A(n176), .ZN(n126) );
  INV_X2 U252 ( .A(n177), .ZN(n127) );
  INV_X2 U253 ( .A(n178), .ZN(n128) );
  INV_X2 U254 ( .A(n179), .ZN(n129) );
  INV_X2 U255 ( .A(n180), .ZN(n130) );
  INV_X2 U256 ( .A(n181), .ZN(n131) );
  INV_X2 U257 ( .A(n149), .ZN(n132) );
  INV_X2 U258 ( .A(n152), .ZN(n133) );
  INV_X2 U259 ( .A(n153), .ZN(n134) );
  INV_X2 U260 ( .A(n154), .ZN(n135) );
  INV_X2 U261 ( .A(n155), .ZN(n136) );
  INV_X2 U262 ( .A(n156), .ZN(n137) );
  INV_X2 U263 ( .A(n157), .ZN(n138) );
  INV_X2 U264 ( .A(n160), .ZN(n139) );
  INV_X2 U265 ( .A(n171), .ZN(n140) );
  INV_X2 U266 ( .A(n182), .ZN(n141) );
  INV_X2 U267 ( .A(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n142) );
  INV_X2 U268 ( .A(\CTRL_WORD[R_TYPE_SEL] ), .ZN(n143) );
  INV_X2 U269 ( .A(\CTRL_WORD[JAL_EN] ), .ZN(n183) );
endmodule


module HU ( CLK, RST_AN, .DP_SIG({\DP_SIG[CMPR_0_IS_0_M] , 
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }), 
    .HZRD_SIG({\HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , 
        \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , 
        \HZRD_SIG[FLUSH_MWB] }) );
  input CLK, RST_AN, \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  output \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] ,
         \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] ;
  wire   \HZRD_SIG[FLUSH_FD] , n2, n3, n4, n1;
  assign \HZRD_SIG[FLUSH_MWB]  = 1'b0;
  assign \HZRD_SIG[STALL_DE]  = 1'b0;
  assign \HZRD_SIG[STALL_FD]  = 1'b0;
  assign \HZRD_SIG[FLUSH_EM]  = \HZRD_SIG[FLUSH_FD] ;
  assign \HZRD_SIG[FLUSH_DE]  = \HZRD_SIG[FLUSH_FD] ;

  NOR4_X2 U3 ( .A1(\DP_SIG[INSTR_OPCODE_M][3] ), .A2(n2), .A3(
        \DP_SIG[INSTR_OPCODE_M][5] ), .A4(\DP_SIG[INSTR_OPCODE_M][4] ), .ZN(
        \HZRD_SIG[FLUSH_FD] ) );
  AOI22_X2 U4 ( .A1(n3), .A2(\DP_SIG[INSTR_OPCODE_M][2] ), .B1(
        \DP_SIG[INSTR_OPCODE_M][1] ), .B2(n1), .ZN(n2) );
  NOR2_X2 U5 ( .A1(\DP_SIG[INSTR_OPCODE_M][1] ), .A2(n4), .ZN(n3) );
  XNOR2_X2 U6 ( .A(\DP_SIG[INSTR_OPCODE_M][0] ), .B(\DP_SIG[CMPR_0_IS_0_M] ), 
        .ZN(n4) );
  INV_X2 U7 ( .A(\DP_SIG[INSTR_OPCODE_M][2] ), .ZN(n1) );
endmodule


module CPU ( CLK, RST_AN, IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, DMEM_WEN, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN;
  output DMEM_WEN;
  wire   \hzrd_sig[FLUSH_FD] , \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] ,
         \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] ,
         \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] ,
         \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] ,
         \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] ,
         \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] ,
         \ctrl_word[COMP_0_INVERT] , \ctrl_word[RF_WB_DMEM_DOUT_SEL] ,
         \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] , \dp_sig[CMPR_0_IS_0_M] ,
         \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] ,
         \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] ,
         \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] ;
  wire   [31:0] instr_cu;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  CU U_CU ( .CLK(CLK), .RST_AN(RST_AN), .INSTR(instr_cu), .HZRD_SIG({1'b0, 
        \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        1'b0}), .CTRL_WORD({\ctrl_word[J_TYPE_IMM_SEL] , 
        \ctrl_word[R_TYPE_SEL] , \ctrl_word[IMM_SEL] , 
        \ctrl_word[PC_PLS_4_SEL] , \ctrl_word[ALU_FUNC][3] , 
        \ctrl_word[ALU_FUNC][2] , \ctrl_word[ALU_FUNC][1] , 
        \ctrl_word[ALU_FUNC][0] , \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }) );
  DATAPATH U_DATAPATH ( .CLK(CLK), .RST_AN(RST_AN), .CTRL_WORD({
        \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] , 
        \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] , 
        \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] , 
        \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] , 
        \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }), .INSTR_CU(instr_cu), 
        .HZRD_SIG({1'b0, \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , 
        \hzrd_sig[FLUSH_EM] , 1'b0}), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), 
        .IMEM_ADDR(IMEM_ADDR), .IMEM_DOUT(IMEM_DOUT), .DMEM_RWADDR(DMEM_RWADDR), .DMEM_DIN(DMEM_DIN), .DMEM_DOUT(DMEM_DOUT) );
  HU U_HU ( .CLK(CLK), .RST_AN(RST_AN), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), .HZRD_SIG(
        {SYNOPSYS_UNCONNECTED__0, \hzrd_sig[FLUSH_FD] , 
        SYNOPSYS_UNCONNECTED__1, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        SYNOPSYS_UNCONNECTED__2}) );
endmodule

