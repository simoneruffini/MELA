
module CU ( CLK, RST_AN, INSTR, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .CTRL_WORD({
        \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] , 
        \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] , 
        \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] , 
        \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] , 
        \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }) );
  input [31:0] INSTR;
  input CLK, RST_AN, \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] ;
  wire   INSTR_31, INSTR_30, INSTR_29, INSTR_28, INSTR_27, INSTR_26,
         \execute_sig_d1[R_TYPE_SEL] , \execute_sig_d1[IMM_SEL] ,
         \execute_sig_d1[PC_PLS_4_SEL] , \execute_sig_d1[ALU_FUNC][3] ,
         \execute_sig_d1[ALU_FUNC][2] , \execute_sig_d1[ALU_FUNC][1] ,
         \execute_sig_d1[ALU_FUNC][0] , \memory_sig_d1[DMEM_WEN] ,
         \memory_sig_d1[BRANCH_EN] , \memory_sig_d1[JUMP_EN] ,
         \memory_sig_d1[COMP_0_INVERT] ,
         \writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d1[JAL_EN] ,
         \writeback_sig_d1[RF_WEN] , \memory_sig_d2[DMEM_WEN] ,
         \memory_sig_d2[BRANCH_EN] , \memory_sig_d2[JUMP_EN] ,
         \memory_sig_d2[COMP_0_INVERT] ,
         \writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] , \writeback_sig_d2[JAL_EN] ,
         \writeback_sig_d2[RF_WEN] , \writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ,
         \writeback_sig_d3[JAL_EN] , \writeback_sig_d3[RF_WEN] , N213, N214,
         N215, N216, N217, N218, N224, N228, N229, N231, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n117,
         n118, n119, n120, n121, n122, n123, n124;
  assign INSTR_31 = INSTR[31];
  assign INSTR_30 = INSTR[30];
  assign INSTR_29 = INSTR[29];
  assign INSTR_28 = INSTR[28];
  assign INSTR_27 = INSTR[27];
  assign INSTR_26 = INSTR[26];

  DFFR_X1 \decode_sig_d1_reg[J_TYPE_IMM_SEL]  ( .D(n38), .CK(CLK), .RN(n30), 
        .Q(\CTRL_WORD[J_TYPE_IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[IMM_SEL]  ( .D(N218), .CK(CLK), .RN(n30), .Q(
        \execute_sig_d1[IMM_SEL] ) );
  DFFR_X1 \execute_sig_d1_reg[PC_PLS_4_SEL]  ( .D(N217), .CK(CLK), .RN(n30), 
        .Q(\execute_sig_d1[PC_PLS_4_SEL] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][3]  ( .D(N216), .CK(CLK), .SN(n33), 
        .Q(\execute_sig_d1[ALU_FUNC][3] ) );
  DFFR_X1 \execute_sig_d1_reg[ALU_FUNC][2]  ( .D(N215), .CK(CLK), .RN(n30), 
        .Q(\execute_sig_d1[ALU_FUNC][2] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][1]  ( .D(N214), .CK(CLK), .SN(n33), 
        .Q(\execute_sig_d1[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d1_reg[ALU_FUNC][0]  ( .D(N213), .CK(CLK), .SN(n33), 
        .Q(\execute_sig_d1[ALU_FUNC][0] ) );
  DFFR_X1 \memory_sig_d1_reg[BRANCH_EN]  ( .D(n39), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d1[BRANCH_EN] ) );
  DFFR_X1 \memory_sig_d1_reg[JUMP_EN]  ( .D(n38), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d1[JUMP_EN] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n36), .CK(CLK), 
        .RN(n30), .Q(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d1_reg[RF_WEN]  ( .D(N224), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d1[RF_WEN] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][3]  ( .D(N231), .CK(CLK), .SN(n32), 
        .Q(\CTRL_WORD[ALU_FUNC][3] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][1]  ( .D(N229), .CK(CLK), .SN(n33), 
        .Q(\CTRL_WORD[ALU_FUNC][1] ) );
  DFFS_X1 \execute_sig_d2_reg[ALU_FUNC][0]  ( .D(N228), .CK(CLK), .SN(n32), 
        .Q(\CTRL_WORD[ALU_FUNC][0] ) );
  NAND3_X1 U118 ( .A1(n68), .A2(n41), .A3(INSTR_31), .ZN(n54) );
  NAND3_X1 U119 ( .A1(INSTR_29), .A2(n117), .A3(n47), .ZN(n71) );
  NAND3_X1 U120 ( .A1(INSTR_26), .A2(n80), .A3(INSTR_29), .ZN(n79) );
  OAI33_X1 U121 ( .A1(n123), .A2(INSTR[5]), .A3(n120), .B1(n124), .B2(INSTR[2]), .B3(n98), .ZN(n97) );
  NAND3_X1 U122 ( .A1(INSTR_26), .A2(n52), .A3(INSTR_27), .ZN(n77) );
  NAND3_X1 U123 ( .A1(INSTR_27), .A2(n46), .A3(INSTR_28), .ZN(n108) );
  NAND3_X1 U124 ( .A1(n96), .A2(n118), .A3(INSTR_30), .ZN(n110) );
  NAND3_X1 U125 ( .A1(n113), .A2(n122), .A3(INSTR[2]), .ZN(n104) );
  NAND3_X1 U126 ( .A1(n113), .A2(n121), .A3(INSTR[3]), .ZN(n98) );
  NAND3_X1 U127 ( .A1(n113), .A2(INSTR[5]), .A3(INSTR[1]), .ZN(n114) );
  NAND3_X1 U128 ( .A1(n40), .A2(INSTR_27), .A3(n116), .ZN(n55) );
  DFFRS_X2 \execute_sig_d2_reg[IMM_SEL]  ( .D(n27), .CK(CLK), .RN(n31), .SN(
        1'b1), .Q(\CTRL_WORD[IMM_SEL] ) );
  SDFFR_X1 \execute_sig_d2_reg[PC_PLS_4_SEL]  ( .D(1'b0), .SI(n35), .SE(
        \execute_sig_d1[PC_PLS_4_SEL] ), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[PC_PLS_4_SEL] ) );
  SDFFR_X1 \writeback_sig_d4_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(1'b0), .SI(n42), 
        .SE(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ), .CK(CLK), .RN(n32), .Q(
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d3_reg[RF_WEN]  ( .D(n23), .CK(CLK), .RN(RST_AN), .Q(
        \writeback_sig_d3[RF_WEN] ) );
  DFFR_X1 \writeback_sig_d3_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n22), .CK(CLK), 
        .RN(n32), .Q(\writeback_sig_d3[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d3_reg[JAL_EN]  ( .D(n21), .CK(CLK), .RN(n32), .Q(
        \writeback_sig_d3[JAL_EN] ) );
  DFFR_X1 \memory_sig_d3_reg[JUMP_EN]  ( .D(n20), .CK(CLK), .RN(n32), .Q(
        \CTRL_WORD[JUMP_EN] ) );
  DFFR_X1 \memory_sig_d3_reg[DMEM_WEN]  ( .D(n19), .CK(CLK), .RN(n32), .Q(
        \CTRL_WORD[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d3_reg[COMP_0_INVERT]  ( .D(n18), .CK(CLK), .RN(n32), 
        .Q(\CTRL_WORD[COMP_0_INVERT] ) );
  DFFR_X1 \memory_sig_d3_reg[BRANCH_EN]  ( .D(n17), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[BRANCH_EN] ) );
  DFFR_X1 \execute_sig_d1_reg[R_TYPE_SEL]  ( .D(n16), .CK(CLK), .RN(n31), .Q(
        \execute_sig_d1[R_TYPE_SEL] ) );
  DFFR_X1 \writeback_sig_d2_reg[RF_WEN]  ( .D(n15), .CK(CLK), .RN(n32), .Q(
        \writeback_sig_d2[RF_WEN] ) );
  DFFR_X1 \writeback_sig_d2_reg[RF_WB_DMEM_DOUT_SEL]  ( .D(n14), .CK(CLK), 
        .RN(n31), .Q(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ) );
  DFFR_X1 \writeback_sig_d2_reg[JAL_EN]  ( .D(n13), .CK(CLK), .RN(n32), .Q(
        \writeback_sig_d2[JAL_EN] ) );
  DFFR_X1 \memory_sig_d2_reg[JUMP_EN]  ( .D(n12), .CK(CLK), .RN(n31), .Q(
        \memory_sig_d2[JUMP_EN] ) );
  DFFR_X1 \memory_sig_d2_reg[DMEM_WEN]  ( .D(n11), .CK(CLK), .RN(n31), .Q(
        \memory_sig_d2[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d2_reg[COMP_0_INVERT]  ( .D(n10), .CK(CLK), .RN(n31), 
        .Q(\memory_sig_d2[COMP_0_INVERT] ) );
  DFFR_X1 \memory_sig_d2_reg[BRANCH_EN]  ( .D(n9), .CK(CLK), .RN(n31), .Q(
        \memory_sig_d2[BRANCH_EN] ) );
  DFFR_X1 \execute_sig_d2_reg[R_TYPE_SEL]  ( .D(n8), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[R_TYPE_SEL] ) );
  DFFR_X1 \execute_sig_d2_reg[ALU_FUNC][2]  ( .D(n7), .CK(CLK), .RN(n31), .Q(
        \CTRL_WORD[ALU_FUNC][2] ) );
  DFFR_X1 \memory_sig_d1_reg[DMEM_WEN]  ( .D(n6), .CK(CLK), .RN(n31), .Q(
        \memory_sig_d1[DMEM_WEN] ) );
  DFFR_X1 \memory_sig_d1_reg[COMP_0_INVERT]  ( .D(n5), .CK(CLK), .RN(n30), .Q(
        \memory_sig_d1[COMP_0_INVERT] ) );
  DFFR_X1 \writeback_sig_d1_reg[JAL_EN]  ( .D(n4), .CK(CLK), .RN(n30), .Q(
        \writeback_sig_d1[JAL_EN] ) );
  DFFR_X1 \writeback_sig_d4_reg[RF_WEN]  ( .D(n3), .CK(CLK), .RN(n30), .Q(
        \CTRL_WORD[RF_WEN] ) );
  DFFRS_X2 \writeback_sig_d4_reg[JAL_EN]  ( .D(n2), .CK(CLK), .RN(RST_AN), 
        .SN(1'b1), .Q(\CTRL_WORD[JAL_EN] ) );
  AND2_X1 U4 ( .A1(\writeback_sig_d3[JAL_EN] ), .A2(n42), .ZN(n2) );
  AND2_X1 U5 ( .A1(\writeback_sig_d3[RF_WEN] ), .A2(n42), .ZN(n3) );
  AND2_X1 U6 ( .A1(INSTR_26), .A2(n38), .ZN(n4) );
  AND2_X1 U7 ( .A1(INSTR_26), .A2(n39), .ZN(n5) );
  AND2_X1 U8 ( .A1(INSTR_29), .A2(n36), .ZN(n6) );
  AND2_X1 U9 ( .A1(\execute_sig_d1[ALU_FUNC][2] ), .A2(n35), .ZN(n7) );
  AND2_X1 U10 ( .A1(\execute_sig_d1[R_TYPE_SEL] ), .A2(n35), .ZN(n8) );
  AND2_X1 U11 ( .A1(\memory_sig_d1[BRANCH_EN] ), .A2(n35), .ZN(n9) );
  AND2_X1 U12 ( .A1(\memory_sig_d1[COMP_0_INVERT] ), .A2(n35), .ZN(n10) );
  AND2_X1 U13 ( .A1(\memory_sig_d1[DMEM_WEN] ), .A2(n35), .ZN(n11) );
  AND2_X1 U14 ( .A1(\memory_sig_d1[JUMP_EN] ), .A2(n35), .ZN(n12) );
  AND2_X1 U15 ( .A1(\writeback_sig_d1[JAL_EN] ), .A2(n35), .ZN(n13) );
  AND2_X1 U16 ( .A1(\writeback_sig_d1[RF_WB_DMEM_DOUT_SEL] ), .A2(n35), .ZN(
        n14) );
  AND2_X1 U17 ( .A1(\writeback_sig_d1[RF_WEN] ), .A2(n35), .ZN(n15) );
  AND2_X1 U18 ( .A1(n44), .A2(n41), .ZN(n16) );
  AND2_X1 U19 ( .A1(\memory_sig_d2[BRANCH_EN] ), .A2(n34), .ZN(n17) );
  AND2_X1 U20 ( .A1(\memory_sig_d2[COMP_0_INVERT] ), .A2(n34), .ZN(n18) );
  AND2_X1 U21 ( .A1(\memory_sig_d2[DMEM_WEN] ), .A2(n34), .ZN(n19) );
  AND2_X1 U22 ( .A1(\memory_sig_d2[JUMP_EN] ), .A2(n34), .ZN(n20) );
  AND2_X1 U23 ( .A1(\writeback_sig_d2[JAL_EN] ), .A2(n34), .ZN(n21) );
  AND2_X1 U24 ( .A1(\writeback_sig_d2[RF_WB_DMEM_DOUT_SEL] ), .A2(n34), .ZN(
        n22) );
  AND2_X1 U25 ( .A1(\writeback_sig_d2[RF_WEN] ), .A2(n34), .ZN(n23) );
  INV_X1 U28 ( .A(n67), .ZN(n40) );
  INV_X1 U29 ( .A(n64), .ZN(n39) );
  INV_X1 U30 ( .A(\HZRD_SIG[FLUSH_FD] ), .ZN(n41) );
  INV_X1 U31 ( .A(\HZRD_SIG[FLUSH_DE] ), .ZN(n35) );
  INV_X1 U32 ( .A(\HZRD_SIG[FLUSH_EM] ), .ZN(n34) );
  AOI21_X1 U33 ( .B1(n56), .B2(n57), .A(\HZRD_SIG[FLUSH_FD] ), .ZN(N224) );
  OAI21_X1 U34 ( .B1(n60), .B2(n61), .A(n43), .ZN(n56) );
  OAI211_X1 U35 ( .C1(n58), .C2(n59), .A(n52), .B(n46), .ZN(n57) );
  OAI22_X1 U36 ( .A1(n52), .A2(n49), .B1(n51), .B2(n62), .ZN(n61) );
  NAND2_X1 U37 ( .A1(n41), .A2(n43), .ZN(n67) );
  NAND4_X1 U38 ( .A1(n50), .A2(n40), .A3(n117), .A4(n46), .ZN(n64) );
  OAI211_X1 U39 ( .C1(n99), .C2(n74), .A(n100), .B(n37), .ZN(N213) );
  OAI211_X1 U40 ( .C1(n106), .C2(n107), .A(n74), .B(n43), .ZN(n100) );
  NOR3_X1 U41 ( .A1(n112), .A2(n81), .A3(n88), .ZN(n99) );
  OAI211_X1 U42 ( .C1(n109), .C2(n117), .A(n110), .B(n95), .ZN(n106) );
  OAI211_X1 U43 ( .C1(n66), .C2(n67), .A(n55), .B(n54), .ZN(N218) );
  AOI21_X1 U44 ( .B1(n53), .B2(n69), .A(n60), .ZN(n66) );
  INV_X1 U45 ( .A(n55), .ZN(n38) );
  INV_X1 U46 ( .A(n101), .ZN(n37) );
  OAI221_X1 U47 ( .B1(n68), .B2(n43), .C1(n102), .C2(n74), .A(n41), .ZN(n101)
         );
  NOR2_X1 U48 ( .A1(n103), .A2(n89), .ZN(n102) );
  NOR3_X1 U49 ( .A1(n104), .A2(n105), .A3(n124), .ZN(n103) );
  NAND2_X1 U50 ( .A1(n64), .A2(n55), .ZN(N217) );
  INV_X1 U51 ( .A(n54), .ZN(n36) );
  BUF_X1 U52 ( .A(n28), .Z(n31) );
  BUF_X1 U53 ( .A(n29), .Z(n32) );
  BUF_X1 U54 ( .A(n28), .Z(n30) );
  INV_X1 U55 ( .A(n74), .ZN(n44) );
  AOI21_X1 U56 ( .B1(n72), .B2(n85), .A(n117), .ZN(n84) );
  INV_X1 U57 ( .A(n96), .ZN(n50) );
  NAND2_X1 U58 ( .A1(n86), .A2(n118), .ZN(n72) );
  INV_X1 U59 ( .A(n69), .ZN(n47) );
  INV_X1 U60 ( .A(n98), .ZN(n119) );
  INV_X1 U61 ( .A(n62), .ZN(n53) );
  INV_X1 U62 ( .A(n87), .ZN(n120) );
  BUF_X1 U63 ( .A(n29), .Z(n33) );
  INV_X1 U64 ( .A(n105), .ZN(n121) );
  INV_X1 U65 ( .A(n63), .ZN(n49) );
  NOR3_X1 U66 ( .A1(INSTR_28), .A2(INSTR_30), .A3(INSTR_29), .ZN(n116) );
  OAI221_X1 U67 ( .B1(n73), .B2(n74), .C1(n44), .C2(n75), .A(n41), .ZN(N216)
         );
  AOI21_X1 U68 ( .B1(INSTR[0]), .B2(n119), .A(n81), .ZN(n73) );
  AOI221_X1 U69 ( .B1(n76), .B2(n51), .C1(INSTR_31), .C2(n77), .A(n78), .ZN(
        n75) );
  OAI221_X1 U70 ( .B1(INSTR_27), .B2(n69), .C1(n50), .C2(n46), .A(n79), .ZN(
        n78) );
  OAI211_X1 U71 ( .C1(n90), .C2(n74), .A(n91), .B(n37), .ZN(N214) );
  AOI21_X1 U72 ( .B1(n87), .B2(n121), .A(n97), .ZN(n90) );
  OAI211_X1 U73 ( .C1(n92), .C2(n48), .A(n74), .B(n43), .ZN(n91) );
  OAI21_X1 U74 ( .B1(n82), .B2(n65), .A(n83), .ZN(N215) );
  AOI211_X1 U75 ( .C1(INSTR[1]), .C2(n87), .A(n88), .B(n89), .ZN(n82) );
  NAND2_X1 U76 ( .A1(n44), .A2(n41), .ZN(n65) );
  OAI211_X1 U77 ( .C1(n84), .C2(n63), .A(n40), .B(INSTR_28), .ZN(n83) );
  OR2_X1 U78 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][0] ), 
        .ZN(N228) );
  OR2_X1 U79 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][1] ), 
        .ZN(N229) );
  OR2_X1 U80 ( .A1(\HZRD_SIG[FLUSH_DE] ), .A2(\execute_sig_d1[ALU_FUNC][3] ), 
        .ZN(N231) );
  NOR4_X1 U81 ( .A1(n123), .A2(n104), .A3(n124), .A4(INSTR[5]), .ZN(n89) );
  NAND4_X1 U82 ( .A1(n117), .A2(n52), .A3(n118), .A4(n111), .ZN(n74) );
  NOR3_X1 U83 ( .A1(INSTR_29), .A2(INSTR_31), .A3(INSTR_30), .ZN(n111) );
  NOR4_X1 U84 ( .A1(INSTR[6]), .A2(INSTR[4]), .A3(INSTR[10]), .A4(n115), .ZN(
        n113) );
  OR3_X1 U85 ( .A1(INSTR[9]), .A2(INSTR[8]), .A3(INSTR[7]), .ZN(n115) );
  NOR4_X1 U86 ( .A1(n114), .A2(INSTR[0]), .A3(INSTR[3]), .A4(INSTR[2]), .ZN(
        n112) );
  NOR3_X1 U87 ( .A1(INSTR[1]), .A2(INSTR[5]), .A3(n120), .ZN(n88) );
  INV_X1 U88 ( .A(INSTR_27), .ZN(n117) );
  INV_X1 U89 ( .A(INSTR[3]), .ZN(n122) );
  AOI211_X1 U90 ( .C1(INSTR_29), .C2(n43), .A(n117), .B(n118), .ZN(n58) );
  NOR2_X1 U91 ( .A1(n104), .A2(INSTR[0]), .ZN(n87) );
  INV_X1 U92 ( .A(INSTR_28), .ZN(n52) );
  NOR2_X1 U93 ( .A1(n51), .A2(INSTR_30), .ZN(n86) );
  OAI22_X1 U94 ( .A1(INSTR_29), .A2(n45), .B1(INSTR_27), .B2(n85), .ZN(n107)
         );
  INV_X1 U95 ( .A(n76), .ZN(n45) );
  OAI211_X1 U96 ( .C1(n46), .C2(n70), .A(n71), .B(n72), .ZN(n60) );
  INV_X1 U97 ( .A(INSTR_31), .ZN(n43) );
  NOR3_X1 U98 ( .A1(INSTR_26), .A2(INSTR_31), .A3(INSTR_27), .ZN(n59) );
  OAI21_X1 U99 ( .B1(INSTR_28), .B2(INSTR_27), .A(n108), .ZN(n76) );
  NOR2_X1 U100 ( .A1(n85), .A2(INSTR_26), .ZN(n63) );
  INV_X1 U101 ( .A(INSTR_29), .ZN(n51) );
  NOR2_X1 U102 ( .A1(n77), .A2(INSTR_30), .ZN(n68) );
  INV_X1 U103 ( .A(INSTR_30), .ZN(n46) );
  AOI21_X1 U104 ( .B1(INSTR_29), .B2(n52), .A(n47), .ZN(n109) );
  OAI211_X1 U105 ( .C1(INSTR_29), .C2(n94), .A(n70), .B(n95), .ZN(n92) );
  AOI21_X1 U106 ( .B1(n117), .B2(n52), .A(n47), .ZN(n94) );
  NAND2_X1 U107 ( .A1(INSTR_30), .A2(n51), .ZN(n85) );
  INV_X1 U108 ( .A(INSTR_26), .ZN(n118) );
  NAND2_X1 U109 ( .A1(INSTR_28), .A2(n117), .ZN(n62) );
  NAND2_X1 U110 ( .A1(INSTR_30), .A2(INSTR_26), .ZN(n69) );
  OAI22_X1 U111 ( .A1(INSTR_31), .A2(INSTR_28), .B1(n117), .B2(n52), .ZN(n80)
         );
  INV_X1 U112 ( .A(INSTR[0]), .ZN(n124) );
  NAND2_X1 U113 ( .A1(n86), .A2(INSTR_26), .ZN(n95) );
  AND3_X1 U114 ( .A1(n119), .A2(n124), .A3(INSTR[2]), .ZN(n81) );
  NAND2_X1 U115 ( .A1(INSTR[5]), .A2(n123), .ZN(n105) );
  NAND2_X1 U116 ( .A1(n50), .A2(INSTR_27), .ZN(n70) );
  INV_X1 U117 ( .A(INSTR[1]), .ZN(n123) );
  NAND2_X1 U129 ( .A1(INSTR_28), .A2(n51), .ZN(n96) );
  INV_X1 U130 ( .A(n93), .ZN(n48) );
  AOI22_X1 U131 ( .A1(n86), .A2(n53), .B1(n62), .B2(INSTR_30), .ZN(n93) );
  BUF_X1 U132 ( .A(RST_AN), .Z(n29) );
  BUF_X1 U133 ( .A(RST_AN), .Z(n28) );
  INV_X1 U134 ( .A(\HZRD_SIG[FLUSH_MWB] ), .ZN(n42) );
  AND2_X1 U136 ( .A1(\execute_sig_d1[IMM_SEL] ), .A2(n35), .ZN(n27) );
endmodule


module REG_PIPO_32_fffffffc_fffffffc ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n17, n18, n19;

  DFFS_X1 \reg_mem_reg[31]  ( .D(n96), .CK(CLK), .SN(n19), .Q(DOUT[31]), .QN(
        n64) );
  DFFS_X1 \reg_mem_reg[30]  ( .D(n95), .CK(CLK), .SN(n19), .Q(DOUT[30]) );
  DFFS_X1 \reg_mem_reg[29]  ( .D(n94), .CK(CLK), .SN(n19), .Q(DOUT[29]) );
  DFFS_X1 \reg_mem_reg[28]  ( .D(n93), .CK(CLK), .SN(n19), .Q(DOUT[28]) );
  DFFS_X1 \reg_mem_reg[27]  ( .D(n92), .CK(CLK), .SN(n19), .Q(DOUT[27]) );
  DFFS_X1 \reg_mem_reg[26]  ( .D(n91), .CK(CLK), .SN(n19), .Q(DOUT[26]) );
  DFFS_X1 \reg_mem_reg[25]  ( .D(n90), .CK(CLK), .SN(n18), .Q(DOUT[25]) );
  DFFS_X1 \reg_mem_reg[24]  ( .D(n89), .CK(CLK), .SN(n18), .Q(DOUT[24]) );
  DFFS_X1 \reg_mem_reg[23]  ( .D(n88), .CK(CLK), .SN(n18), .Q(DOUT[23]) );
  DFFS_X1 \reg_mem_reg[22]  ( .D(n87), .CK(CLK), .SN(n18), .Q(DOUT[22]) );
  DFFS_X1 \reg_mem_reg[21]  ( .D(n86), .CK(CLK), .SN(n18), .Q(DOUT[21]) );
  DFFS_X1 \reg_mem_reg[20]  ( .D(n85), .CK(CLK), .SN(n18), .Q(DOUT[20]) );
  DFFS_X1 \reg_mem_reg[19]  ( .D(n84), .CK(CLK), .SN(n18), .Q(DOUT[19]) );
  DFFS_X1 \reg_mem_reg[18]  ( .D(n83), .CK(CLK), .SN(n18), .Q(DOUT[18]) );
  DFFS_X1 \reg_mem_reg[17]  ( .D(n82), .CK(CLK), .SN(n18), .Q(DOUT[17]) );
  DFFS_X1 \reg_mem_reg[16]  ( .D(n81), .CK(CLK), .SN(n18), .Q(DOUT[16]) );
  DFFS_X1 \reg_mem_reg[15]  ( .D(n80), .CK(CLK), .SN(n18), .Q(DOUT[15]), .QN(
        n48) );
  DFFS_X1 \reg_mem_reg[14]  ( .D(n79), .CK(CLK), .SN(n18), .Q(DOUT[14]), .QN(
        n47) );
  DFFS_X1 \reg_mem_reg[13]  ( .D(n78), .CK(CLK), .SN(n18), .Q(DOUT[13]), .QN(
        n46) );
  DFFS_X1 \reg_mem_reg[12]  ( .D(n77), .CK(CLK), .SN(n17), .Q(DOUT[12]), .QN(
        n45) );
  DFFS_X1 \reg_mem_reg[11]  ( .D(n76), .CK(CLK), .SN(n17), .Q(DOUT[11]), .QN(
        n44) );
  DFFS_X1 \reg_mem_reg[10]  ( .D(n75), .CK(CLK), .SN(n17), .Q(DOUT[10]), .QN(
        n43) );
  DFFS_X1 \reg_mem_reg[9]  ( .D(n74), .CK(CLK), .SN(n17), .Q(DOUT[9]), .QN(n42) );
  DFFS_X1 \reg_mem_reg[8]  ( .D(n73), .CK(CLK), .SN(n17), .Q(DOUT[8]), .QN(n41) );
  DFFS_X1 \reg_mem_reg[7]  ( .D(n72), .CK(CLK), .SN(n17), .Q(DOUT[7]), .QN(n40) );
  DFFS_X1 \reg_mem_reg[6]  ( .D(n71), .CK(CLK), .SN(n17), .Q(DOUT[6]), .QN(n39) );
  DFFS_X1 \reg_mem_reg[5]  ( .D(n70), .CK(CLK), .SN(n17), .Q(DOUT[5]), .QN(n38) );
  DFFS_X1 \reg_mem_reg[4]  ( .D(n69), .CK(CLK), .SN(n17), .Q(DOUT[4]), .QN(n37) );
  DFFS_X1 \reg_mem_reg[3]  ( .D(n68), .CK(CLK), .SN(n17), .Q(DOUT[3]), .QN(n36) );
  DFFS_X1 \reg_mem_reg[2]  ( .D(n67), .CK(CLK), .SN(n17), .Q(DOUT[2]), .QN(n35) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n66), .CK(CLK), .RN(n17), .Q(DOUT[1]), .QN(n34) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n65), .CK(CLK), .RN(n17), .Q(DOUT[0]), .QN(n33) );
  BUF_X1 U2 ( .A(RST_AN), .Z(n17) );
  BUF_X1 U3 ( .A(RST_AN), .Z(n18) );
  BUF_X1 U4 ( .A(RST_AN), .Z(n19) );
  OAI21_X1 U5 ( .B1(n33), .B2(EN), .A(n1), .ZN(n65) );
  NAND2_X1 U6 ( .A1(EN), .A2(DIN[0]), .ZN(n1) );
  OAI21_X1 U7 ( .B1(n40), .B2(EN), .A(n8), .ZN(n72) );
  NAND2_X1 U8 ( .A1(DIN[7]), .A2(EN), .ZN(n8) );
  OAI21_X1 U9 ( .B1(n43), .B2(EN), .A(n11), .ZN(n75) );
  NAND2_X1 U10 ( .A1(DIN[10]), .A2(EN), .ZN(n11) );
  OAI21_X1 U11 ( .B1(n44), .B2(EN), .A(n12), .ZN(n76) );
  NAND2_X1 U12 ( .A1(DIN[11]), .A2(EN), .ZN(n12) );
  OAI21_X1 U13 ( .B1(n46), .B2(EN), .A(n14), .ZN(n78) );
  NAND2_X1 U14 ( .A1(DIN[13]), .A2(EN), .ZN(n14) );
  OAI21_X1 U15 ( .B1(n47), .B2(EN), .A(n15), .ZN(n79) );
  NAND2_X1 U16 ( .A1(DIN[14]), .A2(EN), .ZN(n15) );
  OAI21_X1 U17 ( .B1(n48), .B2(EN), .A(n16), .ZN(n80) );
  NAND2_X1 U18 ( .A1(DIN[15]), .A2(EN), .ZN(n16) );
  OAI21_X1 U19 ( .B1(n37), .B2(EN), .A(n5), .ZN(n69) );
  NAND2_X1 U20 ( .A1(DIN[4]), .A2(EN), .ZN(n5) );
  OAI21_X1 U21 ( .B1(n38), .B2(EN), .A(n6), .ZN(n70) );
  NAND2_X1 U22 ( .A1(DIN[5]), .A2(EN), .ZN(n6) );
  OAI21_X1 U23 ( .B1(n39), .B2(EN), .A(n7), .ZN(n71) );
  NAND2_X1 U24 ( .A1(DIN[6]), .A2(EN), .ZN(n7) );
  OAI21_X1 U25 ( .B1(n41), .B2(EN), .A(n9), .ZN(n73) );
  NAND2_X1 U26 ( .A1(DIN[8]), .A2(EN), .ZN(n9) );
  OAI21_X1 U27 ( .B1(n42), .B2(EN), .A(n10), .ZN(n74) );
  NAND2_X1 U28 ( .A1(DIN[9]), .A2(EN), .ZN(n10) );
  OAI21_X1 U29 ( .B1(n45), .B2(EN), .A(n13), .ZN(n77) );
  NAND2_X1 U30 ( .A1(DIN[12]), .A2(EN), .ZN(n13) );
  OAI21_X1 U31 ( .B1(n64), .B2(EN), .A(n32), .ZN(n96) );
  NAND2_X1 U32 ( .A1(DIN[31]), .A2(EN), .ZN(n32) );
  OAI21_X1 U33 ( .B1(n34), .B2(EN), .A(n2), .ZN(n66) );
  NAND2_X1 U34 ( .A1(DIN[1]), .A2(EN), .ZN(n2) );
  OAI21_X1 U35 ( .B1(n35), .B2(EN), .A(n3), .ZN(n67) );
  NAND2_X1 U36 ( .A1(DIN[2]), .A2(EN), .ZN(n3) );
  OAI21_X1 U37 ( .B1(n36), .B2(EN), .A(n4), .ZN(n68) );
  NAND2_X1 U38 ( .A1(DIN[3]), .A2(EN), .ZN(n4) );
  MUX2_X1 U39 ( .A(DOUT[16]), .B(DIN[16]), .S(EN), .Z(n81) );
  MUX2_X1 U40 ( .A(DOUT[17]), .B(DIN[17]), .S(EN), .Z(n82) );
  MUX2_X1 U41 ( .A(DOUT[18]), .B(DIN[18]), .S(EN), .Z(n83) );
  MUX2_X1 U42 ( .A(DOUT[19]), .B(DIN[19]), .S(EN), .Z(n84) );
  MUX2_X1 U43 ( .A(DOUT[20]), .B(DIN[20]), .S(EN), .Z(n85) );
  MUX2_X1 U44 ( .A(DOUT[21]), .B(DIN[21]), .S(EN), .Z(n86) );
  MUX2_X1 U45 ( .A(DOUT[22]), .B(DIN[22]), .S(EN), .Z(n87) );
  MUX2_X1 U46 ( .A(DOUT[23]), .B(DIN[23]), .S(EN), .Z(n88) );
  MUX2_X1 U47 ( .A(DOUT[24]), .B(DIN[24]), .S(EN), .Z(n89) );
  MUX2_X1 U48 ( .A(DOUT[25]), .B(DIN[25]), .S(EN), .Z(n90) );
  MUX2_X1 U49 ( .A(DOUT[26]), .B(DIN[26]), .S(EN), .Z(n91) );
  MUX2_X1 U50 ( .A(DOUT[27]), .B(DIN[27]), .S(EN), .Z(n92) );
  MUX2_X1 U51 ( .A(DOUT[28]), .B(DIN[28]), .S(EN), .Z(n93) );
  MUX2_X1 U52 ( .A(DOUT[29]), .B(DIN[29]), .S(EN), .Z(n94) );
  MUX2_X1 U53 ( .A(DOUT[30]), .B(DIN[30]), .S(EN), .Z(n95) );
endmodule


module REG_PIPO_32_00000000_00000000_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n99,
         n100, n101, n102;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n98), .CK(CLK), .RN(n4), .Q(DOUT[31]), .QN(
        n66) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n97), .CK(CLK), .RN(n4), .Q(DOUT[30]), .QN(
        n65) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n96), .CK(CLK), .RN(n4), .Q(DOUT[29]), .QN(
        n64) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n95), .CK(CLK), .RN(n4), .Q(DOUT[28]), .QN(
        n63) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n94), .CK(CLK), .RN(n4), .Q(DOUT[27]), .QN(
        n62) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n93), .CK(CLK), .RN(n4), .Q(DOUT[26]), .QN(
        n61) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n92), .CK(CLK), .RN(n4), .Q(DOUT[25]), .QN(
        n60) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n91), .CK(CLK), .RN(n4), .Q(DOUT[24]), .QN(
        n59) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n90), .CK(CLK), .RN(n4), .Q(DOUT[23]), .QN(
        n58) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n89), .CK(CLK), .RN(n4), .Q(DOUT[22]), .QN(
        n57) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n88), .CK(CLK), .RN(n3), .Q(DOUT[21]), .QN(
        n56) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n87), .CK(CLK), .RN(n3), .Q(DOUT[20]), .QN(
        n55) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n86), .CK(CLK), .RN(n3), .Q(DOUT[19]), .QN(
        n54) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n85), .CK(CLK), .RN(n3), .Q(DOUT[18]), .QN(
        n53) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n84), .CK(CLK), .RN(n3), .Q(DOUT[17]), .QN(
        n52) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n83), .CK(CLK), .RN(n3), .Q(DOUT[16]), .QN(
        n51) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n82), .CK(CLK), .RN(n3), .Q(DOUT[15]), .QN(
        n50) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n81), .CK(CLK), .RN(n3), .Q(DOUT[14]), .QN(
        n49) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n80), .CK(CLK), .RN(n3), .Q(DOUT[13]), .QN(
        n48) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n79), .CK(CLK), .RN(n3), .Q(DOUT[12]), .QN(
        n47) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n78), .CK(CLK), .RN(n3), .Q(DOUT[11]), .QN(
        n46) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n77), .CK(CLK), .RN(n2), .Q(DOUT[10]), .QN(
        n45) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n76), .CK(CLK), .RN(n2), .Q(DOUT[9]), .QN(n44)
         );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n75), .CK(CLK), .RN(n2), .Q(DOUT[8]), .QN(n43)
         );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n74), .CK(CLK), .RN(n2), .Q(DOUT[7]), .QN(n42)
         );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n73), .CK(CLK), .RN(n2), .Q(DOUT[6]), .QN(n41)
         );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n72), .CK(CLK), .RN(n2), .Q(DOUT[5]), .QN(n40)
         );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n71), .CK(CLK), .RN(n2), .Q(DOUT[4]), .QN(n39)
         );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n70), .CK(CLK), .RN(n2), .Q(DOUT[3]), .QN(n38)
         );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n69), .CK(CLK), .RN(n2), .Q(DOUT[2]), .QN(n37)
         );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n68), .CK(CLK), .RN(n2), .Q(DOUT[1]), .QN(n36)
         );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n67), .CK(CLK), .RN(n2), .Q(DOUT[0]), .QN(n35)
         );
  BUF_X1 U2 ( .A(RST_AN), .Z(n2) );
  BUF_X1 U3 ( .A(RST_AN), .Z(n3) );
  BUF_X1 U4 ( .A(RST_AN), .Z(n4) );
  OAI22_X1 U5 ( .A1(n35), .A2(EN), .B1(n1), .B2(n101), .ZN(n67) );
  INV_X1 U6 ( .A(DIN[0]), .ZN(n101) );
  OAI22_X1 U7 ( .A1(n36), .A2(EN), .B1(n1), .B2(n100), .ZN(n68) );
  INV_X1 U8 ( .A(DIN[1]), .ZN(n100) );
  OAI22_X1 U9 ( .A1(n37), .A2(EN), .B1(n1), .B2(n99), .ZN(n69) );
  INV_X1 U10 ( .A(DIN[2]), .ZN(n99) );
  OAI22_X1 U11 ( .A1(n38), .A2(EN), .B1(n1), .B2(n34), .ZN(n70) );
  INV_X1 U12 ( .A(DIN[3]), .ZN(n34) );
  OAI22_X1 U13 ( .A1(n39), .A2(EN), .B1(n1), .B2(n33), .ZN(n71) );
  INV_X1 U14 ( .A(DIN[4]), .ZN(n33) );
  OAI22_X1 U15 ( .A1(n40), .A2(EN), .B1(n1), .B2(n32), .ZN(n72) );
  INV_X1 U16 ( .A(DIN[5]), .ZN(n32) );
  OAI22_X1 U17 ( .A1(n41), .A2(EN), .B1(n1), .B2(n31), .ZN(n73) );
  INV_X1 U18 ( .A(DIN[6]), .ZN(n31) );
  OAI22_X1 U19 ( .A1(n42), .A2(EN), .B1(n1), .B2(n30), .ZN(n74) );
  INV_X1 U20 ( .A(DIN[7]), .ZN(n30) );
  OAI22_X1 U21 ( .A1(n43), .A2(EN), .B1(n1), .B2(n29), .ZN(n75) );
  INV_X1 U22 ( .A(DIN[8]), .ZN(n29) );
  OAI22_X1 U23 ( .A1(n44), .A2(EN), .B1(n1), .B2(n28), .ZN(n76) );
  INV_X1 U24 ( .A(DIN[9]), .ZN(n28) );
  OAI22_X1 U25 ( .A1(n45), .A2(EN), .B1(n1), .B2(n27), .ZN(n77) );
  INV_X1 U26 ( .A(DIN[10]), .ZN(n27) );
  OAI22_X1 U27 ( .A1(n46), .A2(EN), .B1(n1), .B2(n26), .ZN(n78) );
  INV_X1 U28 ( .A(DIN[11]), .ZN(n26) );
  OAI22_X1 U29 ( .A1(n47), .A2(EN), .B1(n1), .B2(n25), .ZN(n79) );
  INV_X1 U30 ( .A(DIN[12]), .ZN(n25) );
  OAI22_X1 U31 ( .A1(n48), .A2(EN), .B1(n1), .B2(n24), .ZN(n80) );
  INV_X1 U32 ( .A(DIN[13]), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n49), .A2(EN), .B1(n1), .B2(n23), .ZN(n81) );
  INV_X1 U34 ( .A(DIN[14]), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n50), .A2(EN), .B1(n1), .B2(n22), .ZN(n82) );
  INV_X1 U36 ( .A(DIN[15]), .ZN(n22) );
  OAI22_X1 U37 ( .A1(n66), .A2(EN), .B1(n1), .B2(n102), .ZN(n98) );
  INV_X1 U38 ( .A(DIN[31]), .ZN(n102) );
  INV_X1 U39 ( .A(EN), .ZN(n5) );
  OR2_X1 U40 ( .A1(INIT), .A2(n5), .ZN(n1) );
  INV_X1 U41 ( .A(n1), .ZN(n20) );
  NAND2_X1 U42 ( .A1(DIN[16]), .A2(n20), .ZN(n6) );
  OAI21_X1 U43 ( .B1(n51), .B2(EN), .A(n6), .ZN(n83) );
  NAND2_X1 U44 ( .A1(DIN[17]), .A2(n20), .ZN(n7) );
  OAI21_X1 U45 ( .B1(n52), .B2(EN), .A(n7), .ZN(n84) );
  NAND2_X1 U46 ( .A1(DIN[18]), .A2(n20), .ZN(n8) );
  OAI21_X1 U47 ( .B1(n53), .B2(EN), .A(n8), .ZN(n85) );
  NAND2_X1 U48 ( .A1(DIN[19]), .A2(n20), .ZN(n9) );
  OAI21_X1 U49 ( .B1(n54), .B2(EN), .A(n9), .ZN(n86) );
  NAND2_X1 U50 ( .A1(DIN[20]), .A2(n20), .ZN(n10) );
  OAI21_X1 U51 ( .B1(n55), .B2(EN), .A(n10), .ZN(n87) );
  NAND2_X1 U52 ( .A1(DIN[21]), .A2(n20), .ZN(n11) );
  OAI21_X1 U53 ( .B1(n56), .B2(EN), .A(n11), .ZN(n88) );
  NAND2_X1 U54 ( .A1(DIN[22]), .A2(n20), .ZN(n12) );
  OAI21_X1 U55 ( .B1(n57), .B2(EN), .A(n12), .ZN(n89) );
  NAND2_X1 U56 ( .A1(DIN[23]), .A2(n20), .ZN(n13) );
  OAI21_X1 U57 ( .B1(n58), .B2(EN), .A(n13), .ZN(n90) );
  NAND2_X1 U58 ( .A1(DIN[24]), .A2(n20), .ZN(n14) );
  OAI21_X1 U59 ( .B1(n59), .B2(EN), .A(n14), .ZN(n91) );
  NAND2_X1 U60 ( .A1(DIN[25]), .A2(n20), .ZN(n15) );
  OAI21_X1 U61 ( .B1(n60), .B2(EN), .A(n15), .ZN(n92) );
  NAND2_X1 U62 ( .A1(DIN[26]), .A2(n20), .ZN(n16) );
  OAI21_X1 U63 ( .B1(n61), .B2(EN), .A(n16), .ZN(n93) );
  NAND2_X1 U64 ( .A1(DIN[27]), .A2(n20), .ZN(n17) );
  OAI21_X1 U65 ( .B1(n62), .B2(EN), .A(n17), .ZN(n94) );
  NAND2_X1 U66 ( .A1(DIN[28]), .A2(n20), .ZN(n18) );
  OAI21_X1 U67 ( .B1(n63), .B2(EN), .A(n18), .ZN(n95) );
  NAND2_X1 U68 ( .A1(DIN[29]), .A2(n20), .ZN(n19) );
  OAI21_X1 U69 ( .B1(n64), .B2(EN), .A(n19), .ZN(n96) );
  NAND2_X1 U70 ( .A1(DIN[30]), .A2(n20), .ZN(n21) );
  OAI21_X1 U71 ( .B1(n65), .B2(EN), .A(n21), .ZN(n97) );
endmodule


module REG_PIPO_32_00000000_00000000_11 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module RF_ADDR_W5_DATA_W32 ( CLK, RST_AN, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST_AN, ENABLE, RD1, RD2, WR;
  wire   \registers[1][31] , \registers[1][30] , \registers[1][29] ,
         \registers[1][28] , \registers[1][27] , \registers[1][26] ,
         \registers[1][25] , \registers[1][24] , \registers[1][23] ,
         \registers[1][22] , \registers[1][21] , \registers[1][20] ,
         \registers[1][19] , \registers[1][18] , \registers[1][17] ,
         \registers[1][16] , \registers[1][15] , \registers[1][14] ,
         \registers[1][13] , \registers[1][12] , \registers[1][11] ,
         \registers[1][10] , \registers[1][9] , \registers[1][8] ,
         \registers[1][7] , \registers[1][6] , \registers[1][5] ,
         \registers[1][4] , \registers[1][3] , \registers[1][2] ,
         \registers[1][1] , \registers[1][0] , \registers[6][31] ,
         \registers[6][30] , \registers[6][29] , \registers[6][28] ,
         \registers[6][27] , \registers[6][26] , \registers[6][25] ,
         \registers[6][24] , \registers[6][23] , \registers[6][22] ,
         \registers[6][21] , \registers[6][20] , \registers[6][19] ,
         \registers[6][18] , \registers[6][17] , \registers[6][16] ,
         \registers[6][15] , \registers[6][14] , \registers[6][13] ,
         \registers[6][12] , \registers[6][11] , \registers[6][10] ,
         \registers[6][9] , \registers[6][8] , \registers[6][7] ,
         \registers[6][6] , \registers[6][5] , \registers[6][4] ,
         \registers[6][3] , \registers[6][2] , \registers[6][1] ,
         \registers[6][0] , \registers[7][31] , \registers[7][30] ,
         \registers[7][29] , \registers[7][28] , \registers[7][27] ,
         \registers[7][26] , \registers[7][25] , \registers[7][24] ,
         \registers[7][23] , \registers[7][22] , \registers[7][21] ,
         \registers[7][20] , \registers[7][19] , \registers[7][18] ,
         \registers[7][17] , \registers[7][16] , \registers[7][15] ,
         \registers[7][14] , \registers[7][13] , \registers[7][12] ,
         \registers[7][11] , \registers[7][10] , \registers[7][9] ,
         \registers[7][8] , \registers[7][7] , \registers[7][6] ,
         \registers[7][5] , \registers[7][4] , \registers[7][3] ,
         \registers[7][2] , \registers[7][1] , \registers[7][0] ,
         \registers[8][31] , \registers[8][30] , \registers[8][29] ,
         \registers[8][28] , \registers[8][27] , \registers[8][26] ,
         \registers[8][25] , \registers[8][24] , \registers[8][23] ,
         \registers[8][22] , \registers[8][21] , \registers[8][20] ,
         \registers[8][19] , \registers[8][18] , \registers[8][17] ,
         \registers[8][16] , \registers[8][15] , \registers[8][14] ,
         \registers[8][13] , \registers[8][12] , \registers[8][11] ,
         \registers[8][10] , \registers[8][9] , \registers[8][8] ,
         \registers[8][7] , \registers[8][6] , \registers[8][5] ,
         \registers[8][4] , \registers[8][3] , \registers[8][2] ,
         \registers[8][1] , \registers[8][0] , \registers[9][31] ,
         \registers[9][30] , \registers[9][29] , \registers[9][28] ,
         \registers[9][27] , \registers[9][26] , \registers[9][25] ,
         \registers[9][24] , \registers[9][23] , \registers[9][22] ,
         \registers[9][21] , \registers[9][20] , \registers[9][19] ,
         \registers[9][18] , \registers[9][17] , \registers[9][16] ,
         \registers[9][15] , \registers[9][14] , \registers[9][13] ,
         \registers[9][12] , \registers[9][11] , \registers[9][10] ,
         \registers[9][9] , \registers[9][8] , \registers[9][7] ,
         \registers[9][6] , \registers[9][5] , \registers[9][4] ,
         \registers[9][3] , \registers[9][2] , \registers[9][1] ,
         \registers[9][0] , \registers[12][31] , \registers[12][30] ,
         \registers[12][29] , \registers[12][28] , \registers[12][27] ,
         \registers[12][26] , \registers[12][25] , \registers[12][24] ,
         \registers[12][23] , \registers[12][22] , \registers[12][21] ,
         \registers[12][20] , \registers[12][19] , \registers[12][18] ,
         \registers[12][17] , \registers[12][16] , \registers[12][15] ,
         \registers[12][14] , \registers[12][13] , \registers[12][12] ,
         \registers[12][11] , \registers[12][10] , \registers[12][9] ,
         \registers[12][8] , \registers[12][7] , \registers[12][6] ,
         \registers[12][5] , \registers[12][4] , \registers[12][3] ,
         \registers[12][2] , \registers[12][1] , \registers[12][0] ,
         \registers[13][31] , \registers[13][30] , \registers[13][29] ,
         \registers[13][28] , \registers[13][27] , \registers[13][26] ,
         \registers[13][25] , \registers[13][24] , \registers[13][23] ,
         \registers[13][22] , \registers[13][21] , \registers[13][20] ,
         \registers[13][19] , \registers[13][18] , \registers[13][17] ,
         \registers[13][16] , \registers[13][15] , \registers[13][14] ,
         \registers[13][13] , \registers[13][12] , \registers[13][11] ,
         \registers[13][10] , \registers[13][9] , \registers[13][8] ,
         \registers[13][7] , \registers[13][6] , \registers[13][5] ,
         \registers[13][4] , \registers[13][3] , \registers[13][2] ,
         \registers[13][1] , \registers[13][0] , \registers[18][31] ,
         \registers[18][30] , \registers[18][29] , \registers[18][28] ,
         \registers[18][27] , \registers[18][26] , \registers[18][25] ,
         \registers[18][24] , \registers[18][23] , \registers[18][22] ,
         \registers[18][21] , \registers[18][20] , \registers[18][19] ,
         \registers[18][18] , \registers[18][17] , \registers[18][16] ,
         \registers[18][15] , \registers[18][14] , \registers[18][13] ,
         \registers[18][12] , \registers[18][11] , \registers[18][10] ,
         \registers[18][9] , \registers[18][8] , \registers[18][7] ,
         \registers[18][6] , \registers[18][5] , \registers[18][4] ,
         \registers[18][3] , \registers[18][2] , \registers[18][1] ,
         \registers[18][0] , \registers[19][31] , \registers[19][30] ,
         \registers[19][29] , \registers[19][28] , \registers[19][27] ,
         \registers[19][26] , \registers[19][25] , \registers[19][24] ,
         \registers[19][23] , \registers[19][22] , \registers[19][21] ,
         \registers[19][20] , \registers[19][19] , \registers[19][18] ,
         \registers[19][17] , \registers[19][16] , \registers[19][15] ,
         \registers[19][14] , \registers[19][13] , \registers[19][12] ,
         \registers[19][11] , \registers[19][10] , \registers[19][9] ,
         \registers[19][8] , \registers[19][7] , \registers[19][6] ,
         \registers[19][5] , \registers[19][4] , \registers[19][3] ,
         \registers[19][2] , \registers[19][1] , \registers[19][0] ,
         \registers[22][31] , \registers[22][30] , \registers[22][29] ,
         \registers[22][28] , \registers[22][27] , \registers[22][26] ,
         \registers[22][25] , \registers[22][24] , \registers[22][23] ,
         \registers[22][22] , \registers[22][21] , \registers[22][20] ,
         \registers[22][19] , \registers[22][18] , \registers[22][17] ,
         \registers[22][16] , \registers[22][15] , \registers[22][14] ,
         \registers[22][13] , \registers[22][12] , \registers[22][11] ,
         \registers[22][10] , \registers[22][9] , \registers[22][8] ,
         \registers[22][7] , \registers[22][6] , \registers[22][5] ,
         \registers[22][4] , \registers[22][3] , \registers[22][2] ,
         \registers[22][1] , \registers[22][0] , \registers[23][31] ,
         \registers[23][30] , \registers[23][29] , \registers[23][28] ,
         \registers[23][27] , \registers[23][26] , \registers[23][25] ,
         \registers[23][24] , \registers[23][23] , \registers[23][22] ,
         \registers[23][21] , \registers[23][20] , \registers[23][19] ,
         \registers[23][18] , \registers[23][17] , \registers[23][16] ,
         \registers[23][15] , \registers[23][14] , \registers[23][13] ,
         \registers[23][12] , \registers[23][11] , \registers[23][10] ,
         \registers[23][9] , \registers[23][8] , \registers[23][7] ,
         \registers[23][6] , \registers[23][5] , \registers[23][4] ,
         \registers[23][3] , \registers[23][2] , \registers[23][1] ,
         \registers[23][0] , \registers[24][31] , \registers[24][30] ,
         \registers[24][29] , \registers[24][28] , \registers[24][27] ,
         \registers[24][26] , \registers[24][25] , \registers[24][24] ,
         \registers[24][23] , \registers[24][22] , \registers[24][21] ,
         \registers[24][20] , \registers[24][19] , \registers[24][18] ,
         \registers[24][17] , \registers[24][16] , \registers[24][15] ,
         \registers[24][14] , \registers[24][13] , \registers[24][12] ,
         \registers[24][11] , \registers[24][10] , \registers[24][9] ,
         \registers[24][8] , \registers[24][7] , \registers[24][6] ,
         \registers[24][5] , \registers[24][4] , \registers[24][3] ,
         \registers[24][2] , \registers[24][1] , \registers[24][0] ,
         \registers[25][31] , \registers[25][30] , \registers[25][29] ,
         \registers[25][28] , \registers[25][27] , \registers[25][26] ,
         \registers[25][25] , \registers[25][24] , \registers[25][23] ,
         \registers[25][22] , \registers[25][21] , \registers[25][20] ,
         \registers[25][19] , \registers[25][18] , \registers[25][17] ,
         \registers[25][16] , \registers[25][15] , \registers[25][14] ,
         \registers[25][13] , \registers[25][12] , \registers[25][11] ,
         \registers[25][10] , \registers[25][9] , \registers[25][8] ,
         \registers[25][7] , \registers[25][6] , \registers[25][5] ,
         \registers[25][4] , \registers[25][3] , \registers[25][2] ,
         \registers[25][1] , \registers[25][0] , \registers[28][31] ,
         \registers[28][30] , \registers[28][29] , \registers[28][28] ,
         \registers[28][27] , \registers[28][26] , \registers[28][25] ,
         \registers[28][24] , \registers[28][23] , \registers[28][22] ,
         \registers[28][21] , \registers[28][20] , \registers[28][19] ,
         \registers[28][18] , \registers[28][17] , \registers[28][16] ,
         \registers[28][15] , \registers[28][14] , \registers[28][13] ,
         \registers[28][12] , \registers[28][11] , \registers[28][10] ,
         \registers[28][9] , \registers[28][8] , \registers[28][7] ,
         \registers[28][6] , \registers[28][5] , \registers[28][4] ,
         \registers[28][3] , \registers[28][2] , \registers[28][1] ,
         \registers[28][0] , \registers[29][31] , \registers[29][30] ,
         \registers[29][29] , \registers[29][28] , \registers[29][27] ,
         \registers[29][26] , \registers[29][25] , \registers[29][24] ,
         \registers[29][23] , \registers[29][22] , \registers[29][21] ,
         \registers[29][20] , \registers[29][19] , \registers[29][18] ,
         \registers[29][17] , \registers[29][16] , \registers[29][15] ,
         \registers[29][14] , \registers[29][13] , \registers[29][12] ,
         \registers[29][11] , \registers[29][10] , \registers[29][9] ,
         \registers[29][8] , \registers[29][7] , \registers[29][6] ,
         \registers[29][5] , \registers[29][4] , \registers[29][3] ,
         \registers[29][2] , \registers[29][1] , \registers[29][0] , N83, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n1068, n1069, n1070, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1142, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1202, n1203,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1270, n1272, n1273, n1274, n1275, n1276, n1278, n1279, n1280,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1350, n1351, n1352,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, net17879, net18066,
         net26249, net26247, net26245, net26243, net26429, net26427, net26425,
         net26423, net26421, net26419, net26417, net26415, net26413, net26597,
         net26595, net26593, net26591, net26589, net26585, net26583, net26581,
         net26579, net26747, net26745, net26743, net26753, net26751, net26749,
         net26933, net26931, net26929, net26939, net26937, net26935, net28529,
         net28528, net33812, net38912, net38974, net38973, net38972, net38971,
         net38970, net38969, net38968, net38967, net38966, net38965, net38964,
         net38993, net38992, net39055, net39090, net39089, net39096, net44304,
         net44303, net44322, net44474, net44473, net44605, net44604, net44818,
         net44860, n1277, n1249, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1071, n1098, n1115, n1141,
         n1143, n1201, n1204, n1218, n1261, n1269, n1271, n1281, n1349, n1353,
         n1370, n1400, n1421, n1437, n1474, n1538, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272;

  DFFR_X1 \registers_reg[1][29]  ( .D(n3919), .CK(n4272), .RN(n3748), .Q(
        \registers[1][29] ) );
  DFFR_X1 \registers_reg[1][28]  ( .D(n3918), .CK(n4272), .RN(n3748), .Q(
        \registers[1][28] ) );
  DFFR_X1 \registers_reg[1][26]  ( .D(n3916), .CK(n4272), .RN(n3748), .Q(
        \registers[1][26] ) );
  DFFR_X1 \registers_reg[1][25]  ( .D(n3915), .CK(n4272), .RN(n3748), .Q(
        \registers[1][25] ) );
  DFFR_X1 \registers_reg[1][23]  ( .D(n3913), .CK(n4272), .RN(n3748), .Q(
        \registers[1][23] ) );
  DFFR_X1 \registers_reg[1][22]  ( .D(n3912), .CK(n4272), .RN(n3748), .Q(
        \registers[1][22] ) );
  DFFR_X1 \registers_reg[1][21]  ( .D(n3911), .CK(n4272), .RN(n3748), .Q(
        \registers[1][21] ) );
  DFFR_X1 \registers_reg[1][20]  ( .D(n3910), .CK(n4272), .RN(n3748), .Q(
        \registers[1][20] ) );
  DFFR_X1 \registers_reg[1][18]  ( .D(n3908), .CK(n4272), .RN(n3747), .Q(
        \registers[1][18] ) );
  DFFR_X1 \registers_reg[1][17]  ( .D(n3907), .CK(n4272), .RN(n3747), .Q(
        \registers[1][17] ) );
  DFFR_X1 \registers_reg[1][16]  ( .D(n3906), .CK(n4272), .RN(n3747), .Q(
        \registers[1][16] ) );
  DFFR_X1 \registers_reg[1][13]  ( .D(n3903), .CK(n4272), .RN(n3747), .Q(
        \registers[1][13] ) );
  DFFR_X1 \registers_reg[1][9]  ( .D(n3899), .CK(n4272), .RN(n3747), .Q(
        \registers[1][9] ) );
  DFFR_X1 \registers_reg[1][6]  ( .D(n3896), .CK(n4272), .RN(n3746), .Q(
        \registers[1][6] ) );
  DFFR_X1 \registers_reg[1][5]  ( .D(n3895), .CK(n4272), .RN(n3746), .Q(
        \registers[1][5] ) );
  DFFR_X1 \registers_reg[1][4]  ( .D(n3894), .CK(n4272), .RN(n3746), .Q(
        \registers[1][4] ) );
  DFFR_X1 \registers_reg[1][2]  ( .D(n3892), .CK(n4272), .RN(n3746), .Q(
        \registers[1][2] ) );
  DFFR_X1 \registers_reg[1][1]  ( .D(n3891), .CK(n4272), .RN(n3746), .Q(
        \registers[1][1] ) );
  DFFR_X1 \registers_reg[1][0]  ( .D(n3890), .CK(n4272), .RN(n3746), .Q(
        \registers[1][0] ) );
  DFFR_X1 \registers_reg[2][22]  ( .D(n3276), .CK(n4272), .RN(n3745), .QN(n42)
         );
  DFFR_X1 \registers_reg[2][7]  ( .D(n3261), .CK(n4272), .RN(n3744), .QN(n57)
         );
  DFFR_X1 \registers_reg[3][22]  ( .D(n3244), .CK(n4272), .RN(n3742), .QN(n74)
         );
  DFFR_X1 \registers_reg[3][12]  ( .D(n3234), .CK(n4272), .RN(n3741), .QN(n84)
         );
  DFFR_X1 \registers_reg[3][7]  ( .D(n3229), .CK(n4272), .RN(n3741), .QN(n89)
         );
  DFFR_X1 \registers_reg[4][31]  ( .D(n3221), .CK(n4272), .RN(n3740), .QN(n97)
         );
  DFFR_X1 \registers_reg[4][30]  ( .D(n3220), .CK(n4272), .RN(n3740), .QN(n98)
         );
  DFFR_X1 \registers_reg[4][29]  ( .D(n3219), .CK(n4272), .RN(n3740), .QN(n99)
         );
  DFFR_X1 \registers_reg[4][28]  ( .D(n3218), .CK(n4272), .RN(n3740), .QN(n100) );
  DFFR_X1 \registers_reg[4][26]  ( .D(n3216), .CK(n4272), .RN(n3739), .QN(n102) );
  DFFR_X1 \registers_reg[4][25]  ( .D(n3215), .CK(n4272), .RN(n3739), .QN(n103) );
  DFFR_X1 \registers_reg[4][24]  ( .D(n3214), .CK(n4272), .RN(n3739), .QN(n104) );
  DFFR_X1 \registers_reg[4][22]  ( .D(n3212), .CK(n4272), .RN(n3739), .QN(n106) );
  DFFR_X1 \registers_reg[4][21]  ( .D(n3211), .CK(n4272), .RN(n3739), .QN(n107) );
  DFFR_X1 \registers_reg[4][20]  ( .D(n3210), .CK(n4272), .RN(n3739), .QN(n108) );
  DFFR_X1 \registers_reg[4][19]  ( .D(n3209), .CK(n4272), .RN(n3739), .QN(n109) );
  DFFR_X1 \registers_reg[4][17]  ( .D(n3207), .CK(n4272), .RN(n3739), .QN(n111) );
  DFFR_X1 \registers_reg[4][16]  ( .D(n3206), .CK(n4272), .RN(n3739), .QN(n112) );
  DFFR_X1 \registers_reg[4][15]  ( .D(n3205), .CK(n4272), .RN(n3738), .QN(n113) );
  DFFR_X1 \registers_reg[4][14]  ( .D(n3204), .CK(n4272), .RN(n3738), .QN(n114) );
  DFFR_X1 \registers_reg[4][12]  ( .D(n3202), .CK(n4272), .RN(n3738), .QN(n116) );
  DFFR_X1 \registers_reg[4][11]  ( .D(n3201), .CK(n4272), .RN(n3738), .QN(n117) );
  DFFR_X1 \registers_reg[4][10]  ( .D(n3200), .CK(n4272), .RN(n3738), .QN(n118) );
  DFFR_X1 \registers_reg[4][9]  ( .D(n3199), .CK(n4272), .RN(n3738), .QN(n119)
         );
  DFFR_X1 \registers_reg[4][7]  ( .D(n3197), .CK(n4272), .RN(n3738), .QN(n121)
         );
  DFFR_X1 \registers_reg[4][6]  ( .D(n3196), .CK(n4272), .RN(n3738), .QN(n122)
         );
  DFFR_X1 \registers_reg[4][5]  ( .D(n3195), .CK(n4272), .RN(n3738), .QN(n123)
         );
  DFFR_X1 \registers_reg[4][4]  ( .D(n3194), .CK(n4272), .RN(n3737), .QN(n124)
         );
  DFFR_X1 \registers_reg[4][3]  ( .D(n3193), .CK(n4272), .RN(n3737), .QN(n125)
         );
  DFFR_X1 \registers_reg[4][2]  ( .D(n3192), .CK(n4272), .RN(n3737), .QN(n126)
         );
  DFFR_X1 \registers_reg[4][1]  ( .D(n3191), .CK(n4272), .RN(n3737), .QN(n127)
         );
  DFFR_X1 \registers_reg[4][0]  ( .D(n3190), .CK(n4272), .RN(n3737), .QN(n128)
         );
  DFFR_X1 \registers_reg[5][22]  ( .D(n3180), .CK(n4272), .RN(n3736), .QN(n138) );
  DFFR_X1 \registers_reg[5][17]  ( .D(n3175), .CK(n4272), .RN(n3736), .QN(n143) );
  DFFR_X1 \registers_reg[5][7]  ( .D(n3165), .CK(n4272), .RN(n3735), .QN(n153)
         );
  DFFR_X1 \registers_reg[6][7]  ( .D(n3929), .CK(n4272), .RN(n3732), .Q(
        \registers[6][7] ) );
  DFFR_X1 \registers_reg[6][6]  ( .D(n3928), .CK(n4272), .RN(n3732), .Q(
        \registers[6][6] ) );
  DFFR_X1 \registers_reg[6][5]  ( .D(n3927), .CK(n4272), .RN(n3732), .Q(
        \registers[6][5] ) );
  DFFR_X1 \registers_reg[6][4]  ( .D(n3926), .CK(n4272), .RN(n3732), .Q(
        \registers[6][4] ) );
  DFFR_X1 \registers_reg[6][3]  ( .D(n3925), .CK(n4272), .RN(n3732), .Q(
        \registers[6][3] ) );
  DFFR_X1 \registers_reg[6][2]  ( .D(n3924), .CK(n4272), .RN(n3731), .Q(
        \registers[6][2] ) );
  DFFR_X1 \registers_reg[6][1]  ( .D(n3923), .CK(n4272), .RN(n3731), .Q(
        \registers[6][1] ) );
  DFFR_X1 \registers_reg[6][0]  ( .D(n3922), .CK(n4272), .RN(n3731), .Q(
        \registers[6][0] ) );
  DFFR_X1 \registers_reg[7][31]  ( .D(n3984), .CK(n4272), .RN(n3731), .Q(
        \registers[7][31] ) );
  DFFR_X1 \registers_reg[7][30]  ( .D(n3983), .CK(n4272), .RN(n3731), .Q(
        \registers[7][30] ) );
  DFFR_X1 \registers_reg[7][29]  ( .D(n3982), .CK(n4272), .RN(n3731), .Q(
        \registers[7][29] ) );
  DFFR_X1 \registers_reg[7][28]  ( .D(n3981), .CK(n4272), .RN(n3731), .Q(
        \registers[7][28] ) );
  DFFR_X1 \registers_reg[7][27]  ( .D(n3980), .CK(n4272), .RN(n3731), .Q(
        \registers[7][27] ) );
  DFFR_X1 \registers_reg[7][26]  ( .D(n3979), .CK(n4272), .RN(n3731), .Q(
        \registers[7][26] ) );
  DFFR_X1 \registers_reg[7][25]  ( .D(n3978), .CK(n4272), .RN(n3731), .Q(
        \registers[7][25] ) );
  DFFR_X1 \registers_reg[7][23]  ( .D(n3976), .CK(n4272), .RN(n3730), .Q(
        \registers[7][23] ) );
  DFFR_X1 \registers_reg[7][22]  ( .D(n3975), .CK(n4272), .RN(n3730), .Q(
        \registers[7][22] ) );
  DFFR_X1 \registers_reg[7][21]  ( .D(n3974), .CK(n4272), .RN(n3730), .Q(
        \registers[7][21] ) );
  DFFR_X1 \registers_reg[7][20]  ( .D(n3973), .CK(n4272), .RN(n3730), .Q(
        \registers[7][20] ) );
  DFFR_X1 \registers_reg[7][19]  ( .D(n3972), .CK(n4272), .RN(n3730), .Q(
        \registers[7][19] ) );
  DFFR_X1 \registers_reg[7][18]  ( .D(n3971), .CK(n4272), .RN(n3730), .Q(
        \registers[7][18] ) );
  DFFR_X1 \registers_reg[7][17]  ( .D(n3970), .CK(n4272), .RN(n3730), .Q(
        \registers[7][17] ) );
  DFFR_X1 \registers_reg[7][16]  ( .D(n3969), .CK(n4272), .RN(n3730), .Q(
        \registers[7][16] ) );
  DFFR_X1 \registers_reg[7][15]  ( .D(n3968), .CK(n4272), .RN(n3730), .Q(
        \registers[7][15] ) );
  DFFR_X1 \registers_reg[7][14]  ( .D(n3967), .CK(n4272), .RN(n3730), .Q(
        \registers[7][14] ) );
  DFFR_X1 \registers_reg[7][13]  ( .D(n3966), .CK(n4272), .RN(n3730), .Q(
        \registers[7][13] ) );
  DFFR_X1 \registers_reg[7][12]  ( .D(n3965), .CK(n4272), .RN(n3729), .Q(
        \registers[7][12] ) );
  DFFR_X1 \registers_reg[7][11]  ( .D(n3964), .CK(n4272), .RN(n3729), .Q(
        \registers[7][11] ) );
  DFFR_X1 \registers_reg[7][10]  ( .D(n3963), .CK(n4272), .RN(n3729), .Q(
        \registers[7][10] ) );
  DFFR_X1 \registers_reg[7][9]  ( .D(n3962), .CK(n4272), .RN(n3729), .Q(
        \registers[7][9] ) );
  DFFR_X1 \registers_reg[7][8]  ( .D(n3961), .CK(n4272), .RN(n3729), .Q(
        \registers[7][8] ) );
  DFFR_X1 \registers_reg[7][7]  ( .D(n3960), .CK(n4272), .RN(n3729), .Q(
        \registers[7][7] ) );
  DFFR_X1 \registers_reg[7][6]  ( .D(n3959), .CK(n4272), .RN(n3729), .Q(
        \registers[7][6] ) );
  DFFR_X1 \registers_reg[7][5]  ( .D(n3958), .CK(n4272), .RN(n3729), .Q(
        \registers[7][5] ) );
  DFFR_X1 \registers_reg[7][4]  ( .D(n3957), .CK(n4272), .RN(n3729), .Q(
        \registers[7][4] ) );
  DFFR_X1 \registers_reg[7][3]  ( .D(n3956), .CK(n4272), .RN(n3729), .Q(
        \registers[7][3] ) );
  DFFR_X1 \registers_reg[7][2]  ( .D(n3955), .CK(n4272), .RN(n3729), .Q(
        \registers[7][2] ) );
  DFFR_X1 \registers_reg[7][1]  ( .D(n3954), .CK(n4272), .RN(n3728), .Q(
        \registers[7][1] ) );
  DFFR_X1 \registers_reg[7][0]  ( .D(n3953), .CK(n4272), .RN(n3728), .Q(
        \registers[7][0] ) );
  DFFR_X1 \registers_reg[8][31]  ( .D(n3796), .CK(n4272), .RN(n3728), .Q(
        \registers[8][31] ) );
  DFFR_X1 \registers_reg[8][30]  ( .D(n3795), .CK(n4272), .RN(n3728), .Q(
        \registers[8][30] ) );
  DFFR_X1 \registers_reg[8][29]  ( .D(n3794), .CK(n4272), .RN(n3728), .Q(
        \registers[8][29] ) );
  DFFR_X1 \registers_reg[8][28]  ( .D(n3793), .CK(n4272), .RN(n3728), .Q(
        \registers[8][28] ) );
  DFFR_X1 \registers_reg[8][27]  ( .D(n3792), .CK(n4272), .RN(n3728), .Q(
        \registers[8][27] ) );
  DFFR_X1 \registers_reg[8][26]  ( .D(n3791), .CK(n4272), .RN(n3728), .Q(
        \registers[8][26] ) );
  DFFR_X1 \registers_reg[8][25]  ( .D(n3790), .CK(n4272), .RN(n3728), .Q(
        \registers[8][25] ) );
  DFFR_X1 \registers_reg[8][23]  ( .D(n3788), .CK(n4272), .RN(n3728), .Q(
        \registers[8][23] ) );
  DFFR_X1 \registers_reg[8][22]  ( .D(n3787), .CK(n4272), .RN(n3727), .Q(
        \registers[8][22] ) );
  DFFR_X1 \registers_reg[8][21]  ( .D(n3786), .CK(n4272), .RN(n3727), .Q(
        \registers[8][21] ) );
  DFFR_X1 \registers_reg[8][20]  ( .D(n3785), .CK(n4272), .RN(n3727), .Q(
        \registers[8][20] ) );
  DFFR_X1 \registers_reg[8][19]  ( .D(n3784), .CK(n4272), .RN(n3727), .Q(
        \registers[8][19] ) );
  DFFR_X1 \registers_reg[8][17]  ( .D(n3783), .CK(n4272), .RN(n3727), .Q(
        \registers[8][17] ) );
  DFFR_X1 \registers_reg[8][16]  ( .D(n3782), .CK(n4272), .RN(n3727), .Q(
        \registers[8][16] ) );
  DFFR_X1 \registers_reg[8][15]  ( .D(n3781), .CK(n4272), .RN(n3727), .Q(
        \registers[8][15] ) );
  DFFR_X1 \registers_reg[8][14]  ( .D(n3780), .CK(n4272), .RN(n3727), .Q(
        \registers[8][14] ) );
  DFFR_X1 \registers_reg[8][13]  ( .D(n3779), .CK(n4272), .RN(n3727), .Q(
        \registers[8][13] ) );
  DFFR_X1 \registers_reg[8][12]  ( .D(n3778), .CK(n4272), .RN(n3727), .Q(
        \registers[8][12] ) );
  DFFR_X1 \registers_reg[8][11]  ( .D(n3777), .CK(n4272), .RN(n3726), .Q(
        \registers[8][11] ) );
  DFFR_X1 \registers_reg[8][10]  ( .D(n3776), .CK(n4272), .RN(n3726), .Q(
        \registers[8][10] ) );
  DFFR_X1 \registers_reg[8][9]  ( .D(n3775), .CK(n4272), .RN(n3726), .Q(
        \registers[8][9] ) );
  DFFR_X1 \registers_reg[8][8]  ( .D(n3774), .CK(n4272), .RN(n3726), .Q(
        \registers[8][8] ) );
  DFFR_X1 \registers_reg[8][7]  ( .D(n3773), .CK(n4272), .RN(n3726), .Q(
        \registers[8][7] ) );
  DFFR_X1 \registers_reg[8][6]  ( .D(n3772), .CK(n4272), .RN(n3726), .Q(
        \registers[8][6] ) );
  DFFR_X1 \registers_reg[8][5]  ( .D(n3771), .CK(n4272), .RN(n3726), .Q(
        \registers[8][5] ) );
  DFFR_X1 \registers_reg[8][4]  ( .D(n3770), .CK(n4272), .RN(n3726), .Q(
        \registers[8][4] ) );
  DFFR_X1 \registers_reg[8][3]  ( .D(n3769), .CK(n4272), .RN(n3726), .Q(
        \registers[8][3] ) );
  DFFR_X1 \registers_reg[8][2]  ( .D(n3768), .CK(n4272), .RN(n3726), .Q(
        \registers[8][2] ) );
  DFFR_X1 \registers_reg[8][1]  ( .D(n3767), .CK(n4272), .RN(n3726), .Q(
        \registers[8][1] ) );
  DFFR_X1 \registers_reg[8][0]  ( .D(n3766), .CK(n4272), .RN(n3725), .Q(
        \registers[8][0] ) );
  DFFR_X1 \registers_reg[9][29]  ( .D(n3825), .CK(n4272), .RN(n3725), .Q(
        \registers[9][29] ) );
  DFFR_X1 \registers_reg[9][28]  ( .D(n3824), .CK(n4272), .RN(n3725), .Q(
        \registers[9][28] ) );
  DFFR_X1 \registers_reg[9][26]  ( .D(n3822), .CK(n4272), .RN(n3725), .Q(
        \registers[9][26] ) );
  DFFR_X1 \registers_reg[9][25]  ( .D(n3821), .CK(n4272), .RN(n3725), .Q(
        \registers[9][25] ) );
  DFFR_X1 \registers_reg[9][23]  ( .D(n3819), .CK(n4272), .RN(n3725), .Q(
        \registers[9][23] ) );
  DFFR_X1 \registers_reg[9][22]  ( .D(n3818), .CK(n4272), .RN(n3725), .Q(
        \registers[9][22] ) );
  DFFR_X1 \registers_reg[9][21]  ( .D(n3817), .CK(n4272), .RN(n3724), .Q(
        \registers[9][21] ) );
  DFFR_X1 \registers_reg[9][20]  ( .D(n3816), .CK(n4272), .RN(n3724), .Q(
        \registers[9][20] ) );
  DFFR_X1 \registers_reg[9][18]  ( .D(n3814), .CK(n4272), .RN(n3724), .Q(
        \registers[9][18] ) );
  DFFR_X1 \registers_reg[9][17]  ( .D(n3813), .CK(n4272), .RN(n3724), .Q(
        \registers[9][17] ) );
  DFFR_X1 \registers_reg[9][16]  ( .D(n3812), .CK(n4272), .RN(n3724), .Q(
        \registers[9][16] ) );
  DFFR_X1 \registers_reg[9][13]  ( .D(n3810), .CK(n4272), .RN(n3724), .Q(
        \registers[9][13] ) );
  DFFR_X1 \registers_reg[9][9]  ( .D(n3806), .CK(n4272), .RN(n3723), .Q(
        \registers[9][9] ) );
  DFFR_X1 \registers_reg[9][6]  ( .D(n3803), .CK(n4272), .RN(n3723), .Q(
        \registers[9][6] ) );
  DFFR_X1 \registers_reg[9][5]  ( .D(n3802), .CK(n4272), .RN(n3723), .Q(
        \registers[9][5] ) );
  DFFR_X1 \registers_reg[9][4]  ( .D(n3801), .CK(n4272), .RN(n3723), .Q(
        \registers[9][4] ) );
  DFFR_X1 \registers_reg[9][2]  ( .D(n3799), .CK(n4272), .RN(n3723), .Q(
        \registers[9][2] ) );
  DFFR_X1 \registers_reg[9][1]  ( .D(n3798), .CK(n4272), .RN(n3723), .Q(
        \registers[9][1] ) );
  DFFR_X1 \registers_reg[9][0]  ( .D(n3797), .CK(n4272), .RN(n3723), .Q(
        \registers[9][0] ) );
  DFFR_X1 \registers_reg[10][23]  ( .D(n3149), .CK(n4272), .RN(n3722), .QN(
        n297) );
  DFFR_X1 \registers_reg[11][23]  ( .D(n3117), .CK(n4272), .RN(n3719), .QN(
        n329) );
  DFFR_X1 \registers_reg[11][18]  ( .D(n3112), .CK(n4272), .RN(n3718), .QN(
        n334) );
  DFFR_X1 \registers_reg[11][17]  ( .D(n3111), .CK(n4272), .RN(n3718), .QN(
        n335) );
  DFFR_X1 \registers_reg[11][16]  ( .D(n3110), .CK(n4272), .RN(n3718), .QN(
        n336) );
  DFFR_X1 \registers_reg[11][15]  ( .D(n3109), .CK(n4272), .RN(n3718), .QN(
        n337) );
  DFFR_X1 \registers_reg[11][14]  ( .D(n3108), .CK(n4272), .RN(n3718), .QN(
        n338) );
  DFFR_X1 \registers_reg[11][13]  ( .D(n3107), .CK(n4272), .RN(n3718), .QN(
        n339) );
  DFFR_X1 \registers_reg[11][12]  ( .D(n3106), .CK(n4272), .RN(n3718), .QN(
        n340) );
  DFFR_X1 \registers_reg[11][11]  ( .D(n3105), .CK(n4272), .RN(n3718), .QN(
        n341) );
  DFFR_X1 \registers_reg[11][4]  ( .D(n3098), .CK(n4272), .RN(n3717), .QN(n348) );
  DFFR_X1 \registers_reg[11][3]  ( .D(n3097), .CK(n4272), .RN(n3717), .QN(n349) );
  DFFR_X1 \registers_reg[12][31]  ( .D(n3858), .CK(n4272), .RN(n3717), .Q(
        \registers[12][31] ) );
  DFFR_X1 \registers_reg[12][30]  ( .D(n3857), .CK(n4272), .RN(n3717), .Q(
        \registers[12][30] ) );
  DFFR_X1 \registers_reg[12][29]  ( .D(n3856), .CK(n4272), .RN(n3716), .Q(
        \registers[12][29] ) );
  DFFR_X1 \registers_reg[12][28]  ( .D(n3855), .CK(n4272), .RN(n3716), .Q(
        \registers[12][28] ) );
  DFFR_X1 \registers_reg[12][27]  ( .D(n3854), .CK(n4272), .RN(n3716), .Q(
        \registers[12][27] ) );
  DFFR_X1 \registers_reg[12][26]  ( .D(n3853), .CK(n4272), .RN(n3716), .Q(
        \registers[12][26] ) );
  DFFR_X1 \registers_reg[12][25]  ( .D(n3852), .CK(n4272), .RN(n3716), .Q(
        \registers[12][25] ) );
  DFFR_X1 \registers_reg[12][24]  ( .D(n3851), .CK(n4272), .RN(n3716), .Q(
        \registers[12][24] ) );
  DFFR_X1 \registers_reg[12][23]  ( .D(n3850), .CK(n4272), .RN(n3716), .Q(
        \registers[12][23] ) );
  DFFR_X1 \registers_reg[12][22]  ( .D(n3849), .CK(n4272), .RN(n3716), .Q(
        \registers[12][22] ) );
  DFFR_X1 \registers_reg[12][21]  ( .D(n3848), .CK(n4272), .RN(n3716), .Q(
        \registers[12][21] ) );
  DFFR_X1 \registers_reg[12][20]  ( .D(n3847), .CK(n4272), .RN(n3716), .Q(
        \registers[12][20] ) );
  DFFR_X1 \registers_reg[12][19]  ( .D(n3846), .CK(n4272), .RN(n3716), .Q(
        \registers[12][19] ) );
  DFFR_X1 \registers_reg[12][18]  ( .D(n3845), .CK(n4272), .RN(n3715), .Q(
        \registers[12][18] ) );
  DFFR_X1 \registers_reg[12][17]  ( .D(n3844), .CK(n4272), .RN(n3715), .Q(
        \registers[12][17] ) );
  DFFR_X1 \registers_reg[12][16]  ( .D(n3843), .CK(n4272), .RN(n3715), .Q(
        \registers[12][16] ) );
  DFFR_X1 \registers_reg[12][15]  ( .D(n3842), .CK(n4272), .RN(n3715), .Q(
        \registers[12][15] ) );
  DFFR_X1 \registers_reg[12][14]  ( .D(n3841), .CK(n4272), .RN(n3715), .Q(
        \registers[12][14] ) );
  DFFR_X1 \registers_reg[12][13]  ( .D(n3840), .CK(n4272), .RN(n3715), .Q(
        \registers[12][13] ) );
  DFFR_X1 \registers_reg[12][11]  ( .D(n3839), .CK(n4272), .RN(n3715), .Q(
        \registers[12][11] ) );
  DFFR_X1 \registers_reg[12][10]  ( .D(n3838), .CK(n4272), .RN(n3715), .Q(
        \registers[12][10] ) );
  DFFR_X1 \registers_reg[12][9]  ( .D(n3837), .CK(n4272), .RN(n3715), .Q(
        \registers[12][9] ) );
  DFFR_X1 \registers_reg[12][8]  ( .D(n3836), .CK(n4272), .RN(n3715), .Q(
        \registers[12][8] ) );
  DFFR_X1 \registers_reg[12][7]  ( .D(n3835), .CK(n4272), .RN(n3714), .Q(
        \registers[12][7] ) );
  DFFR_X1 \registers_reg[12][6]  ( .D(n3834), .CK(n4272), .RN(n3714), .Q(
        \registers[12][6] ) );
  DFFR_X1 \registers_reg[12][5]  ( .D(n3833), .CK(n4272), .RN(n3714), .Q(
        \registers[12][5] ) );
  DFFR_X1 \registers_reg[12][4]  ( .D(n3832), .CK(n4272), .RN(n3714), .Q(
        \registers[12][4] ) );
  DFFR_X1 \registers_reg[12][3]  ( .D(n3831), .CK(n4272), .RN(n3714), .Q(
        \registers[12][3] ) );
  DFFR_X1 \registers_reg[12][2]  ( .D(n3830), .CK(n4272), .RN(n3714), .Q(
        \registers[12][2] ) );
  DFFR_X1 \registers_reg[12][1]  ( .D(n3829), .CK(n4272), .RN(n3714), .Q(
        \registers[12][1] ) );
  DFFR_X1 \registers_reg[12][0]  ( .D(n3828), .CK(n4272), .RN(n3714), .Q(
        \registers[12][0] ) );
  DFFR_X1 \registers_reg[13][30]  ( .D(n3888), .CK(n4272), .RN(n3714), .Q(
        \registers[13][30] ) );
  DFFR_X1 \registers_reg[13][29]  ( .D(n3887), .CK(n4272), .RN(n3714), .Q(
        \registers[13][29] ) );
  DFFR_X1 \registers_reg[13][28]  ( .D(n3886), .CK(n4272), .RN(n3713), .Q(
        \registers[13][28] ) );
  DFFR_X1 \registers_reg[13][26]  ( .D(n3884), .CK(n4272), .RN(n3713), .Q(
        \registers[13][26] ) );
  DFFR_X1 \registers_reg[13][25]  ( .D(n3883), .CK(n4272), .RN(n3713), .Q(
        \registers[13][25] ) );
  DFFR_X1 \registers_reg[13][24]  ( .D(n3882), .CK(n4272), .RN(n3713), .Q(
        \registers[13][24] ) );
  DFFR_X1 \registers_reg[13][23]  ( .D(n3881), .CK(n4272), .RN(n3713), .Q(
        \registers[13][23] ) );
  DFFR_X1 \registers_reg[13][22]  ( .D(n3880), .CK(n4272), .RN(n3713), .Q(
        \registers[13][22] ) );
  DFFR_X1 \registers_reg[13][21]  ( .D(n3879), .CK(n4272), .RN(n3713), .Q(
        \registers[13][21] ) );
  DFFR_X1 \registers_reg[13][20]  ( .D(n3878), .CK(n4272), .RN(n3713), .Q(
        \registers[13][20] ) );
  DFFR_X1 \registers_reg[13][18]  ( .D(n3876), .CK(n4272), .RN(n3713), .Q(
        \registers[13][18] ) );
  DFFR_X1 \registers_reg[13][17]  ( .D(n3875), .CK(n4272), .RN(n3712), .Q(
        \registers[13][17] ) );
  DFFR_X1 \registers_reg[13][16]  ( .D(n3874), .CK(n4272), .RN(n3712), .Q(
        \registers[13][16] ) );
  DFFR_X1 \registers_reg[13][13]  ( .D(n3872), .CK(n4272), .RN(n3712), .Q(
        \registers[13][13] ) );
  DFFR_X1 \registers_reg[13][9]  ( .D(n3868), .CK(n4272), .RN(n3712), .Q(
        \registers[13][9] ) );
  DFFR_X1 \registers_reg[13][6]  ( .D(n3865), .CK(n4272), .RN(n3711), .Q(
        \registers[13][6] ) );
  DFFR_X1 \registers_reg[13][5]  ( .D(n3864), .CK(n4272), .RN(n3711), .Q(
        \registers[13][5] ) );
  DFFR_X1 \registers_reg[13][4]  ( .D(n3863), .CK(n4272), .RN(n3711), .Q(
        \registers[13][4] ) );
  DFFR_X1 \registers_reg[13][2]  ( .D(n3861), .CK(n4272), .RN(n3711), .Q(
        \registers[13][2] ) );
  DFFR_X1 \registers_reg[13][1]  ( .D(n3860), .CK(n4272), .RN(n3711), .Q(
        \registers[13][1] ) );
  DFFR_X1 \registers_reg[13][0]  ( .D(n3859), .CK(n4272), .RN(n3711), .Q(
        \registers[13][0] ) );
  DFFR_X1 \registers_reg[15][25]  ( .D(n3055), .CK(n4272), .RN(n3707), .QN(
        n455) );
  DFFR_X1 \registers_reg[15][23]  ( .D(n3053), .CK(n4272), .RN(n3707), .QN(
        n457) );
  DFFR_X1 \registers_reg[15][3]  ( .D(n3033), .CK(n4272), .RN(n3705), .QN(n477) );
  DFFR_X1 \registers_reg[16][23]  ( .D(n3021), .CK(n4272), .RN(n3704), .QN(
        n489) );
  DFFR_X1 \registers_reg[18][31]  ( .D(n4017), .CK(n4272), .RN(n3699), .Q(
        \registers[18][31] ) );
  DFFR_X1 \registers_reg[18][30]  ( .D(n4016), .CK(n4272), .RN(n3699), .Q(
        \registers[18][30] ) );
  DFFR_X1 \registers_reg[18][29]  ( .D(n4015), .CK(n4272), .RN(n3699), .Q(
        \registers[18][29] ) );
  DFFR_X1 \registers_reg[18][28]  ( .D(n4014), .CK(n4272), .RN(n3699), .Q(
        \registers[18][28] ) );
  DFFR_X1 \registers_reg[18][27]  ( .D(n4013), .CK(n4272), .RN(n3699), .Q(
        \registers[18][27] ) );
  DFFR_X1 \registers_reg[18][26]  ( .D(n4012), .CK(n4272), .RN(n3699), .Q(
        \registers[18][26] ) );
  DFFR_X1 \registers_reg[18][25]  ( .D(n4011), .CK(n4272), .RN(n3699), .Q(
        \registers[18][25] ) );
  DFFR_X1 \registers_reg[18][24]  ( .D(n4010), .CK(n4272), .RN(n3699), .Q(
        \registers[18][24] ) );
  DFFR_X1 \registers_reg[18][23]  ( .D(n4009), .CK(n4272), .RN(n3698), .Q(
        \registers[18][23] ) );
  DFFR_X1 \registers_reg[18][22]  ( .D(n4008), .CK(n4272), .RN(n3698), .Q(
        \registers[18][22] ) );
  DFFR_X1 \registers_reg[18][21]  ( .D(n4007), .CK(n4272), .RN(n3698), .Q(
        \registers[18][21] ) );
  DFFR_X1 \registers_reg[18][20]  ( .D(n4006), .CK(n4272), .RN(n3698), .Q(
        \registers[18][20] ) );
  DFFR_X1 \registers_reg[18][19]  ( .D(n4005), .CK(n4272), .RN(n3698), .Q(
        \registers[18][19] ) );
  DFFR_X1 \registers_reg[18][18]  ( .D(n4004), .CK(n4272), .RN(n3698), .Q(
        \registers[18][18] ) );
  DFFR_X1 \registers_reg[18][17]  ( .D(n4003), .CK(n4272), .RN(n3698), .Q(
        \registers[18][17] ) );
  DFFR_X1 \registers_reg[18][16]  ( .D(n4002), .CK(n4272), .RN(n3698), .Q(
        \registers[18][16] ) );
  DFFR_X1 \registers_reg[18][15]  ( .D(n4001), .CK(n4272), .RN(n3698), .Q(
        \registers[18][15] ) );
  DFFR_X1 \registers_reg[18][14]  ( .D(n4000), .CK(n4272), .RN(n3698), .Q(
        \registers[18][14] ) );
  DFFR_X1 \registers_reg[18][13]  ( .D(n3999), .CK(n4272), .RN(n3698), .Q(
        \registers[18][13] ) );
  DFFR_X1 \registers_reg[18][12]  ( .D(n3998), .CK(n4272), .RN(n3697), .Q(
        \registers[18][12] ) );
  DFFR_X1 \registers_reg[18][11]  ( .D(n3997), .CK(n4272), .RN(n3697), .Q(
        \registers[18][11] ) );
  DFFR_X1 \registers_reg[18][10]  ( .D(n3996), .CK(n4272), .RN(n3697), .Q(
        \registers[18][10] ) );
  DFFR_X1 \registers_reg[18][9]  ( .D(n3995), .CK(n4272), .RN(n3697), .Q(
        \registers[18][9] ) );
  DFFR_X1 \registers_reg[18][8]  ( .D(n3994), .CK(n4272), .RN(n3697), .Q(
        \registers[18][8] ) );
  DFFR_X1 \registers_reg[18][7]  ( .D(n3993), .CK(n4272), .RN(n3697), .Q(
        \registers[18][7] ) );
  DFFR_X1 \registers_reg[18][6]  ( .D(n3992), .CK(n4272), .RN(n3697), .Q(
        \registers[18][6] ) );
  DFFR_X1 \registers_reg[18][5]  ( .D(n3991), .CK(n4272), .RN(n3697), .Q(
        \registers[18][5] ) );
  DFFR_X1 \registers_reg[18][4]  ( .D(n3990), .CK(n4272), .RN(n3697), .Q(
        \registers[18][4] ) );
  DFFR_X1 \registers_reg[18][3]  ( .D(n3989), .CK(n4272), .RN(n3697), .Q(
        \registers[18][3] ) );
  DFFR_X1 \registers_reg[18][2]  ( .D(n3988), .CK(n4272), .RN(n3697), .Q(
        \registers[18][2] ) );
  DFFR_X1 \registers_reg[18][1]  ( .D(n3987), .CK(n4272), .RN(n3696), .Q(
        \registers[18][1] ) );
  DFFR_X1 \registers_reg[18][0]  ( .D(n3986), .CK(n4272), .RN(n3696), .Q(
        \registers[18][0] ) );
  DFFR_X1 \registers_reg[19][31]  ( .D(n4049), .CK(n4272), .RN(n3696), .Q(
        \registers[19][31] ) );
  DFFR_X1 \registers_reg[19][30]  ( .D(n4048), .CK(n4272), .RN(n3696), .Q(
        \registers[19][30] ) );
  DFFR_X1 \registers_reg[19][29]  ( .D(n4047), .CK(n4272), .RN(n3696), .Q(
        \registers[19][29] ) );
  DFFR_X1 \registers_reg[19][28]  ( .D(n4046), .CK(n4272), .RN(n3696), .Q(
        \registers[19][28] ) );
  DFFR_X1 \registers_reg[19][27]  ( .D(n4045), .CK(n4272), .RN(n3696), .Q(
        \registers[19][27] ) );
  DFFR_X1 \registers_reg[19][26]  ( .D(n4044), .CK(n4272), .RN(n3696), .Q(
        \registers[19][26] ) );
  DFFR_X1 \registers_reg[19][25]  ( .D(n4043), .CK(n4272), .RN(n3696), .Q(
        \registers[19][25] ) );
  DFFR_X1 \registers_reg[19][23]  ( .D(n4041), .CK(n4272), .RN(n3696), .Q(
        \registers[19][23] ) );
  DFFR_X1 \registers_reg[19][22]  ( .D(n4040), .CK(n4272), .RN(n3695), .Q(
        \registers[19][22] ) );
  DFFR_X1 \registers_reg[19][21]  ( .D(n4039), .CK(n4272), .RN(n3695), .Q(
        \registers[19][21] ) );
  DFFR_X1 \registers_reg[19][20]  ( .D(n4038), .CK(n4272), .RN(n3695), .Q(
        \registers[19][20] ) );
  DFFR_X1 \registers_reg[19][19]  ( .D(n4037), .CK(n4272), .RN(n3695), .Q(
        \registers[19][19] ) );
  DFFR_X1 \registers_reg[19][18]  ( .D(n4036), .CK(n4272), .RN(n3695), .Q(
        \registers[19][18] ) );
  DFFR_X1 \registers_reg[19][17]  ( .D(n4035), .CK(n4272), .RN(n3695), .Q(
        \registers[19][17] ) );
  DFFR_X1 \registers_reg[19][16]  ( .D(n4034), .CK(n4272), .RN(n3695), .Q(
        \registers[19][16] ) );
  DFFR_X1 \registers_reg[19][15]  ( .D(n4033), .CK(n4272), .RN(n3695), .Q(
        \registers[19][15] ) );
  DFFR_X1 \registers_reg[19][14]  ( .D(n4032), .CK(n4272), .RN(n3695), .Q(
        \registers[19][14] ) );
  DFFR_X1 \registers_reg[19][13]  ( .D(n4031), .CK(n4272), .RN(n3695), .Q(
        \registers[19][13] ) );
  DFFR_X1 \registers_reg[19][12]  ( .D(n4030), .CK(n4272), .RN(n3695), .Q(
        \registers[19][12] ) );
  DFFR_X1 \registers_reg[19][11]  ( .D(n4029), .CK(n4272), .RN(n3694), .Q(
        \registers[19][11] ) );
  DFFR_X1 \registers_reg[19][10]  ( .D(n4028), .CK(n4272), .RN(n3694), .Q(
        \registers[19][10] ) );
  DFFR_X1 \registers_reg[19][9]  ( .D(n4027), .CK(n4272), .RN(n3694), .Q(
        \registers[19][9] ) );
  DFFR_X1 \registers_reg[19][8]  ( .D(n4026), .CK(n4272), .RN(n3694), .Q(
        \registers[19][8] ) );
  DFFR_X1 \registers_reg[19][7]  ( .D(n4025), .CK(n4272), .RN(n3694), .Q(
        \registers[19][7] ) );
  DFFR_X1 \registers_reg[19][6]  ( .D(n4024), .CK(n4272), .RN(n3694), .Q(
        \registers[19][6] ) );
  DFFR_X1 \registers_reg[19][5]  ( .D(n4023), .CK(n4272), .RN(n3694), .Q(
        \registers[19][5] ) );
  DFFR_X1 \registers_reg[19][4]  ( .D(n4022), .CK(n4272), .RN(n3694), .Q(
        \registers[19][4] ) );
  DFFR_X1 \registers_reg[19][3]  ( .D(n4021), .CK(n4272), .RN(n3694), .Q(
        \registers[19][3] ) );
  DFFR_X1 \registers_reg[19][2]  ( .D(n4020), .CK(n4272), .RN(n3694), .Q(
        \registers[19][2] ) );
  DFFR_X1 \registers_reg[19][1]  ( .D(n4019), .CK(n4272), .RN(n3694), .Q(
        \registers[19][1] ) );
  DFFR_X1 \registers_reg[19][0]  ( .D(n4018), .CK(n4272), .RN(n3693), .Q(
        \registers[19][0] ) );
  DFFR_X1 \registers_reg[20][23]  ( .D(n2957), .CK(n4272), .RN(n3693), .QN(
        n617) );
  DFFR_X1 \registers_reg[20][22]  ( .D(n2956), .CK(n4272), .RN(n3693), .QN(
        n618) );
  DFFR_X1 \registers_reg[21][23]  ( .D(n2925), .CK(n4272), .RN(n3690), .QN(
        n649) );
  DFFR_X1 \registers_reg[21][22]  ( .D(n2924), .CK(n4272), .RN(n3690), .QN(
        n650) );
  DFFR_X1 \registers_reg[21][12]  ( .D(n2914), .CK(n4272), .RN(n3689), .QN(
        n660) );
  DFFR_X1 \registers_reg[22][7]  ( .D(n4057), .CK(n4272), .RN(n3685), .Q(
        \registers[22][7] ) );
  DFFR_X1 \registers_reg[22][6]  ( .D(n4056), .CK(n4272), .RN(n3685), .Q(
        \registers[22][6] ) );
  DFFR_X1 \registers_reg[22][5]  ( .D(n4055), .CK(n4272), .RN(n3685), .Q(
        \registers[22][5] ) );
  DFFR_X1 \registers_reg[22][4]  ( .D(n4054), .CK(n4272), .RN(n3685), .Q(
        \registers[22][4] ) );
  DFFR_X1 \registers_reg[22][3]  ( .D(n4053), .CK(n4272), .RN(n3685), .Q(
        \registers[22][3] ) );
  DFFR_X1 \registers_reg[22][2]  ( .D(n4052), .CK(n4272), .RN(n3685), .Q(
        \registers[22][2] ) );
  DFFR_X1 \registers_reg[22][1]  ( .D(n4051), .CK(n4272), .RN(n3685), .Q(
        \registers[22][1] ) );
  DFFR_X1 \registers_reg[22][0]  ( .D(n4050), .CK(n4272), .RN(n3685), .Q(
        \registers[22][0] ) );
  DFFR_X1 \registers_reg[23][31]  ( .D(n4108), .CK(n4272), .RN(n3685), .Q(
        \registers[23][31] ) );
  DFFR_X1 \registers_reg[23][30]  ( .D(n4107), .CK(n4272), .RN(n3685), .Q(
        \registers[23][30] ) );
  DFFR_X1 \registers_reg[23][29]  ( .D(n4106), .CK(n4272), .RN(n3684), .Q(
        \registers[23][29] ) );
  DFFR_X1 \registers_reg[23][28]  ( .D(n4105), .CK(n4272), .RN(n3684), .Q(
        \registers[23][28] ) );
  DFFR_X1 \registers_reg[23][27]  ( .D(n4104), .CK(n4272), .RN(n3684), .Q(
        \registers[23][27] ) );
  DFFR_X1 \registers_reg[23][26]  ( .D(n4103), .CK(n4272), .RN(n3684), .Q(
        \registers[23][26] ) );
  DFFR_X1 \registers_reg[23][25]  ( .D(n4102), .CK(n4272), .RN(n3684), .Q(
        \registers[23][25] ) );
  DFFR_X1 \registers_reg[23][23]  ( .D(n4100), .CK(n4272), .RN(n3684), .Q(
        \registers[23][23] ) );
  DFFR_X1 \registers_reg[23][22]  ( .D(n4099), .CK(n4272), .RN(n3684), .Q(
        \registers[23][22] ) );
  DFFR_X1 \registers_reg[23][21]  ( .D(n4098), .CK(n4272), .RN(n3684), .Q(
        \registers[23][21] ) );
  DFFR_X1 \registers_reg[23][20]  ( .D(n4097), .CK(n4272), .RN(n3684), .Q(
        \registers[23][20] ) );
  DFFR_X1 \registers_reg[23][19]  ( .D(n4096), .CK(n4272), .RN(n3684), .Q(
        \registers[23][19] ) );
  DFFR_X1 \registers_reg[23][18]  ( .D(n4095), .CK(n4272), .RN(n3683), .Q(
        \registers[23][18] ) );
  DFFR_X1 \registers_reg[23][17]  ( .D(n4094), .CK(n4272), .RN(n3683), .Q(
        \registers[23][17] ) );
  DFFR_X1 \registers_reg[23][16]  ( .D(n4093), .CK(n4272), .RN(n3683), .Q(
        \registers[23][16] ) );
  DFFR_X1 \registers_reg[23][15]  ( .D(n4092), .CK(n4272), .RN(n3683), .Q(
        \registers[23][15] ) );
  DFFR_X1 \registers_reg[23][14]  ( .D(n4091), .CK(n4272), .RN(n3683), .Q(
        \registers[23][14] ) );
  DFFR_X1 \registers_reg[23][13]  ( .D(n4090), .CK(n4272), .RN(n3683), .Q(
        \registers[23][13] ) );
  DFFR_X1 \registers_reg[23][12]  ( .D(n4089), .CK(n4272), .RN(n3683), .Q(
        \registers[23][12] ) );
  DFFR_X1 \registers_reg[23][11]  ( .D(n4088), .CK(n4272), .RN(n3683), .Q(
        \registers[23][11] ) );
  DFFR_X1 \registers_reg[23][10]  ( .D(n4087), .CK(n4272), .RN(n3683), .Q(
        \registers[23][10] ) );
  DFFR_X1 \registers_reg[23][9]  ( .D(n4086), .CK(n4272), .RN(n3683), .Q(
        \registers[23][9] ) );
  DFFR_X1 \registers_reg[23][8]  ( .D(n4085), .CK(n4272), .RN(n3683), .Q(
        \registers[23][8] ) );
  DFFR_X1 \registers_reg[23][7]  ( .D(n4084), .CK(n4272), .RN(n3682), .Q(
        \registers[23][7] ) );
  DFFR_X1 \registers_reg[23][6]  ( .D(n4083), .CK(n4272), .RN(n3682), .Q(
        \registers[23][6] ) );
  DFFR_X1 \registers_reg[23][5]  ( .D(n4082), .CK(n4272), .RN(n3682), .Q(
        \registers[23][5] ) );
  DFFR_X1 \registers_reg[23][4]  ( .D(n4081), .CK(n4272), .RN(n3682), .Q(
        \registers[23][4] ) );
  DFFR_X1 \registers_reg[23][2]  ( .D(n4080), .CK(n4272), .RN(n3682), .Q(
        \registers[23][2] ) );
  DFFR_X1 \registers_reg[23][1]  ( .D(n4079), .CK(n4272), .RN(n3682), .Q(
        \registers[23][1] ) );
  DFFR_X1 \registers_reg[23][0]  ( .D(n4078), .CK(n4272), .RN(n3682), .Q(
        \registers[23][0] ) );
  DFFR_X1 \registers_reg[24][31]  ( .D(n4138), .CK(n4272), .RN(n3682), .Q(
        \registers[24][31] ) );
  DFFR_X1 \registers_reg[24][30]  ( .D(n4137), .CK(n4272), .RN(n3682), .Q(
        \registers[24][30] ) );
  DFFR_X1 \registers_reg[24][29]  ( .D(n4136), .CK(n4272), .RN(n3682), .Q(
        \registers[24][29] ) );
  DFFR_X1 \registers_reg[24][28]  ( .D(n4135), .CK(n4272), .RN(n3681), .Q(
        \registers[24][28] ) );
  DFFR_X1 \registers_reg[24][27]  ( .D(n4134), .CK(n4272), .RN(n3681), .Q(
        \registers[24][27] ) );
  DFFR_X1 \registers_reg[24][26]  ( .D(n4133), .CK(n4272), .RN(n3681), .Q(
        \registers[24][26] ) );
  DFFR_X1 \registers_reg[24][25]  ( .D(n4132), .CK(n4272), .RN(n3681), .Q(
        \registers[24][25] ) );
  DFFR_X1 \registers_reg[24][24]  ( .D(n226), .CK(n4272), .RN(n3681), .Q(
        \registers[24][24] ), .QN(n227) );
  DFFR_X1 \registers_reg[24][23]  ( .D(n4131), .CK(n4272), .RN(n3681), .Q(
        \registers[24][23] ) );
  DFFR_X1 \registers_reg[24][22]  ( .D(n4130), .CK(n4272), .RN(n3681), .Q(
        \registers[24][22] ) );
  DFFR_X1 \registers_reg[24][20]  ( .D(n4129), .CK(n4272), .RN(n3681), .Q(
        \registers[24][20] ) );
  DFFR_X1 \registers_reg[24][19]  ( .D(n4128), .CK(n4272), .RN(n3681), .Q(
        \registers[24][19] ) );
  DFFR_X1 \registers_reg[24][18]  ( .D(n4127), .CK(n4272), .RN(n3681), .Q(
        \registers[24][18] ) );
  DFFR_X1 \registers_reg[24][17]  ( .D(n4126), .CK(n4272), .RN(n3680), .Q(
        \registers[24][17] ) );
  DFFR_X1 \registers_reg[24][16]  ( .D(n4125), .CK(n4272), .RN(n3680), .Q(
        \registers[24][16] ) );
  DFFR_X1 \registers_reg[24][15]  ( .D(n4124), .CK(n4272), .RN(n3680), .Q(
        \registers[24][15] ) );
  DFFR_X1 \registers_reg[24][14]  ( .D(n4123), .CK(n4272), .RN(n3680), .Q(
        \registers[24][14] ) );
  DFFR_X1 \registers_reg[24][13]  ( .D(n4122), .CK(n4272), .RN(n3680), .Q(
        \registers[24][13] ) );
  DFFR_X1 \registers_reg[24][12]  ( .D(n4121), .CK(n4272), .RN(n3680), .Q(
        \registers[24][12] ) );
  DFFR_X1 \registers_reg[24][11]  ( .D(n4120), .CK(n4272), .RN(n3680), .Q(
        \registers[24][11] ) );
  DFFR_X1 \registers_reg[24][10]  ( .D(n4119), .CK(n4272), .RN(n3680), .Q(
        \registers[24][10] ) );
  DFFR_X1 \registers_reg[24][9]  ( .D(n4118), .CK(n4272), .RN(n3680), .Q(
        \registers[24][9] ) );
  DFFR_X1 \registers_reg[24][8]  ( .D(n4117), .CK(n4272), .RN(n3680), .Q(
        \registers[24][8] ) );
  DFFR_X1 \registers_reg[24][7]  ( .D(n4116), .CK(n4272), .RN(n3680), .Q(
        \registers[24][7] ) );
  DFFR_X1 \registers_reg[24][6]  ( .D(n4115), .CK(n4272), .RN(n3679), .Q(
        \registers[24][6] ) );
  DFFR_X1 \registers_reg[24][5]  ( .D(n4114), .CK(n4272), .RN(n3679), .Q(
        \registers[24][5] ) );
  DFFR_X1 \registers_reg[24][4]  ( .D(n4113), .CK(n4272), .RN(n3679), .Q(
        \registers[24][4] ) );
  DFFR_X1 \registers_reg[24][3]  ( .D(n4112), .CK(n4272), .RN(n3679), .Q(
        \registers[24][3] ) );
  DFFR_X1 \registers_reg[24][2]  ( .D(n4111), .CK(n4272), .RN(n3679), .Q(
        \registers[24][2] ) );
  DFFR_X1 \registers_reg[24][1]  ( .D(n4110), .CK(n4272), .RN(n3679), .Q(
        \registers[24][1] ) );
  DFFR_X1 \registers_reg[24][0]  ( .D(n4109), .CK(n4272), .RN(n3679), .Q(
        \registers[24][0] ) );
  DFFR_X1 \registers_reg[25][31]  ( .D(n4170), .CK(n4272), .RN(n3679), .Q(
        \registers[25][31] ) );
  DFFR_X1 \registers_reg[25][29]  ( .D(n4168), .CK(n4272), .RN(n3679), .Q(
        \registers[25][29] ) );
  DFFR_X1 \registers_reg[25][28]  ( .D(n4167), .CK(n4272), .RN(n3679), .Q(
        \registers[25][28] ) );
  DFFR_X1 \registers_reg[25][27]  ( .D(n4166), .CK(n4272), .RN(n3678), .Q(
        \registers[25][27] ) );
  DFFR_X1 \registers_reg[25][26]  ( .D(n4165), .CK(n4272), .RN(n3678), .Q(
        \registers[25][26] ) );
  DFFR_X1 \registers_reg[25][25]  ( .D(n4164), .CK(n4272), .RN(n3678), .Q(
        \registers[25][25] ) );
  DFFR_X1 \registers_reg[25][24]  ( .D(n4163), .CK(n4272), .RN(n3678), .Q(
        \registers[25][24] ) );
  DFFR_X1 \registers_reg[25][23]  ( .D(n4162), .CK(n4272), .RN(n3678), .Q(
        \registers[25][23] ) );
  DFFR_X1 \registers_reg[25][22]  ( .D(n4161), .CK(n4272), .RN(n3678), .Q(
        \registers[25][22] ) );
  DFFR_X1 \registers_reg[25][21]  ( .D(n4160), .CK(n4272), .RN(n3678), .Q(
        \registers[25][21] ) );
  DFFR_X1 \registers_reg[25][20]  ( .D(n4159), .CK(n4272), .RN(n3678), .Q(
        \registers[25][20] ) );
  DFFR_X1 \registers_reg[25][19]  ( .D(n4158), .CK(n4272), .RN(n3678), .Q(
        \registers[25][19] ) );
  DFFR_X1 \registers_reg[25][18]  ( .D(n4157), .CK(n4272), .RN(n3678), .Q(
        \registers[25][18] ) );
  DFFR_X1 \registers_reg[25][17]  ( .D(n4156), .CK(n4272), .RN(n3678), .Q(
        \registers[25][17] ) );
  DFFR_X1 \registers_reg[25][16]  ( .D(n4155), .CK(n4272), .RN(n3677), .Q(
        \registers[25][16] ) );
  DFFR_X1 \registers_reg[25][15]  ( .D(n4154), .CK(n4272), .RN(n3677), .Q(
        \registers[25][15] ) );
  DFFR_X1 \registers_reg[25][14]  ( .D(n4153), .CK(n4272), .RN(n3677), .Q(
        \registers[25][14] ) );
  DFFR_X1 \registers_reg[25][13]  ( .D(n4152), .CK(n4272), .RN(n3677), .Q(
        \registers[25][13] ) );
  DFFR_X1 \registers_reg[25][12]  ( .D(n4151), .CK(n4272), .RN(n3677), .Q(
        \registers[25][12] ) );
  DFFR_X1 \registers_reg[25][11]  ( .D(n4150), .CK(n4272), .RN(n3677), .Q(
        \registers[25][11] ) );
  DFFR_X1 \registers_reg[25][10]  ( .D(n4149), .CK(n4272), .RN(n3677), .Q(
        \registers[25][10] ) );
  DFFR_X1 \registers_reg[25][9]  ( .D(n4148), .CK(n4272), .RN(n3677), .Q(
        \registers[25][9] ) );
  DFFR_X1 \registers_reg[25][8]  ( .D(n4147), .CK(n4272), .RN(n3677), .Q(
        \registers[25][8] ) );
  DFFR_X1 \registers_reg[25][7]  ( .D(n4146), .CK(n4272), .RN(n3677), .Q(
        \registers[25][7] ) );
  DFFR_X1 \registers_reg[25][6]  ( .D(n4145), .CK(n4272), .RN(n3677), .Q(
        \registers[25][6] ) );
  DFFR_X1 \registers_reg[25][5]  ( .D(n4144), .CK(n4272), .RN(n3676), .Q(
        \registers[25][5] ) );
  DFFR_X1 \registers_reg[25][4]  ( .D(n4143), .CK(n4272), .RN(n3676), .Q(
        \registers[25][4] ) );
  DFFR_X1 \registers_reg[25][3]  ( .D(n4142), .CK(n4272), .RN(n3676), .Q(
        \registers[25][3] ) );
  DFFR_X1 \registers_reg[25][2]  ( .D(n4141), .CK(n4272), .RN(n3676), .Q(
        \registers[25][2] ) );
  DFFR_X1 \registers_reg[25][1]  ( .D(n4140), .CK(n4272), .RN(n3676), .Q(
        \registers[25][1] ) );
  DFFR_X1 \registers_reg[25][0]  ( .D(n4139), .CK(n4272), .RN(n3676), .Q(
        \registers[25][0] ) );
  DFFR_X1 \registers_reg[26][30]  ( .D(n2900), .CK(n4272), .RN(n3676), .QN(
        n802) );
  DFFR_X1 \registers_reg[26][3]  ( .D(n2873), .CK(n4272), .RN(n3673), .QN(n829) );
  DFFR_X1 \registers_reg[27][12]  ( .D(n2850), .CK(n4272), .RN(n3671), .QN(
        n852) );
  DFFR_X1 \registers_reg[28][31]  ( .D(n4201), .CK(n4272), .RN(n3670), .Q(
        \registers[28][31] ) );
  DFFR_X1 \registers_reg[28][29]  ( .D(n4199), .CK(n4272), .RN(n3670), .Q(
        \registers[28][29] ) );
  DFFR_X1 \registers_reg[28][28]  ( .D(n4198), .CK(n4272), .RN(n3670), .Q(
        \registers[28][28] ) );
  DFFR_X1 \registers_reg[28][27]  ( .D(n4197), .CK(n4272), .RN(n3670), .Q(
        \registers[28][27] ) );
  DFFR_X1 \registers_reg[28][26]  ( .D(n4196), .CK(n4272), .RN(n3670), .Q(
        \registers[28][26] ) );
  DFFR_X1 \registers_reg[28][25]  ( .D(n4195), .CK(n4272), .RN(n3670), .Q(
        \registers[28][25] ) );
  DFFR_X1 \registers_reg[28][23]  ( .D(n4193), .CK(n4272), .RN(n3669), .Q(
        \registers[28][23] ) );
  DFFR_X1 \registers_reg[28][22]  ( .D(n4192), .CK(n4272), .RN(n3669), .Q(
        \registers[28][22] ) );
  DFFR_X1 \registers_reg[28][21]  ( .D(n4191), .CK(n4272), .RN(n3669), .Q(
        \registers[28][21] ) );
  DFFR_X1 \registers_reg[28][20]  ( .D(n4190), .CK(n4272), .RN(n3669), .Q(
        \registers[28][20] ) );
  DFFR_X1 \registers_reg[28][19]  ( .D(n4189), .CK(n4272), .RN(n3669), .Q(
        \registers[28][19] ) );
  DFFR_X1 \registers_reg[28][18]  ( .D(n4188), .CK(n4272), .RN(n3669), .Q(
        \registers[28][18] ) );
  DFFR_X1 \registers_reg[28][17]  ( .D(n4187), .CK(n4272), .RN(n3669), .Q(
        \registers[28][17] ) );
  DFFR_X1 \registers_reg[28][16]  ( .D(n4186), .CK(n4272), .RN(n3669), .Q(
        \registers[28][16] ) );
  DFFR_X1 \registers_reg[28][15]  ( .D(n4185), .CK(n4272), .RN(n3669), .Q(
        \registers[28][15] ) );
  DFFR_X1 \registers_reg[28][14]  ( .D(n4184), .CK(n4272), .RN(n3669), .Q(
        \registers[28][14] ) );
  DFFR_X1 \registers_reg[28][13]  ( .D(n4183), .CK(n4272), .RN(n3668), .Q(
        \registers[28][13] ) );
  DFFR_X1 \registers_reg[28][12]  ( .D(n4182), .CK(n4272), .RN(n3668), .Q(
        \registers[28][12] ) );
  DFFR_X1 \registers_reg[28][11]  ( .D(n4181), .CK(n4272), .RN(n3668), .Q(
        \registers[28][11] ) );
  DFFR_X1 \registers_reg[28][10]  ( .D(n4180), .CK(n4272), .RN(n3668), .Q(
        \registers[28][10] ) );
  DFFR_X1 \registers_reg[28][9]  ( .D(n4179), .CK(n4272), .RN(n3668), .Q(
        \registers[28][9] ) );
  DFFR_X1 \registers_reg[28][8]  ( .D(n4178), .CK(n4272), .RN(n3668), .Q(
        \registers[28][8] ) );
  DFFR_X1 \registers_reg[28][7]  ( .D(n236), .CK(n4272), .RN(n3668), .Q(
        \registers[28][7] ), .QN(n237) );
  DFFR_X1 \registers_reg[28][6]  ( .D(n4177), .CK(n4272), .RN(n3668), .Q(
        \registers[28][6] ) );
  DFFR_X1 \registers_reg[28][5]  ( .D(n4176), .CK(n4272), .RN(n3668), .Q(
        \registers[28][5] ) );
  DFFR_X1 \registers_reg[28][4]  ( .D(n4175), .CK(n4272), .RN(n3668), .Q(
        \registers[28][4] ) );
  DFFR_X1 \registers_reg[28][3]  ( .D(n4174), .CK(n4272), .RN(n3668), .Q(
        \registers[28][3] ) );
  DFFR_X1 \registers_reg[28][2]  ( .D(n4173), .CK(n4272), .RN(n3667), .Q(
        \registers[28][2] ) );
  DFFR_X1 \registers_reg[28][1]  ( .D(n4172), .CK(n4272), .RN(n3667), .Q(
        \registers[28][1] ) );
  DFFR_X1 \registers_reg[28][0]  ( .D(n4171), .CK(n4272), .RN(n3667), .Q(
        \registers[28][0] ) );
  DFFR_X1 \registers_reg[29][31]  ( .D(n4232), .CK(n4272), .RN(n3667), .Q(
        \registers[29][31] ) );
  DFFR_X1 \registers_reg[29][30]  ( .D(n4231), .CK(n4272), .RN(n3667), .Q(
        \registers[29][30] ) );
  DFFR_X1 \registers_reg[29][29]  ( .D(n4230), .CK(n4272), .RN(n3667), .Q(
        \registers[29][29] ) );
  DFFR_X1 \registers_reg[29][28]  ( .D(n4229), .CK(n4272), .RN(n3667), .Q(
        \registers[29][28] ) );
  DFFR_X1 \registers_reg[29][27]  ( .D(n4228), .CK(n4272), .RN(n3667), .Q(
        \registers[29][27] ) );
  DFFR_X1 \registers_reg[29][26]  ( .D(n4227), .CK(n4272), .RN(n3667), .Q(
        \registers[29][26] ) );
  DFFR_X1 \registers_reg[29][25]  ( .D(n4226), .CK(n4272), .RN(n3667), .Q(
        \registers[29][25] ) );
  DFFR_X1 \registers_reg[29][23]  ( .D(n4225), .CK(n4272), .RN(n3666), .Q(
        \registers[29][23] ) );
  DFFR_X1 \registers_reg[29][22]  ( .D(n4224), .CK(n4272), .RN(n3666), .Q(
        \registers[29][22] ) );
  DFFR_X1 \registers_reg[29][21]  ( .D(n4223), .CK(n4272), .RN(n3666), .Q(
        \registers[29][21] ) );
  DFFR_X1 \registers_reg[29][20]  ( .D(n4222), .CK(n4272), .RN(n3666), .Q(
        \registers[29][20] ) );
  DFFR_X1 \registers_reg[29][19]  ( .D(n4221), .CK(n4272), .RN(n3666), .Q(
        \registers[29][19] ) );
  DFFR_X1 \registers_reg[29][18]  ( .D(n4220), .CK(n4272), .RN(n3666), .Q(
        \registers[29][18] ) );
  DFFR_X1 \registers_reg[29][17]  ( .D(n4219), .CK(n4272), .RN(n3666), .Q(
        \registers[29][17] ) );
  DFFR_X1 \registers_reg[29][16]  ( .D(n4218), .CK(n4272), .RN(n3666), .Q(
        \registers[29][16] ) );
  DFFR_X1 \registers_reg[29][15]  ( .D(n4217), .CK(n4272), .RN(n3666), .Q(
        \registers[29][15] ) );
  DFFR_X1 \registers_reg[29][14]  ( .D(n4216), .CK(n4272), .RN(n3666), .Q(
        \registers[29][14] ) );
  DFFR_X1 \registers_reg[29][13]  ( .D(n4215), .CK(n4272), .RN(n3666), .Q(
        \registers[29][13] ) );
  DFFR_X1 \registers_reg[29][12]  ( .D(n4214), .CK(n4272), .RN(n3665), .Q(
        \registers[29][12] ) );
  DFFR_X1 \registers_reg[29][11]  ( .D(n4213), .CK(n4272), .RN(n3665), .Q(
        \registers[29][11] ) );
  DFFR_X1 \registers_reg[29][10]  ( .D(n4212), .CK(n4272), .RN(n3665), .Q(
        \registers[29][10] ) );
  DFFR_X1 \registers_reg[29][9]  ( .D(n4211), .CK(n4272), .RN(n3665), .Q(
        \registers[29][9] ) );
  DFFR_X1 \registers_reg[29][8]  ( .D(n4210), .CK(n4272), .RN(n3665), .Q(
        \registers[29][8] ) );
  DFFR_X1 \registers_reg[29][7]  ( .D(n4209), .CK(n4272), .RN(n3665), .Q(
        \registers[29][7] ) );
  DFFR_X1 \registers_reg[29][6]  ( .D(n4208), .CK(n4272), .RN(n3665), .Q(
        \registers[29][6] ) );
  DFFR_X1 \registers_reg[29][5]  ( .D(n4207), .CK(n4272), .RN(n3665), .Q(
        \registers[29][5] ) );
  DFFR_X1 \registers_reg[29][4]  ( .D(n4206), .CK(n4272), .RN(n3665), .Q(
        \registers[29][4] ) );
  DFFR_X1 \registers_reg[29][3]  ( .D(n4205), .CK(n4272), .RN(n3665), .Q(
        \registers[29][3] ) );
  DFFR_X1 \registers_reg[29][2]  ( .D(n4204), .CK(n4272), .RN(n3665), .Q(
        \registers[29][2] ) );
  DFFR_X1 \registers_reg[29][1]  ( .D(n4203), .CK(n4272), .RN(n3664), .Q(
        \registers[29][1] ) );
  DFFR_X1 \registers_reg[29][0]  ( .D(n4202), .CK(n4272), .RN(n3664), .Q(
        \registers[29][0] ) );
  DFFR_X1 \registers_reg[30][19]  ( .D(n2825), .CK(n4272), .RN(n3663), .QN(
        n941) );
  DFFR_X1 \registers_reg[30][12]  ( .D(n2818), .CK(n4272), .RN(n3663), .QN(
        n948) );
  DFFR_X1 \registers_reg[31][24]  ( .D(n2798), .CK(n4272), .RN(n3661), .QN(
        n968) );
  DFFR_X1 \registers_reg[31][4]  ( .D(n2778), .CK(n4272), .RN(n3659), .QN(n988) );
  DLH_X1 \OUT1_reg[31]  ( .G(n3644), .D(N217), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n3644), .D(N216), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n3644), .D(N215), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n3644), .D(N214), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n3644), .D(N213), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n3644), .D(N212), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n3644), .D(N211), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n3644), .D(N210), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n3644), .D(N209), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n3644), .D(N208), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n3645), .D(N207), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n3645), .D(N206), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n3645), .D(N205), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n3645), .D(N204), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n3645), .D(N203), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n3645), .D(N202), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n3645), .D(N201), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n3645), .D(N200), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n3645), .D(N199), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n3645), .D(N198), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n3646), .D(N197), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n3646), .D(N196), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n3646), .D(N195), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n3646), .D(N194), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n3646), .D(N193), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n3646), .D(N192), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n3646), .D(N191), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n3646), .D(N190), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n3646), .D(N189), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n3646), .D(N188), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n3647), .D(N187), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n3647), .D(N186), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(n3640), .D(N352), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n3640), .D(N351), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n3640), .D(N350), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n3640), .D(N349), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n3640), .D(N348), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n3640), .D(N347), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n3640), .D(N346), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n3640), .D(N345), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n3640), .D(N344), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n3640), .D(N343), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n3641), .D(N342), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n3641), .D(N341), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n3641), .D(N340), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n3641), .D(N339), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n3641), .D(N338), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n3641), .D(N337), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n3641), .D(N336), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n3641), .D(N335), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n3641), .D(N334), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n3641), .D(N333), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n3642), .D(N332), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n3642), .D(N331), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n3642), .D(N330), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n3642), .D(N329), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n3642), .D(N328), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n3642), .D(N327), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n3642), .D(N326), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n3642), .D(N325), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n3642), .D(N324), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n3642), .D(N323), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n3643), .D(N322), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n3643), .D(N321), .Q(OUT2[0]) );
  AND3_X2 U531 ( .A1(n1213), .A2(n4233), .A3(ADD_WR[4]), .ZN(n1247) );
  AND3_X2 U796 ( .A1(n3985), .A2(n1213), .A3(ADD_WR[3]), .ZN(n1352) );
  NOR3_X2 U864 ( .A1(n393), .A2(n681), .A3(n4234), .ZN(n1072) );
  NOR3_X2 U966 ( .A1(ADD_WR[2]), .A2(n4236), .A3(n4235), .ZN(n1142) );
  NOR3_X2 U1000 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(n4235), .ZN(n1144) );
  AND3_X2 U1036 ( .A1(n4233), .A2(n3985), .A3(n1213), .ZN(n1521) );
  AND2_X2 U1037 ( .A1(WR), .A2(ENABLE), .ZN(n1213) );
  DFFR_X2 \registers_reg[22][8]  ( .D(n4058), .CK(n4272), .RN(n3685), .Q(
        \registers[22][8] ) );
  DFFR_X2 \registers_reg[22][9]  ( .D(n4059), .CK(n4272), .RN(n3686), .Q(
        \registers[22][9] ) );
  DFFR_X2 \registers_reg[22][10]  ( .D(n4060), .CK(n4272), .RN(n3686), .Q(
        \registers[22][10] ) );
  DFFR_X2 \registers_reg[22][11]  ( .D(n4061), .CK(n4272), .RN(n3686), .Q(
        \registers[22][11] ) );
  DFFR_X2 \registers_reg[22][13]  ( .D(n4062), .CK(n4272), .RN(n3686), .Q(
        \registers[22][13] ) );
  DFFR_X2 \registers_reg[22][14]  ( .D(n4063), .CK(n4272), .RN(n3686), .Q(
        \registers[22][14] ) );
  DFFR_X2 \registers_reg[22][15]  ( .D(n4064), .CK(n4272), .RN(n3686), .Q(
        \registers[22][15] ) );
  DFFR_X2 \registers_reg[22][16]  ( .D(n4065), .CK(n4272), .RN(n3686), .Q(
        \registers[22][16] ) );
  DFFR_X2 \registers_reg[22][17]  ( .D(n4066), .CK(n4272), .RN(n3686), .Q(
        \registers[22][17] ) );
  DFFR_X2 \registers_reg[22][18]  ( .D(n4067), .CK(n4272), .RN(n3686), .Q(
        \registers[22][18] ) );
  DFFR_X2 \registers_reg[22][19]  ( .D(n4068), .CK(n4272), .RN(n3686), .Q(
        \registers[22][19] ) );
  DFFR_X2 \registers_reg[22][21]  ( .D(n4069), .CK(n4272), .RN(n3687), .Q(
        \registers[22][21] ) );
  DFFR_X2 \registers_reg[22][23]  ( .D(n4070), .CK(n4272), .RN(n3687), .Q(
        \registers[22][23] ) );
  DFFR_X2 \registers_reg[22][24]  ( .D(n4071), .CK(n4272), .RN(n3687), .Q(
        \registers[22][24] ) );
  DFFR_X2 \registers_reg[22][25]  ( .D(n4072), .CK(n4272), .RN(n3687), .Q(
        \registers[22][25] ) );
  DFFR_X2 \registers_reg[22][26]  ( .D(n4073), .CK(n4272), .RN(n3687), .Q(
        \registers[22][26] ) );
  DFFR_X2 \registers_reg[22][27]  ( .D(n4074), .CK(n4272), .RN(n3687), .Q(
        \registers[22][27] ) );
  DFFR_X2 \registers_reg[22][29]  ( .D(n4075), .CK(n4272), .RN(n3687), .Q(
        \registers[22][29] ) );
  DFFR_X2 \registers_reg[22][30]  ( .D(n4076), .CK(n4272), .RN(n3687), .Q(
        \registers[22][30] ) );
  DFFR_X2 \registers_reg[22][31]  ( .D(n4077), .CK(n4272), .RN(n3688), .Q(
        \registers[22][31] ) );
  DFFR_X2 \registers_reg[6][8]  ( .D(n3930), .CK(n4272), .RN(n3732), .Q(
        \registers[6][8] ) );
  DFFR_X2 \registers_reg[6][10]  ( .D(n3932), .CK(n4272), .RN(n3732), .Q(
        \registers[6][10] ) );
  DFFR_X2 \registers_reg[6][13]  ( .D(n3935), .CK(n4272), .RN(n3732), .Q(
        \registers[6][13] ) );
  DFFR_X2 \registers_reg[6][16]  ( .D(n3937), .CK(n4272), .RN(n3733), .Q(
        \registers[6][16] ) );
  DFFR_X2 \registers_reg[6][18]  ( .D(n3939), .CK(n4272), .RN(n3733), .Q(
        \registers[6][18] ) );
  DFFR_X2 \registers_reg[6][21]  ( .D(n3942), .CK(n4272), .RN(n3733), .Q(
        \registers[6][21] ) );
  DFFR_X2 \registers_reg[6][23]  ( .D(n3944), .CK(n4272), .RN(n3733), .Q(
        \registers[6][23] ) );
  DFFR_X2 \registers_reg[6][24]  ( .D(n3945), .CK(n4272), .RN(n3733), .Q(
        \registers[6][24] ) );
  DFFR_X2 \registers_reg[6][25]  ( .D(n3946), .CK(n4272), .RN(n3734), .Q(
        \registers[6][25] ) );
  DFFR_X2 \registers_reg[6][26]  ( .D(n3947), .CK(n4272), .RN(n3734), .Q(
        \registers[6][26] ) );
  DFFR_X2 \registers_reg[6][27]  ( .D(n3948), .CK(n4272), .RN(n3734), .Q(
        \registers[6][27] ) );
  DFFR_X2 \registers_reg[6][29]  ( .D(n3950), .CK(n4272), .RN(n3734), .Q(
        \registers[6][29] ) );
  DFFR_X2 \registers_reg[6][30]  ( .D(n3951), .CK(n4272), .RN(n3734), .Q(
        \registers[6][30] ) );
  DFFR_X2 \registers_reg[9][3]  ( .D(n3800), .CK(n4272), .RN(n3723), .Q(
        \registers[9][3] ) );
  DFFR_X2 \registers_reg[9][7]  ( .D(n3804), .CK(n4272), .RN(n3723), .Q(
        \registers[9][7] ) );
  DFFR_X2 \registers_reg[9][8]  ( .D(n3805), .CK(n4272), .RN(n3723), .Q(
        \registers[9][8] ) );
  DFFR_X2 \registers_reg[9][10]  ( .D(n3807), .CK(n4272), .RN(n3723), .Q(
        \registers[9][10] ) );
  DFFR_X2 \registers_reg[9][11]  ( .D(n3808), .CK(n4272), .RN(n3724), .Q(
        \registers[9][11] ) );
  DFFR_X2 \registers_reg[9][15]  ( .D(n3811), .CK(n4272), .RN(n3724), .Q(
        \registers[9][15] ) );
  DFFR_X2 \registers_reg[9][19]  ( .D(n3815), .CK(n4272), .RN(n3724), .Q(
        \registers[9][19] ) );
  DFFR_X2 \registers_reg[9][27]  ( .D(n3823), .CK(n4272), .RN(n3725), .Q(
        \registers[9][27] ) );
  DFFR_X2 \registers_reg[9][31]  ( .D(n3827), .CK(n4272), .RN(n3725), .Q(
        \registers[9][31] ) );
  DFFR_X2 \registers_reg[1][3]  ( .D(n3893), .CK(n4272), .RN(n3746), .Q(
        \registers[1][3] ) );
  DFFR_X2 \registers_reg[1][8]  ( .D(n3898), .CK(n4272), .RN(n3747), .Q(
        \registers[1][8] ) );
  DFFR_X2 \registers_reg[1][10]  ( .D(n3900), .CK(n4272), .RN(n3747), .Q(
        \registers[1][10] ) );
  DFFR_X2 \registers_reg[1][11]  ( .D(n3901), .CK(n4272), .RN(n3747), .Q(
        \registers[1][11] ) );
  DFFR_X2 \registers_reg[1][12]  ( .D(n3902), .CK(n4272), .RN(n3747), .Q(
        \registers[1][12] ) );
  DFFR_X2 \registers_reg[1][14]  ( .D(n3904), .CK(n4272), .RN(n3747), .Q(
        \registers[1][14] ) );
  DFFR_X2 \registers_reg[1][15]  ( .D(n3905), .CK(n4272), .RN(n3747), .Q(
        \registers[1][15] ) );
  DFFR_X2 \registers_reg[1][19]  ( .D(n3909), .CK(n4272), .RN(n3748), .Q(
        \registers[1][19] ) );
  DFFR_X2 \registers_reg[1][27]  ( .D(n3917), .CK(n4272), .RN(n3748), .Q(
        \registers[1][27] ) );
  DFFR_X2 \registers_reg[1][31]  ( .D(n3921), .CK(n4272), .RN(n3749), .Q(
        \registers[1][31] ) );
  DFFR_X2 \registers_reg[13][10]  ( .D(n3869), .CK(n4272), .RN(n3712), .Q(
        \registers[13][10] ) );
  DFFR_X2 \registers_reg[13][11]  ( .D(n3870), .CK(n4272), .RN(n3712), .Q(
        \registers[13][11] ) );
  DFFR_X2 \registers_reg[13][14]  ( .D(n3873), .CK(n4272), .RN(n3712), .Q(
        \registers[13][14] ) );
  DFFR_X2 \registers_reg[13][19]  ( .D(n3877), .CK(n4272), .RN(n3713), .Q(
        \registers[13][19] ) );
  DFFR_X2 \registers_reg[13][31]  ( .D(n3889), .CK(n4272), .RN(n3714), .Q(
        \registers[13][31] ) );
  DFFR_X2 \registers_reg[13][3]  ( .D(n3862), .CK(n4272), .RN(n3711), .Q(
        \registers[13][3] ) );
  DFFR_X2 \registers_reg[13][8]  ( .D(n3867), .CK(n4272), .RN(n3712), .Q(
        \registers[13][8] ) );
  DFFR_X2 \registers_reg[13][27]  ( .D(n3885), .CK(n4272), .RN(n3713), .Q(
        \registers[13][27] ) );
  DFFR_X1 \registers_reg[22][28]  ( .D(net18066), .CK(n4272), .RN(n3687), .Q(
        \registers[22][28] ) );
  DFFR_X1 \registers_reg[6][14]  ( .D(n3936), .CK(n4272), .RN(n3733), .Q(
        \registers[6][14] ) );
  DFFR_X1 \registers_reg[6][28]  ( .D(n3949), .CK(n4272), .RN(n3734), .Q(
        \registers[6][28] ) );
  DFFR_X1 \registers_reg[6][12]  ( .D(n3934), .CK(n4272), .RN(n3732), .Q(
        \registers[6][12] ) );
  DFFR_X1 \registers_reg[13][7]  ( .D(n3866), .CK(n4272), .RN(n3712), .Q(
        \registers[13][7] ) );
  DFFR_X1 \registers_reg[13][12]  ( .D(n3871), .CK(n4272), .RN(n3712), .Q(
        \registers[13][12] ) );
  DFFR_X1 \registers_reg[9][12]  ( .D(n3809), .CK(n4272), .RN(n3724), .Q(
        \registers[9][12] ) );
  DFFR_X1 \registers_reg[1][7]  ( .D(n3897), .CK(n4272), .RN(n3746), .Q(
        \registers[1][7] ) );
  DFFR_X1 \registers_reg[16][12]  ( .D(n3010), .CK(n4272), .RN(n3703), .QN(
        n500) );
  DFFR_X1 \registers_reg[5][12]  ( .D(n3170), .CK(n4272), .RN(n3735), .QN(n148) );
  DFFR_X1 \registers_reg[26][12]  ( .D(n2882), .CK(n4272), .RN(n3674), .QN(
        n820) );
  DFFR_X1 \registers_reg[14][30]  ( .D(n3092), .CK(n4272), .RN(n3711), .QN(
        n418) );
  DFFR_X1 \registers_reg[3][30]  ( .D(n3252), .CK(n4272), .RN(n3743), .QN(n66)
         );
  DFFR_X1 \registers_reg[2][12]  ( .D(n3266), .CK(n4272), .RN(n3744), .QN(n52)
         );
  DFFR_X1 \registers_reg[14][25]  ( .D(n3087), .CK(n4272), .RN(n3710), .QN(
        n423) );
  DFFR_X1 \registers_reg[14][21]  ( .D(n3083), .CK(n4272), .RN(n3710), .QN(
        n427) );
  DFFR_X1 \registers_reg[15][19]  ( .D(n3049), .CK(n4272), .RN(n3707), .QN(
        n461) );
  DFFR_X1 \registers_reg[20][12]  ( .D(n2946), .CK(n4272), .RN(n3692), .QN(
        n628) );
  DFFR_X1 \registers_reg[3][25]  ( .D(n3247), .CK(n4272), .RN(n3742), .QN(n71)
         );
  DFFR_X1 \registers_reg[2][25]  ( .D(n3279), .CK(n4272), .RN(n3745), .QN(n39)
         );
  DFFR_X1 \registers_reg[15][31]  ( .D(n3061), .CK(n4272), .RN(n3708), .QN(
        n449) );
  DFFR_X1 \registers_reg[17][31]  ( .D(n2997), .CK(n4272), .RN(n3702), .QN(
        n513) );
  DFFR_X1 \registers_reg[26][25]  ( .D(n2895), .CK(n4272), .RN(n3675), .QN(
        n807) );
  DFFR_X1 \registers_reg[26][21]  ( .D(n2891), .CK(n4272), .RN(n3675), .QN(
        n811) );
  DFFR_X1 \registers_reg[14][19]  ( .D(n3081), .CK(n4272), .RN(n3710), .QN(
        n429) );
  DFFR_X1 \registers_reg[30][25]  ( .D(n2831), .CK(n4272), .RN(n3664), .QN(
        n935) );
  DFFR_X1 \registers_reg[11][20]  ( .D(n3114), .CK(n4272), .RN(n3719), .QN(
        n332) );
  DFFR_X1 \registers_reg[2][19]  ( .D(n3273), .CK(n4272), .RN(n3745), .QN(n45)
         );
  DFFR_X1 \registers_reg[30][21]  ( .D(n2827), .CK(n4272), .RN(n3663), .QN(
        n939) );
  DFFR_X1 \registers_reg[2][15]  ( .D(n3269), .CK(n4272), .RN(n3744), .QN(n49)
         );
  DFFR_X1 \registers_reg[21][30]  ( .D(n2932), .CK(n4272), .RN(n3690), .QN(
        n642) );
  DFFR_X1 \registers_reg[5][30]  ( .D(n3188), .CK(n4272), .RN(n3737), .QN(n130) );
  DFFR_X1 \registers_reg[17][30]  ( .D(n2996), .CK(n4272), .RN(n3702), .QN(
        n514) );
  DFFR_X1 \registers_reg[10][29]  ( .D(n3155), .CK(n4272), .RN(n3722), .QN(
        n291) );
  DFFR_X1 \registers_reg[17][29]  ( .D(n2995), .CK(n4272), .RN(n3702), .QN(
        n515) );
  DFFR_X1 \registers_reg[15][29]  ( .D(n3059), .CK(n4272), .RN(n3708), .QN(
        n451) );
  DFFR_X1 \registers_reg[21][15]  ( .D(n2917), .CK(n4272), .RN(n3689), .QN(
        n657) );
  DFFR_X1 \registers_reg[30][14]  ( .D(n2820), .CK(n4272), .RN(n3663), .QN(
        n946) );
  DFFR_X1 \registers_reg[5][19]  ( .D(n3177), .CK(n4272), .RN(n3736), .QN(n141) );
  DFFR_X1 \registers_reg[14][29]  ( .D(n3091), .CK(n4272), .RN(n3711), .QN(
        n419) );
  DFFR_X1 \registers_reg[21][31]  ( .D(n2933), .CK(n4272), .RN(n3690), .QN(
        n641) );
  DFFR_X1 \registers_reg[30][13]  ( .D(n2819), .CK(n4272), .RN(n3663), .QN(
        n947) );
  DFFR_X1 \registers_reg[30][9]  ( .D(n2815), .CK(n4272), .RN(n3662), .QN(n951) );
  DFFR_X1 \registers_reg[30][6]  ( .D(n2812), .CK(n4272), .RN(n3662), .QN(n954) );
  DFFR_X1 \registers_reg[26][19]  ( .D(n2889), .CK(n4272), .RN(n3675), .QN(
        n813) );
  DFFR_X1 \registers_reg[10][30]  ( .D(n3156), .CK(n4272), .RN(n3722), .QN(
        n290) );
  DFFR_X1 \registers_reg[30][18]  ( .D(n2824), .CK(n4272), .RN(n3663), .QN(
        n942) );
  DFFR_X1 \registers_reg[14][13]  ( .D(n3075), .CK(n4272), .RN(n3709), .QN(
        n435) );
  DFFR_X1 \registers_reg[14][10]  ( .D(n3072), .CK(n4272), .RN(n3709), .QN(
        n438) );
  DFFR_X1 \registers_reg[14][9]  ( .D(n3071), .CK(n4272), .RN(n3709), .QN(n439) );
  DFFR_X1 \registers_reg[14][6]  ( .D(n3068), .CK(n4272), .RN(n3709), .QN(n442) );
  DFFR_X1 \registers_reg[21][25]  ( .D(n2927), .CK(n4272), .RN(n3690), .QN(
        n647) );
  DFFR_X1 \registers_reg[21][19]  ( .D(n2921), .CK(n4272), .RN(n3689), .QN(
        n653) );
  DFFR_X1 \registers_reg[31][25]  ( .D(n2799), .CK(n4272), .RN(n3661), .QN(
        n967) );
  DFFR_X1 \registers_reg[14][20]  ( .D(n3082), .CK(n4272), .RN(n3710), .QN(
        n428) );
  DFFR_X1 \registers_reg[26][15]  ( .D(n2885), .CK(n4272), .RN(n3674), .QN(
        n817) );
  DFFR_X1 \registers_reg[21][28]  ( .D(n2930), .CK(n4272), .RN(n3690), .QN(
        n644) );
  DFFR_X1 \registers_reg[5][28]  ( .D(n3186), .CK(n4272), .RN(n3737), .QN(n132) );
  DFFR_X1 \registers_reg[5][14]  ( .D(n3172), .CK(n4272), .RN(n3735), .QN(n146) );
  DFFR_X1 \registers_reg[21][14]  ( .D(n2916), .CK(n4272), .RN(n3689), .QN(
        n658) );
  DFFR_X1 \registers_reg[15][10]  ( .D(n3040), .CK(n4272), .RN(n3706), .QN(
        n470) );
  DFFR_X1 \registers_reg[15][28]  ( .D(n3058), .CK(n4272), .RN(n3708), .QN(
        n452) );
  DFFR_X1 \registers_reg[15][1]  ( .D(n3031), .CK(n4272), .RN(n3705), .QN(n479) );
  DFFR_X1 \registers_reg[3][6]  ( .D(n3228), .CK(n4272), .RN(n3741), .QN(n90)
         );
  DFFR_X1 \registers_reg[3][1]  ( .D(n3223), .CK(n4272), .RN(n3740), .QN(n95)
         );
  DFFR_X1 \registers_reg[2][1]  ( .D(n3255), .CK(n4272), .RN(n3743), .QN(n63)
         );
  DFFR_X1 \registers_reg[3][13]  ( .D(n3235), .CK(n4272), .RN(n3741), .QN(n83)
         );
  DFFR_X1 \registers_reg[3][10]  ( .D(n3232), .CK(n4272), .RN(n3741), .QN(n86)
         );
  DFFR_X1 \registers_reg[3][9]  ( .D(n3231), .CK(n4272), .RN(n3741), .QN(n87)
         );
  DFFR_X1 \registers_reg[2][13]  ( .D(n3267), .CK(n4272), .RN(n3744), .QN(n51)
         );
  DFFR_X1 \registers_reg[2][10]  ( .D(n3264), .CK(n4272), .RN(n3744), .QN(n54)
         );
  DFFR_X1 \registers_reg[20][9]  ( .D(n2943), .CK(n4272), .RN(n3691), .QN(n631) );
  DFFR_X1 \registers_reg[4][18]  ( .D(n3208), .CK(n4272), .RN(n3739), .QN(n110) );
  DFFR_X1 \registers_reg[4][13]  ( .D(n3203), .CK(n4272), .RN(n3738), .QN(n115) );
  DFFR_X1 \registers_reg[21][13]  ( .D(n2915), .CK(n4272), .RN(n3689), .QN(
        n659) );
  DFFR_X1 \registers_reg[21][6]  ( .D(n2908), .CK(n4272), .RN(n3688), .QN(n666) );
  DFFR_X1 \registers_reg[5][18]  ( .D(n3176), .CK(n4272), .RN(n3736), .QN(n142) );
  DFFR_X1 \registers_reg[5][10]  ( .D(n3168), .CK(n4272), .RN(n3735), .QN(n150) );
  DFFR_X1 \registers_reg[5][9]  ( .D(n3167), .CK(n4272), .RN(n3735), .QN(n151)
         );
  DFFR_X1 \registers_reg[5][1]  ( .D(n3159), .CK(n4272), .RN(n3734), .QN(n159)
         );
  DFFR_X1 \registers_reg[16][10]  ( .D(n3008), .CK(n4272), .RN(n3703), .QN(
        n502) );
  DFFR_X1 \registers_reg[16][9]  ( .D(n3007), .CK(n4272), .RN(n3703), .QN(n503) );
  DFFR_X1 \registers_reg[17][1]  ( .D(n2967), .CK(n4272), .RN(n3699), .QN(n543) );
  DFFR_X1 \registers_reg[16][13]  ( .D(n3011), .CK(n4272), .RN(n3703), .QN(
        n499) );
  DFFR_X1 \registers_reg[26][13]  ( .D(n2883), .CK(n4272), .RN(n3674), .QN(
        n819) );
  DFFR_X1 \registers_reg[26][10]  ( .D(n2880), .CK(n4272), .RN(n3674), .QN(
        n822) );
  DFFR_X1 \registers_reg[26][9]  ( .D(n2879), .CK(n4272), .RN(n3674), .QN(n823) );
  DFFR_X1 \registers_reg[26][6]  ( .D(n2876), .CK(n4272), .RN(n3674), .QN(n826) );
  DFFR_X1 \registers_reg[14][1]  ( .D(n3063), .CK(n4272), .RN(n3708), .QN(n447) );
  DFFR_X1 \registers_reg[14][28]  ( .D(n3090), .CK(n4272), .RN(n3711), .QN(
        n420) );
  DFFR_X1 \registers_reg[3][20]  ( .D(n3242), .CK(n4272), .RN(n3742), .QN(n76)
         );
  DFFR_X1 \registers_reg[2][20]  ( .D(n3274), .CK(n4272), .RN(n3745), .QN(n44)
         );
  DFFR_X1 \registers_reg[26][1]  ( .D(n2871), .CK(n4272), .RN(n3673), .QN(n831) );
  DFFR_X1 \registers_reg[30][11]  ( .D(n2817), .CK(n4272), .RN(n3662), .QN(
        n949) );
  DFFR_X1 \registers_reg[5][11]  ( .D(n3169), .CK(n4272), .RN(n3735), .QN(n149) );
  DFFR_X1 \registers_reg[15][12]  ( .D(n3042), .CK(n4272), .RN(n3706), .QN(
        n468) );
  DFFR_X1 \registers_reg[10][12]  ( .D(n3138), .CK(n4272), .RN(n3721), .QN(
        n308) );
  DFFR_X1 \registers_reg[27][29]  ( .D(n2867), .CK(n4272), .RN(n3673), .QN(
        n835) );
  DFFR_X1 \registers_reg[27][28]  ( .D(n2866), .CK(n4272), .RN(n3673), .QN(
        n836) );
  DFFR_X1 \registers_reg[27][25]  ( .D(n2863), .CK(n4272), .RN(n3672), .QN(
        n839) );
  DFFR_X1 \registers_reg[27][21]  ( .D(n2859), .CK(n4272), .RN(n3672), .QN(
        n843) );
  DFFR_X1 \registers_reg[27][20]  ( .D(n2858), .CK(n4272), .RN(n3672), .QN(
        n844) );
  DFFR_X1 \registers_reg[27][19]  ( .D(n2857), .CK(n4272), .RN(n3672), .QN(
        n845) );
  DFFR_X1 \registers_reg[27][10]  ( .D(n2848), .CK(n4272), .RN(n3671), .QN(
        n854) );
  DFFR_X1 \registers_reg[27][1]  ( .D(n2839), .CK(n4272), .RN(n3670), .QN(n863) );
  DFFR_X1 \registers_reg[17][19]  ( .D(n2985), .CK(n4272), .RN(n3701), .QN(
        n525) );
  DFFR_X1 \registers_reg[10][7]  ( .D(n3133), .CK(n4272), .RN(n3720), .QN(n313) );
  DFFR_X1 \registers_reg[3][24]  ( .D(n3246), .CK(n4272), .RN(n3742), .QN(n72)
         );
  DFFR_X1 \registers_reg[3][29]  ( .D(n3251), .CK(n4272), .RN(n3743), .QN(n67)
         );
  DFFR_X1 \registers_reg[11][29]  ( .D(n3123), .CK(n4272), .RN(n3719), .QN(
        n323) );
  DFFR_X1 \registers_reg[2][29]  ( .D(n3283), .CK(n4272), .RN(n3746), .QN(n35)
         );
  DFFR_X1 \registers_reg[17][12]  ( .D(n2978), .CK(n4272), .RN(n3700), .QN(
        n532) );
  DFFR_X1 \registers_reg[17][14]  ( .D(n2980), .CK(n4272), .RN(n3701), .QN(
        n530) );
  DFFR_X1 \registers_reg[27][22]  ( .D(n2860), .CK(n4272), .RN(n3672), .QN(
        n842) );
  DFFR_X1 \registers_reg[27][7]  ( .D(n2845), .CK(n4272), .RN(n3671), .QN(n857) );
  DFFR_X1 \registers_reg[30][20]  ( .D(n2826), .CK(n4272), .RN(n3663), .QN(
        n940) );
  DFFR_X1 \registers_reg[21][20]  ( .D(n2922), .CK(n4272), .RN(n3689), .QN(
        n652) );
  DFFR_X1 \registers_reg[5][20]  ( .D(n3178), .CK(n4272), .RN(n3736), .QN(n140) );
  DFFR_X1 \registers_reg[11][9]  ( .D(n3103), .CK(n4272), .RN(n3718), .QN(n343) );
  DFFR_X1 \registers_reg[11][28]  ( .D(n3122), .CK(n4272), .RN(n3719), .QN(
        n324) );
  DFFR_X1 \registers_reg[10][2]  ( .D(n3128), .CK(n4272), .RN(n3720), .QN(n318) );
  DFFR_X1 \registers_reg[17][2]  ( .D(n2968), .CK(n4272), .RN(n3699), .QN(n542) );
  DFFR_X1 \registers_reg[15][30]  ( .D(n3060), .CK(n4272), .RN(n3708), .QN(
        n450) );
  DFFR_X1 \registers_reg[17][3]  ( .D(n2969), .CK(n4272), .RN(n3700), .QN(n541) );
  DFFR_X1 \registers_reg[15][2]  ( .D(n3032), .CK(n4272), .RN(n3705), .QN(n478) );
  DFFR_X1 \registers_reg[26][20]  ( .D(n2890), .CK(n4272), .RN(n3675), .QN(
        n812) );
  DFFR_X1 \registers_reg[15][8]  ( .D(n3038), .CK(n4272), .RN(n3706), .QN(n472) );
  DFFR_X1 \registers_reg[14][8]  ( .D(n3070), .CK(n4272), .RN(n3709), .QN(n440) );
  DFFR_X1 \registers_reg[10][8]  ( .D(n3134), .CK(n4272), .RN(n3720), .QN(n312) );
  DFFR_X1 \registers_reg[10][5]  ( .D(n3131), .CK(n4272), .RN(n3720), .QN(n315) );
  DFFR_X1 \registers_reg[5][29]  ( .D(n3187), .CK(n4272), .RN(n3737), .QN(n131) );
  DFFR_X1 \registers_reg[11][30]  ( .D(n3124), .CK(n4272), .RN(n3719), .QN(
        n322) );
  DFFR_X1 \registers_reg[14][31]  ( .D(n3093), .CK(n4272), .RN(n3711), .QN(
        n417) );
  DFFR_X1 \registers_reg[14][22]  ( .D(n3084), .CK(n4272), .RN(n3710), .QN(
        n426) );
  DFFR_X1 \registers_reg[14][7]  ( .D(n3069), .CK(n4272), .RN(n3709), .QN(n441) );
  DFFR_X1 \registers_reg[14][12]  ( .D(n3074), .CK(n4272), .RN(n3709), .QN(
        n436) );
  DFFR_X1 \registers_reg[16][11]  ( .D(n3009), .CK(n4272), .RN(n3703), .QN(
        n501) );
  DFFR_X1 \registers_reg[10][11]  ( .D(n3137), .CK(n4272), .RN(n3721), .QN(
        n309) );
  DFFR_X1 \registers_reg[14][3]  ( .D(n3065), .CK(n4272), .RN(n3708), .QN(n445) );
  DFFR_X1 \registers_reg[16][27]  ( .D(n3025), .CK(n4272), .RN(n3705), .QN(
        n485) );
  DFFR_X1 \registers_reg[16][26]  ( .D(n3024), .CK(n4272), .RN(n3705), .QN(
        n486) );
  DFFR_X1 \registers_reg[10][27]  ( .D(n3153), .CK(n4272), .RN(n3722), .QN(
        n293) );
  DFFR_X1 \registers_reg[10][26]  ( .D(n3152), .CK(n4272), .RN(n3722), .QN(
        n294) );
  DFFR_X1 \registers_reg[21][29]  ( .D(n2931), .CK(n4272), .RN(n3690), .QN(
        n643) );
  DFFR_X1 \registers_reg[17][5]  ( .D(n2971), .CK(n4272), .RN(n3700), .QN(n539) );
  DFFR_X1 \registers_reg[14][27]  ( .D(n3089), .CK(n4272), .RN(n3710), .QN(
        n421) );
  DFFR_X1 \registers_reg[15][11]  ( .D(n3041), .CK(n4272), .RN(n3706), .QN(
        n469) );
  DFFR_X1 \registers_reg[26][29]  ( .D(n2899), .CK(n4272), .RN(n3676), .QN(
        n803) );
  DFFR_X1 \registers_reg[15][27]  ( .D(n3057), .CK(n4272), .RN(n3708), .QN(
        n453) );
  DFFR_X1 \registers_reg[15][26]  ( .D(n3056), .CK(n4272), .RN(n3707), .QN(
        n454) );
  DFFR_X1 \registers_reg[15][5]  ( .D(n3035), .CK(n4272), .RN(n3706), .QN(n475) );
  DFFR_X1 \registers_reg[17][11]  ( .D(n2977), .CK(n4272), .RN(n3700), .QN(
        n533) );
  DFFR_X1 \registers_reg[26][7]  ( .D(n2877), .CK(n4272), .RN(n3674), .QN(n825) );
  DFFR_X1 \registers_reg[10][20]  ( .D(n3146), .CK(n4272), .RN(n3721), .QN(
        n300) );
  DFFR_X1 \registers_reg[10][19]  ( .D(n3145), .CK(n4272), .RN(n3721), .QN(
        n301) );
  DFFR_X1 \registers_reg[10][24]  ( .D(n3150), .CK(n4272), .RN(n3722), .QN(
        n296) );
  DFFR_X1 \registers_reg[11][8]  ( .D(n3102), .CK(n4272), .RN(n3717), .QN(n344) );
  DFFR_X1 \registers_reg[17][8]  ( .D(n2974), .CK(n4272), .RN(n3700), .QN(n536) );
  DFFR_X1 \registers_reg[16][8]  ( .D(n3006), .CK(n4272), .RN(n3703), .QN(n504) );
  DFFR_X1 \registers_reg[10][4]  ( .D(n3130), .CK(n4272), .RN(n3720), .QN(n316) );
  DFFR_X1 \registers_reg[27][2]  ( .D(n2840), .CK(n4272), .RN(n3670), .QN(n862) );
  DFFR_X1 \registers_reg[3][8]  ( .D(n3230), .CK(n4272), .RN(n3741), .QN(n88)
         );
  DFFR_X1 \registers_reg[2][8]  ( .D(n3262), .CK(n4272), .RN(n3744), .QN(n56)
         );
  DFFR_X1 \registers_reg[27][26]  ( .D(n2864), .CK(n4272), .RN(n3673), .QN(
        n838) );
  DFFR_X1 \registers_reg[31][7]  ( .D(n2781), .CK(n4272), .RN(n3659), .QN(n985) );
  DFFR_X1 \registers_reg[30][22]  ( .D(n2828), .CK(n4272), .RN(n3663), .QN(
        n938) );
  DFFR_X1 \registers_reg[30][29]  ( .D(n2835), .CK(n4272), .RN(n3664), .QN(
        n931) );
  DFFR_X1 \registers_reg[11][27]  ( .D(n3121), .CK(n4272), .RN(n3719), .QN(
        n325) );
  DFFR_X1 \registers_reg[11][26]  ( .D(n3120), .CK(n4272), .RN(n3719), .QN(
        n326) );
  DFFR_X1 \registers_reg[11][5]  ( .D(n3099), .CK(n4272), .RN(n3717), .QN(n347) );
  DFFR_X1 \registers_reg[30][0]  ( .D(n2806), .CK(n4272), .RN(n3661), .QN(n960) );
  DFFR_X1 \registers_reg[16][25]  ( .D(n3023), .CK(n4272), .RN(n3704), .QN(
        n487) );
  DFFR_X1 \registers_reg[10][25]  ( .D(n3151), .CK(n4272), .RN(n3722), .QN(
        n295) );
  DFFR_X1 \registers_reg[21][7]  ( .D(n2909), .CK(n4272), .RN(n3688), .QN(n665) );
  DFFR_X1 \registers_reg[14][0]  ( .D(n3062), .CK(n4272), .RN(n3708), .QN(n448) );
  DFFR_X1 \registers_reg[14][11]  ( .D(n3073), .CK(n4272), .RN(n3709), .QN(
        n437) );
  DFFR_X1 \registers_reg[31][22]  ( .D(n2796), .CK(n4272), .RN(n3661), .QN(
        n970) );
  DFFR_X1 \registers_reg[14][26]  ( .D(n3088), .CK(n4272), .RN(n3710), .QN(
        n422) );
  DFFR_X1 \registers_reg[26][2]  ( .D(n2872), .CK(n4272), .RN(n3673), .QN(n830) );
  DFFR_X1 \registers_reg[17][21]  ( .D(n2987), .CK(n4272), .RN(n3701), .QN(
        n523) );
  DFFR_X1 \registers_reg[16][21]  ( .D(n3019), .CK(n4272), .RN(n3704), .QN(
        n491) );
  DFFR_X1 \registers_reg[15][21]  ( .D(n3051), .CK(n4272), .RN(n3707), .QN(
        n459) );
  DFFR_X1 \registers_reg[11][21]  ( .D(n3115), .CK(n4272), .RN(n3719), .QN(
        n331) );
  DFFR_X1 \registers_reg[10][21]  ( .D(n3147), .CK(n4272), .RN(n3722), .QN(
        n299) );
  DFFR_X1 \registers_reg[20][7]  ( .D(n2941), .CK(n4272), .RN(n3691), .QN(n633) );
  DFFR_X1 \registers_reg[30][8]  ( .D(n2814), .CK(n4272), .RN(n3662), .QN(n952) );
  DFFR_X1 \registers_reg[27][4]  ( .D(n2842), .CK(n4272), .RN(n3671), .QN(n860) );
  DFFR_X1 \registers_reg[2][2]  ( .D(n3256), .CK(n4272), .RN(n3743), .QN(n62)
         );
  DFFR_X1 \registers_reg[14][5]  ( .D(n3067), .CK(n4272), .RN(n3708), .QN(n443) );
  DFFR_X1 \registers_reg[26][22]  ( .D(n2892), .CK(n4272), .RN(n3675), .QN(
        n810) );
  DFFR_X1 \registers_reg[3][3]  ( .D(n3225), .CK(n4272), .RN(n3740), .QN(n93)
         );
  DFFR_X1 \registers_reg[11][25]  ( .D(n3119), .CK(n4272), .RN(n3719), .QN(
        n327) );
  DFFR_X1 \registers_reg[17][15]  ( .D(n2981), .CK(n4272), .RN(n3701), .QN(
        n529) );
  DFFR_X1 \registers_reg[30][7]  ( .D(n2813), .CK(n4272), .RN(n3662), .QN(n953) );
  DFFR_X1 \registers_reg[3][31]  ( .D(n3253), .CK(n4272), .RN(n3743), .QN(n65)
         );
  DFFR_X1 \registers_reg[20][0]  ( .D(n2934), .CK(n4272), .RN(n3691), .QN(n640) );
  DFFR_X1 \registers_reg[10][0]  ( .D(n3126), .CK(n4272), .RN(n3720), .QN(n320) );
  DFFR_X1 \registers_reg[21][0]  ( .D(n2902), .CK(n4272), .RN(n3688), .QN(n672) );
  DFFR_X1 \registers_reg[11][0]  ( .D(n3094), .CK(n4272), .RN(n3717), .QN(n352) );
  DFFR_X1 \registers_reg[26][5]  ( .D(n2875), .CK(n4272), .RN(n3674), .QN(n827) );
  DFFR_X1 \registers_reg[10][15]  ( .D(n3141), .CK(n4272), .RN(n3721), .QN(
        n305) );
  DFFR_X1 \registers_reg[10][31]  ( .D(n3157), .CK(n4272), .RN(n3722), .QN(
        n289) );
  DFFR_X1 \registers_reg[27][3]  ( .D(n2841), .CK(n4272), .RN(n3670), .QN(n861) );
  DFFR_X1 \registers_reg[15][15]  ( .D(n3045), .CK(n4272), .RN(n3706), .QN(
        n465) );
  DFFR_X1 \registers_reg[3][11]  ( .D(n3233), .CK(n4272), .RN(n3741), .QN(n85)
         );
  DFFR_X1 \registers_reg[2][11]  ( .D(n3265), .CK(n4272), .RN(n3744), .QN(n53)
         );
  DFFR_X1 \registers_reg[27][0]  ( .D(n2838), .CK(n4272), .RN(n3670), .QN(n864) );
  DFFR_X1 \registers_reg[21][3]  ( .D(n2905), .CK(n4272), .RN(n3688), .QN(n669) );
  DFFR_X1 \registers_reg[3][27]  ( .D(n3249), .CK(n4272), .RN(n3742), .QN(n69)
         );
  DFFR_X1 \registers_reg[3][26]  ( .D(n3248), .CK(n4272), .RN(n3742), .QN(n70)
         );
  DFFR_X1 \registers_reg[3][5]  ( .D(n3227), .CK(n4272), .RN(n3740), .QN(n91)
         );
  DFFR_X1 \registers_reg[2][27]  ( .D(n3281), .CK(n4272), .RN(n3745), .QN(n37)
         );
  DFFR_X1 \registers_reg[2][26]  ( .D(n3280), .CK(n4272), .RN(n3745), .QN(n38)
         );
  DFFR_X1 \registers_reg[2][5]  ( .D(n3259), .CK(n4272), .RN(n3743), .QN(n59)
         );
  DFFR_X1 \registers_reg[31][5]  ( .D(n2779), .CK(n4272), .RN(n3659), .QN(n987) );
  DFFR_X1 \registers_reg[26][0]  ( .D(n2870), .CK(n4272), .RN(n3673), .QN(n832) );
  DFFR_X1 \registers_reg[10][16]  ( .D(n3142), .CK(n4272), .RN(n3721), .QN(
        n304) );
  DFFR_X1 \registers_reg[31][3]  ( .D(n2777), .CK(n4272), .RN(n3659), .QN(n989) );
  DFFR_X1 \registers_reg[5][3]  ( .D(n3161), .CK(n4272), .RN(n3734), .QN(n157)
         );
  DFFR_X1 \registers_reg[14][16]  ( .D(n3078), .CK(n4272), .RN(n3709), .QN(
        n432) );
  DFFR_X1 \registers_reg[14][15]  ( .D(n3077), .CK(n4272), .RN(n3709), .QN(
        n433) );
  DFFR_X1 \registers_reg[26][4]  ( .D(n2874), .CK(n4272), .RN(n3673), .QN(n828) );
  DFFR_X1 \registers_reg[15][16]  ( .D(n3046), .CK(n4272), .RN(n3707), .QN(
        n464) );
  DFFR_X1 \registers_reg[21][2]  ( .D(n2904), .CK(n4272), .RN(n3688), .QN(n670) );
  DFFR_X1 \registers_reg[5][2]  ( .D(n3160), .CK(n4272), .RN(n3734), .QN(n158)
         );
  DFFR_X1 \registers_reg[16][31]  ( .D(n3029), .CK(n4272), .RN(n3705), .QN(
        n481) );
  DFFR_X1 \registers_reg[16][29]  ( .D(n3027), .CK(n4272), .RN(n3705), .QN(
        n483) );
  DFFR_X1 \registers_reg[16][15]  ( .D(n3013), .CK(n4272), .RN(n3704), .QN(
        n497) );
  DFFR_X1 \registers_reg[16][2]  ( .D(n3000), .CK(n4272), .RN(n3702), .QN(n510) );
  DFFR_X1 \registers_reg[3][4]  ( .D(n3226), .CK(n4272), .RN(n3740), .QN(n92)
         );
  DFFR_X1 \registers_reg[2][4]  ( .D(n3258), .CK(n4272), .RN(n3743), .QN(n60)
         );
  DFFR_X1 \registers_reg[17][16]  ( .D(n2982), .CK(n4272), .RN(n3701), .QN(
        n528) );
  DFFR_X1 \registers_reg[21][26]  ( .D(n2928), .CK(n4272), .RN(n3690), .QN(
        n646) );
  DFFR_X1 \registers_reg[21][5]  ( .D(n2907), .CK(n4272), .RN(n3688), .QN(n667) );
  DFFR_X1 \registers_reg[5][27]  ( .D(n3185), .CK(n4272), .RN(n3737), .QN(n133) );
  DFFR_X1 \registers_reg[5][5]  ( .D(n3163), .CK(n4272), .RN(n3735), .QN(n155)
         );
  DFFR_X1 \registers_reg[30][10]  ( .D(n2816), .CK(n4272), .RN(n3662), .QN(
        n950) );
  DFFR_X1 \registers_reg[30][31]  ( .D(n2837), .CK(n4272), .RN(n3664), .QN(
        n929) );
  DFFR_X1 \registers_reg[14][14]  ( .D(n3076), .CK(n4272), .RN(n3709), .QN(
        n434) );
  DFFR_X1 \registers_reg[3][21]  ( .D(n3243), .CK(n4272), .RN(n3742), .QN(n75)
         );
  DFFR_X1 \registers_reg[2][21]  ( .D(n3275), .CK(n4272), .RN(n3745), .QN(n43)
         );
  DFFR_X1 \registers_reg[14][18]  ( .D(n3080), .CK(n4272), .RN(n3710), .QN(
        n430) );
  DFFR_X1 \registers_reg[16][7]  ( .D(n3005), .CK(n4272), .RN(n3703), .QN(n505) );
  DFFR_X1 \registers_reg[16][6]  ( .D(n3004), .CK(n4272), .RN(n3703), .QN(n506) );
  DFFR_X1 \registers_reg[16][0]  ( .D(n2998), .CK(n4272), .RN(n3702), .QN(n512) );
  DFFR_X1 \registers_reg[16][28]  ( .D(n3026), .CK(n4272), .RN(n3705), .QN(
        n484) );
  DFFR_X1 \registers_reg[26][31]  ( .D(n2901), .CK(n4272), .RN(n3676), .QN(
        n801) );
  DFFR_X1 \registers_reg[16][17]  ( .D(n3015), .CK(n4272), .RN(n3704), .QN(
        n495) );
  DFFR_X1 \registers_reg[17][27]  ( .D(n2993), .CK(n4272), .RN(n3702), .QN(
        n517) );
  DFFR_X1 \registers_reg[17][26]  ( .D(n2992), .CK(n4272), .RN(n3702), .QN(
        n518) );
  DFFR_X1 \registers_reg[21][11]  ( .D(n2913), .CK(n4272), .RN(n3689), .QN(
        n661) );
  DFFR_X1 \registers_reg[17][25]  ( .D(n2991), .CK(n4272), .RN(n3702), .QN(
        n519) );
  DFFR_X1 \registers_reg[17][24]  ( .D(n2990), .CK(n4272), .RN(n3701), .QN(
        n520) );
  DFFR_X1 \registers_reg[4][27]  ( .D(n3217), .CK(n4272), .RN(n3740), .QN(n101) );
  DFFR_X1 \registers_reg[30][5]  ( .D(n2811), .CK(n4272), .RN(n3662), .QN(n955) );
  DFFR_X1 \registers_reg[21][27]  ( .D(n2929), .CK(n4272), .RN(n3690), .QN(
        n645) );
  DFFR_X1 \registers_reg[5][26]  ( .D(n3184), .CK(n4272), .RN(n3737), .QN(n134) );
  DFFR_X1 \registers_reg[20][27]  ( .D(n2961), .CK(n4272), .RN(n3693), .QN(
        n613) );
  DFFR_X1 \registers_reg[2][3]  ( .D(n3257), .CK(n4272), .RN(n3743), .QN(n61)
         );
  DFFR_X1 \registers_reg[5][25]  ( .D(n3183), .CK(n4272), .RN(n3736), .QN(n135) );
  DFFR_X1 \registers_reg[26][11]  ( .D(n2881), .CK(n4272), .RN(n3674), .QN(
        n821) );
  DFFR_X1 \registers_reg[30][4]  ( .D(n2810), .CK(n4272), .RN(n3662), .QN(n956) );
  DFFR_X1 \registers_reg[21][8]  ( .D(n2910), .CK(n4272), .RN(n3688), .QN(n664) );
  DFFR_X1 \registers_reg[5][8]  ( .D(n3166), .CK(n4272), .RN(n3735), .QN(n152)
         );
  DFFR_X1 \registers_reg[20][8]  ( .D(n2942), .CK(n4272), .RN(n3691), .QN(n632) );
  DFFR_X1 \registers_reg[15][17]  ( .D(n3047), .CK(n4272), .RN(n3707), .QN(
        n463) );
  DFFR_X1 \registers_reg[16][30]  ( .D(n3028), .CK(n4272), .RN(n3705), .QN(
        n482) );
  DFFR_X1 \registers_reg[17][17]  ( .D(n2983), .CK(n4272), .RN(n3701), .QN(
        n527) );
  DFFR_X1 \registers_reg[30][23]  ( .D(n2829), .CK(n4272), .RN(n3664), .QN(
        n937) );
  DFFR_X1 \registers_reg[30][26]  ( .D(n2832), .CK(n4272), .RN(n3664), .QN(
        n934) );
  DFFR_X1 \registers_reg[30][28]  ( .D(n2834), .CK(n4272), .RN(n3664), .QN(
        n932) );
  DFFR_X1 \registers_reg[3][28]  ( .D(n3250), .CK(n4272), .RN(n3743), .QN(n68)
         );
  DFFR_X1 \registers_reg[3][14]  ( .D(n3236), .CK(n4272), .RN(n3741), .QN(n82)
         );
  DFFR_X1 \registers_reg[2][28]  ( .D(n3282), .CK(n4272), .RN(n3745), .QN(n36)
         );
  DFFR_X1 \registers_reg[2][14]  ( .D(n3268), .CK(n4272), .RN(n3744), .QN(n50)
         );
  DFFR_X1 \registers_reg[10][14]  ( .D(n3140), .CK(n4272), .RN(n3721), .QN(
        n306) );
  DFFR_X1 \registers_reg[16][14]  ( .D(n3012), .CK(n4272), .RN(n3703), .QN(
        n498) );
  DFFR_X1 \registers_reg[10][28]  ( .D(n3154), .CK(n4272), .RN(n3722), .QN(
        n292) );
  DFFR_X1 \registers_reg[26][27]  ( .D(n2897), .CK(n4272), .RN(n3676), .QN(
        n805) );
  DFFR_X1 \registers_reg[26][26]  ( .D(n2896), .CK(n4272), .RN(n3675), .QN(
        n806) );
  DFFR_X1 \registers_reg[16][18]  ( .D(n3016), .CK(n4272), .RN(n3704), .QN(
        n494) );
  DFFR_X1 \registers_reg[15][14]  ( .D(n3044), .CK(n4272), .RN(n3706), .QN(
        n466) );
  DFFR_X1 \registers_reg[17][28]  ( .D(n2994), .CK(n4272), .RN(n3702), .QN(
        n516) );
  DFFR_X1 \registers_reg[3][23]  ( .D(n3245), .CK(n4272), .RN(n3742), .QN(n73)
         );
  DFFR_X1 \registers_reg[2][23]  ( .D(n3277), .CK(n4272), .RN(n3745), .QN(n41)
         );
  DFFR_X1 \registers_reg[4][23]  ( .D(n3213), .CK(n4272), .RN(n3739), .QN(n105) );
  DFFR_X1 \registers_reg[5][23]  ( .D(n3181), .CK(n4272), .RN(n3736), .QN(n137) );
  DFFR_X1 \registers_reg[17][23]  ( .D(n2989), .CK(n4272), .RN(n3701), .QN(
        n521) );
  DFFR_X1 \registers_reg[15][18]  ( .D(n3048), .CK(n4272), .RN(n3707), .QN(
        n462) );
  DFFR_X1 \registers_reg[21][4]  ( .D(n2906), .CK(n4272), .RN(n3688), .QN(n668) );
  DFFR_X1 \registers_reg[5][4]  ( .D(n3162), .CK(n4272), .RN(n3735), .QN(n156)
         );
  DFFR_X1 \registers_reg[26][8]  ( .D(n2878), .CK(n4272), .RN(n3674), .QN(n824) );
  DFFR_X1 \registers_reg[30][1]  ( .D(n2807), .CK(n4272), .RN(n3662), .QN(n959) );
  DFFR_X1 \registers_reg[2][6]  ( .D(n3260), .CK(n4272), .RN(n3743), .QN(n58)
         );
  DFFR_X1 \registers_reg[3][18]  ( .D(n3240), .CK(n4272), .RN(n3742), .QN(n78)
         );
  DFFR_X1 \registers_reg[2][18]  ( .D(n3272), .CK(n4272), .RN(n3745), .QN(n46)
         );
  DFFR_X1 \registers_reg[2][9]  ( .D(n3263), .CK(n4272), .RN(n3744), .QN(n55)
         );
  DFFR_X1 \registers_reg[10][1]  ( .D(n3127), .CK(n4272), .RN(n3720), .QN(n319) );
  DFFR_X1 \registers_reg[21][18]  ( .D(n2920), .CK(n4272), .RN(n3689), .QN(
        n654) );
  DFFR_X1 \registers_reg[21][10]  ( .D(n2912), .CK(n4272), .RN(n3689), .QN(
        n662) );
  DFFR_X1 \registers_reg[21][9]  ( .D(n2911), .CK(n4272), .RN(n3688), .QN(n663) );
  DFFR_X1 \registers_reg[21][1]  ( .D(n2903), .CK(n4272), .RN(n3688), .QN(n671) );
  DFFR_X1 \registers_reg[5][13]  ( .D(n3171), .CK(n4272), .RN(n3735), .QN(n147) );
  DFFR_X1 \registers_reg[5][6]  ( .D(n3164), .CK(n4272), .RN(n3735), .QN(n154)
         );
  DFFR_X1 \registers_reg[17][18]  ( .D(n2984), .CK(n4272), .RN(n3701), .QN(
        n526) );
  DFFR_X1 \registers_reg[17][13]  ( .D(n2979), .CK(n4272), .RN(n3700), .QN(
        n531) );
  DFFR_X1 \registers_reg[17][9]  ( .D(n2975), .CK(n4272), .RN(n3700), .QN(n535) );
  DFFR_X1 \registers_reg[17][6]  ( .D(n2972), .CK(n4272), .RN(n3700), .QN(n538) );
  DFFR_X1 \registers_reg[11][1]  ( .D(n3095), .CK(n4272), .RN(n3717), .QN(n351) );
  DFFR_X1 \registers_reg[10][18]  ( .D(n3144), .CK(n4272), .RN(n3721), .QN(
        n302) );
  DFFR_X1 \registers_reg[10][13]  ( .D(n3139), .CK(n4272), .RN(n3721), .QN(
        n307) );
  DFFR_X1 \registers_reg[17][10]  ( .D(n2976), .CK(n4272), .RN(n3700), .QN(
        n534) );
  DFFR_X1 \registers_reg[16][1]  ( .D(n2999), .CK(n4272), .RN(n3702), .QN(n511) );
  DFFR_X1 \registers_reg[11][10]  ( .D(n3104), .CK(n4272), .RN(n3718), .QN(
        n342) );
  DFFR_X1 \registers_reg[10][10]  ( .D(n3136), .CK(n4272), .RN(n3721), .QN(
        n310) );
  DFFR_X1 \registers_reg[10][9]  ( .D(n3135), .CK(n4272), .RN(n3720), .QN(n311) );
  DFFR_X1 \registers_reg[10][6]  ( .D(n3132), .CK(n4272), .RN(n3720), .QN(n314) );
  DFFR_X1 \registers_reg[26][23]  ( .D(n2893), .CK(n4272), .RN(n3675), .QN(
        n809) );
  DFFR_X1 \registers_reg[14][23]  ( .D(n3085), .CK(n4272), .RN(n3710), .QN(
        n425) );
  DFFR_X1 \registers_reg[15][9]  ( .D(n3039), .CK(n4272), .RN(n3706), .QN(n471) );
  DFFR_X1 \registers_reg[15][13]  ( .D(n3043), .CK(n4272), .RN(n3706), .QN(
        n467) );
  DFFR_X1 \registers_reg[16][16]  ( .D(n3014), .CK(n4272), .RN(n3704), .QN(
        n496) );
  DFFR_X1 \registers_reg[15][6]  ( .D(n3036), .CK(n4272), .RN(n3706), .QN(n474) );
  DFFR_X1 \registers_reg[26][28]  ( .D(n2898), .CK(n4272), .RN(n3676), .QN(
        n804) );
  DFFR_X1 \registers_reg[26][14]  ( .D(n2884), .CK(n4272), .RN(n3674), .QN(
        n818) );
  DFFR_X1 \registers_reg[27][18]  ( .D(n2856), .CK(n4272), .RN(n3672), .QN(
        n846) );
  DFFR_X1 \registers_reg[17][20]  ( .D(n2986), .CK(n4272), .RN(n3701), .QN(
        n524) );
  DFFR_X1 \registers_reg[16][20]  ( .D(n3018), .CK(n4272), .RN(n3704), .QN(
        n492) );
  DFFR_X1 \registers_reg[15][20]  ( .D(n3050), .CK(n4272), .RN(n3707), .QN(
        n460) );
  DFFR_X1 \registers_reg[30][27]  ( .D(n2833), .CK(n4272), .RN(n3664), .QN(
        n933) );
  DFFR_X1 \registers_reg[21][21]  ( .D(n2923), .CK(n4272), .RN(n3690), .QN(
        n651) );
  DFFR_X1 \registers_reg[5][21]  ( .D(n3179), .CK(n4272), .RN(n3736), .QN(n139) );
  DFFR_X1 \registers_reg[26][18]  ( .D(n2888), .CK(n4272), .RN(n3675), .QN(
        n814) );
  DFFR_X1 \registers_reg[16][5]  ( .D(n3003), .CK(n4272), .RN(n3703), .QN(n507) );
  DFFR_X1 \registers_reg[16][3]  ( .D(n3001), .CK(n4272), .RN(n3702), .QN(n509) );
  DFFR_X1 \registers_reg[2][31]  ( .D(n3285), .CK(n4272), .RN(n3746), .QN(n33)
         );
  DFFR_X1 \registers_reg[20][31]  ( .D(n2965), .CK(n4272), .RN(n3693), .QN(
        n609) );
  DFFR_X1 \registers_reg[20][25]  ( .D(n2959), .CK(n4272), .RN(n3693), .QN(
        n615) );
  DFFR_X1 \registers_reg[20][21]  ( .D(n2955), .CK(n4272), .RN(n3692), .QN(
        n619) );
  DFFR_X1 \registers_reg[20][20]  ( .D(n2954), .CK(n4272), .RN(n3692), .QN(
        n620) );
  DFFR_X1 \registers_reg[20][15]  ( .D(n2949), .CK(n4272), .RN(n3692), .QN(
        n625) );
  DFFR_X1 \registers_reg[20][13]  ( .D(n2947), .CK(n4272), .RN(n3692), .QN(
        n627) );
  DFFR_X1 \registers_reg[20][6]  ( .D(n2940), .CK(n4272), .RN(n3691), .QN(n634) );
  DFFR_X1 \registers_reg[20][5]  ( .D(n2939), .CK(n4272), .RN(n3691), .QN(n635) );
  DFFR_X1 \registers_reg[3][15]  ( .D(n3237), .CK(n4272), .RN(n3741), .QN(n81)
         );
  DFFR_X1 \registers_reg[2][24]  ( .D(n3278), .CK(n4272), .RN(n3745), .QN(n40)
         );
  DFFR_X1 \registers_reg[20][24]  ( .D(n2958), .CK(n4272), .RN(n3693), .QN(
        n616) );
  DFFR_X1 \registers_reg[21][24]  ( .D(n2926), .CK(n4272), .RN(n3690), .QN(
        n648) );
  DFFR_X1 \registers_reg[5][24]  ( .D(n3182), .CK(n4272), .RN(n3736), .QN(n136) );
  DFFR_X1 \registers_reg[11][24]  ( .D(n3118), .CK(n4272), .RN(n3719), .QN(
        n328) );
  DFFR_X1 \registers_reg[14][17]  ( .D(n3079), .CK(n4272), .RN(n3710), .QN(
        n431) );
  DFFR_X1 \registers_reg[5][31]  ( .D(n3189), .CK(n4272), .RN(n3737), .QN(n129) );
  DFFR_X1 \registers_reg[20][30]  ( .D(n2964), .CK(n4272), .RN(n3693), .QN(
        n610) );
  DFFR_X1 \registers_reg[20][29]  ( .D(n2963), .CK(n4272), .RN(n3693), .QN(
        n611) );
  DFFR_X1 \registers_reg[20][28]  ( .D(n2962), .CK(n4272), .RN(n3693), .QN(
        n612) );
  DFFR_X1 \registers_reg[20][26]  ( .D(n2960), .CK(n4272), .RN(n3693), .QN(
        n614) );
  DFFR_X1 \registers_reg[20][19]  ( .D(n2953), .CK(n4272), .RN(n3692), .QN(
        n621) );
  DFFR_X1 \registers_reg[20][18]  ( .D(n2952), .CK(n4272), .RN(n3692), .QN(
        n622) );
  DFFR_X1 \registers_reg[20][14]  ( .D(n2948), .CK(n4272), .RN(n3692), .QN(
        n626) );
  DFFR_X1 \registers_reg[20][11]  ( .D(n2945), .CK(n4272), .RN(n3692), .QN(
        n629) );
  DFFR_X1 \registers_reg[20][10]  ( .D(n2944), .CK(n4272), .RN(n3691), .QN(
        n630) );
  DFFR_X1 \registers_reg[20][4]  ( .D(n2938), .CK(n4272), .RN(n3691), .QN(n636) );
  DFFR_X1 \registers_reg[20][3]  ( .D(n2937), .CK(n4272), .RN(n3691), .QN(n637) );
  DFFR_X1 \registers_reg[20][2]  ( .D(n2936), .CK(n4272), .RN(n3691), .QN(n638) );
  DFFR_X1 \registers_reg[20][1]  ( .D(n2935), .CK(n4272), .RN(n3691), .QN(n639) );
  DFFR_X1 \registers_reg[30][3]  ( .D(n2809), .CK(n4272), .RN(n3662), .QN(n957) );
  DFFR_X1 \registers_reg[16][24]  ( .D(n3022), .CK(n4272), .RN(n3704), .QN(
        n488) );
  DFFR_X1 \registers_reg[11][2]  ( .D(n3096), .CK(n4272), .RN(n3717), .QN(n350) );
  DFFR_X1 \registers_reg[14][2]  ( .D(n3064), .CK(n4272), .RN(n3708), .QN(n446) );
  DFFR_X1 \registers_reg[30][16]  ( .D(n2822), .CK(n4272), .RN(n3663), .QN(
        n944) );
  DFFR_X1 \registers_reg[30][15]  ( .D(n2821), .CK(n4272), .RN(n3663), .QN(
        n945) );
  DFFR_X1 \registers_reg[5][15]  ( .D(n3173), .CK(n4272), .RN(n3736), .QN(n145) );
  DFFR_X1 \registers_reg[3][17]  ( .D(n3239), .CK(n4272), .RN(n3742), .QN(n79)
         );
  DFFR_X1 \registers_reg[10][17]  ( .D(n3143), .CK(n4272), .RN(n3721), .QN(
        n303) );
  DFFR_X1 \registers_reg[16][19]  ( .D(n3017), .CK(n4272), .RN(n3704), .QN(
        n493) );
  DFFR_X1 \registers_reg[11][19]  ( .D(n3113), .CK(n4272), .RN(n3718), .QN(
        n333) );
  DFFR_X1 \registers_reg[21][16]  ( .D(n2918), .CK(n4272), .RN(n3689), .QN(
        n656) );
  DFFR_X1 \registers_reg[5][16]  ( .D(n3174), .CK(n4272), .RN(n3736), .QN(n144) );
  DFFR_X1 \registers_reg[31][16]  ( .D(n2790), .CK(n4272), .RN(n3660), .QN(
        n976) );
  DFFR_X1 \registers_reg[31][8]  ( .D(n2782), .CK(n4272), .RN(n3659), .QN(n984) );
  DFFR_X1 \registers_reg[31][9]  ( .D(n2783), .CK(n4272), .RN(n3659), .QN(n983) );
  DFFR_X1 \registers_reg[31][31]  ( .D(n2805), .CK(n4272), .RN(n3661), .QN(
        n961) );
  DFFR_X1 \registers_reg[31][27]  ( .D(n2801), .CK(n4272), .RN(n3661), .QN(
        n965) );
  DFFR_X1 \registers_reg[31][21]  ( .D(n2795), .CK(n4272), .RN(n3660), .QN(
        n971) );
  DFFR_X1 \registers_reg[31][19]  ( .D(n2793), .CK(n4272), .RN(n3660), .QN(
        n973) );
  DFFR_X1 \registers_reg[31][17]  ( .D(n2791), .CK(n4272), .RN(n3660), .QN(
        n975) );
  DFFR_X1 \registers_reg[31][14]  ( .D(n2788), .CK(n4272), .RN(n3660), .QN(
        n978) );
  DFFR_X1 \registers_reg[31][0]  ( .D(n2774), .CK(n4272), .RN(n3659), .QN(n992) );
  DFFR_X1 \registers_reg[30][24]  ( .D(n2830), .CK(n4272), .RN(n3664), .QN(
        n936) );
  DFFR_X1 \registers_reg[26][16]  ( .D(n2886), .CK(n4272), .RN(n3675), .QN(
        n816) );
  DFFR_X1 \registers_reg[16][4]  ( .D(n3002), .CK(n4272), .RN(n3703), .QN(n508) );
  DFFR_X1 \registers_reg[17][4]  ( .D(n2970), .CK(n4272), .RN(n3700), .QN(n540) );
  DFFR_X1 \registers_reg[20][17]  ( .D(n2951), .CK(n4272), .RN(n3692), .QN(
        n623) );
  DFFR_X1 \registers_reg[3][16]  ( .D(n3238), .CK(n4272), .RN(n3741), .QN(n80)
         );
  DFFR_X1 \registers_reg[2][16]  ( .D(n3270), .CK(n4272), .RN(n3744), .QN(n48)
         );
  DFFR_X1 \registers_reg[27][31]  ( .D(n2869), .CK(n4272), .RN(n3673), .QN(
        n833) );
  DFFR_X1 \registers_reg[31][30]  ( .D(n2804), .CK(n4272), .RN(n3661), .QN(
        n962) );
  DFFR_X1 \registers_reg[15][4]  ( .D(n3034), .CK(n4272), .RN(n3705), .QN(n476) );
  DFFR_X1 \registers_reg[31][29]  ( .D(n2803), .CK(n4272), .RN(n3661), .QN(
        n963) );
  DFFR_X1 \registers_reg[31][28]  ( .D(n2802), .CK(n4272), .RN(n3661), .QN(
        n964) );
  DFFR_X1 \registers_reg[31][26]  ( .D(n2800), .CK(n4272), .RN(n3661), .QN(
        n966) );
  DFFR_X1 \registers_reg[31][15]  ( .D(n2789), .CK(n4272), .RN(n3660), .QN(
        n977) );
  DFFR_X1 \registers_reg[31][13]  ( .D(n2787), .CK(n4272), .RN(n3660), .QN(
        n979) );
  DFFR_X1 \registers_reg[31][12]  ( .D(n2786), .CK(n4272), .RN(n3660), .QN(
        n980) );
  DFFR_X1 \registers_reg[31][11]  ( .D(n2785), .CK(n4272), .RN(n3660), .QN(
        n981) );
  DFFR_X1 \registers_reg[31][10]  ( .D(n2784), .CK(n4272), .RN(n3659), .QN(
        n982) );
  DFFR_X1 \registers_reg[31][6]  ( .D(n2780), .CK(n4272), .RN(n3659), .QN(n986) );
  DFFR_X1 \registers_reg[31][1]  ( .D(n2775), .CK(n4272), .RN(n3659), .QN(n991) );
  DFFR_X1 \registers_reg[27][27]  ( .D(n2865), .CK(n4272), .RN(n3673), .QN(
        n837) );
  DFFR_X1 \registers_reg[27][23]  ( .D(n2861), .CK(n4272), .RN(n3672), .QN(
        n841) );
  DFFR_X1 \registers_reg[27][17]  ( .D(n2855), .CK(n4272), .RN(n3672), .QN(
        n847) );
  DFFR_X1 \registers_reg[27][16]  ( .D(n2854), .CK(n4272), .RN(n3672), .QN(
        n848) );
  DFFR_X1 \registers_reg[27][15]  ( .D(n2853), .CK(n4272), .RN(n3672), .QN(
        n849) );
  DFFR_X1 \registers_reg[27][14]  ( .D(n2852), .CK(n4272), .RN(n3671), .QN(
        n850) );
  DFFR_X1 \registers_reg[27][13]  ( .D(n2851), .CK(n4272), .RN(n3671), .QN(
        n851) );
  DFFR_X1 \registers_reg[27][11]  ( .D(n2849), .CK(n4272), .RN(n3671), .QN(
        n853) );
  DFFR_X1 \registers_reg[27][9]  ( .D(n2847), .CK(n4272), .RN(n3671), .QN(n855) );
  DFFR_X1 \registers_reg[27][8]  ( .D(n2846), .CK(n4272), .RN(n3671), .QN(n856) );
  DFFR_X1 \registers_reg[27][6]  ( .D(n2844), .CK(n4272), .RN(n3671), .QN(n858) );
  DFFR_X1 \registers_reg[27][5]  ( .D(n2843), .CK(n4272), .RN(n3671), .QN(n859) );
  DFFR_X1 \registers_reg[31][20]  ( .D(n2794), .CK(n4272), .RN(n3660), .QN(
        n972) );
  DFFR_X1 \registers_reg[30][17]  ( .D(n2823), .CK(n4272), .RN(n3663), .QN(
        n943) );
  DFFR_X1 \registers_reg[21][17]  ( .D(n2919), .CK(n4272), .RN(n3689), .QN(
        n655) );
  DFFR_X1 \registers_reg[26][17]  ( .D(n2887), .CK(n4272), .RN(n3675), .QN(
        n815) );
  DFFR_X1 \registers_reg[15][24]  ( .D(n3054), .CK(n4272), .RN(n3707), .QN(
        n456) );
  DFFR_X1 \registers_reg[26][24]  ( .D(n2894), .CK(n4272), .RN(n3675), .QN(
        n808) );
  DFFR_X1 \registers_reg[27][24]  ( .D(n2862), .CK(n4272), .RN(n3672), .QN(
        n840) );
  DFFR_X1 \registers_reg[14][24]  ( .D(n3086), .CK(n4272), .RN(n3710), .QN(
        n424) );
  DFFR_X1 \registers_reg[20][16]  ( .D(n2950), .CK(n4272), .RN(n3692), .QN(
        n624) );
  DFFR_X1 \registers_reg[31][2]  ( .D(n2776), .CK(n4272), .RN(n3659), .QN(n990) );
  DFFR_X1 \registers_reg[3][2]  ( .D(n3224), .CK(n4272), .RN(n3740), .QN(n94)
         );
  DFFR_X1 \registers_reg[31][23]  ( .D(n2797), .CK(n4272), .RN(n3661), .QN(
        n969) );
  DFFR_X1 \registers_reg[31][18]  ( .D(n2792), .CK(n4272), .RN(n3660), .QN(
        n974) );
  DFFR_X1 \registers_reg[14][4]  ( .D(n3066), .CK(n4272), .RN(n3708), .QN(n444) );
  DFFR_X1 \registers_reg[10][3]  ( .D(n3129), .CK(n4272), .RN(n3720), .QN(n317) );
  DFFR_X1 \registers_reg[3][0]  ( .D(n3222), .CK(n4272), .RN(n3740), .QN(n96)
         );
  DFFR_X1 \registers_reg[2][0]  ( .D(n3254), .CK(n4272), .RN(n3743), .QN(n64)
         );
  DFFR_X1 \registers_reg[5][0]  ( .D(n3158), .CK(n4272), .RN(n3734), .QN(n160)
         );
  DFFR_X1 \registers_reg[17][0]  ( .D(n2966), .CK(n4272), .RN(n3699), .QN(n544) );
  DFFR_X1 \registers_reg[17][22]  ( .D(n2988), .CK(n4272), .RN(n3701), .QN(
        n522) );
  DFFR_X1 \registers_reg[17][7]  ( .D(n2973), .CK(n4272), .RN(n3700), .QN(n537) );
  DFFR_X1 \registers_reg[16][22]  ( .D(n3020), .CK(n4272), .RN(n3704), .QN(
        n490) );
  DFFR_X1 \registers_reg[15][22]  ( .D(n3052), .CK(n4272), .RN(n3707), .QN(
        n458) );
  DFFR_X1 \registers_reg[15][7]  ( .D(n3037), .CK(n4272), .RN(n3706), .QN(n473) );
  DFFR_X1 \registers_reg[11][22]  ( .D(n3116), .CK(n4272), .RN(n3719), .QN(
        n330) );
  DFFR_X1 \registers_reg[10][22]  ( .D(n3148), .CK(n4272), .RN(n3722), .QN(
        n298) );
  DFFR_X1 \registers_reg[15][0]  ( .D(n3030), .CK(n4272), .RN(n3705), .QN(n480) );
  DFFR_X1 \registers_reg[11][31]  ( .D(n3125), .CK(n4272), .RN(n3720), .QN(
        n321) );
  DFFR_X1 \registers_reg[2][17]  ( .D(n3271), .CK(n4272), .RN(n3744), .QN(n47)
         );
  DFFR_X1 \registers_reg[3][19]  ( .D(n3241), .CK(n4272), .RN(n3742), .QN(n77)
         );
  DFFR_X1 \registers_reg[30][30]  ( .D(n2836), .CK(n4272), .RN(n3664), .QN(
        n930) );
  DFFR_X1 \registers_reg[27][30]  ( .D(n2868), .CK(n4272), .RN(n3673), .QN(
        n834) );
  DFFR_X1 \registers_reg[2][30]  ( .D(n3284), .CK(n4272), .RN(n3746), .QN(n34)
         );
  DFFR_X1 \registers_reg[11][7]  ( .D(n3101), .CK(n4272), .RN(n3717), .QN(n345) );
  DFFR_X1 \registers_reg[11][6]  ( .D(n3100), .CK(n4272), .RN(n3717), .QN(n346) );
  DFFR_X1 \registers_reg[30][2]  ( .D(n2808), .CK(n4272), .RN(n3662), .QN(n958) );
  DFFR_X1 \registers_reg[22][12]  ( .D(n251), .CK(n4272), .RN(n3686), .Q(
        \registers[22][12] ), .QN(n252) );
  DFFR_X1 \registers_reg[6][15]  ( .D(n406), .CK(n4272), .RN(n3733), .Q(
        \registers[6][15] ), .QN(n407) );
  DFFR_X1 \registers_reg[8][18]  ( .D(n385), .CK(n4272), .RN(n3727), .Q(
        \registers[8][18] ), .QN(n386) );
  DFFR_X1 \registers_reg[29][24]  ( .D(n272), .CK(n4272), .RN(n3667), .Q(
        \registers[29][24] ), .QN(n273) );
  DFFR_X1 \registers_reg[9][14]  ( .D(n257), .CK(n4272), .RN(n3724), .Q(
        \registers[9][14] ), .QN(n258) );
  DFFR_X1 \registers_reg[24][21]  ( .D(n255), .CK(n4272), .RN(n3681), .Q(
        \registers[24][21] ), .QN(n256) );
  DFFR_X1 \registers_reg[13][15]  ( .D(n391), .CK(n4272), .RN(n3712), .Q(
        \registers[13][15] ), .QN(n392) );
  DFFR_X1 \registers_reg[22][20]  ( .D(n404), .CK(n4272), .RN(n3687), .Q(
        \registers[22][20] ), .QN(n405) );
  DFFR_X1 \registers_reg[22][22]  ( .D(n253), .CK(n4272), .RN(n3687), .Q(
        \registers[22][22] ), .QN(n254) );
  DFFR_X1 \registers_reg[12][12]  ( .D(n694), .CK(n4272), .RN(n3715), .Q(
        \registers[12][12] ), .QN(n695) );
  DFFR_X1 \registers_reg[23][3]  ( .D(n685), .CK(n4272), .RN(n3682), .Q(
        \registers[23][3] ), .QN(n686) );
  DFFR_X2 \registers_reg[28][24]  ( .D(n4194), .CK(n4272), .RN(n3669), .Q(
        \registers[28][24] ) );
  DFFR_X2 \registers_reg[8][24]  ( .D(n3789), .CK(n4272), .RN(n3728), .Q(
        \registers[8][24] ) );
  DFFR_X2 \registers_reg[23][24]  ( .D(n4101), .CK(n4272), .RN(n3684), .Q(
        \registers[23][24] ) );
  DFFR_X2 \registers_reg[19][24]  ( .D(n4042), .CK(n4272), .RN(n3696), .Q(
        \registers[19][24] ) );
  DFFR_X1 \registers_reg[6][9]  ( .D(n3931), .CK(n4272), .RN(n3732), .Q(
        \registers[6][9] ) );
  DFFR_X1 \registers_reg[6][11]  ( .D(n3933), .CK(n4272), .RN(n3732), .Q(
        \registers[6][11] ) );
  DFFR_X1 \registers_reg[6][17]  ( .D(n3938), .CK(n4272), .RN(n3733), .Q(
        \registers[6][17] ) );
  DFFR_X1 \registers_reg[6][19]  ( .D(n3940), .CK(n4272), .RN(n3733), .Q(
        \registers[6][19] ) );
  DFFR_X1 \registers_reg[6][20]  ( .D(n3941), .CK(n4272), .RN(n3733), .Q(
        \registers[6][20] ) );
  DFFR_X1 \registers_reg[6][22]  ( .D(n3943), .CK(n4272), .RN(n3733), .Q(
        \registers[6][22] ) );
  DFFR_X1 \registers_reg[6][31]  ( .D(n3952), .CK(n4272), .RN(n3734), .Q(
        \registers[6][31] ) );
  DFFR_X2 \registers_reg[7][24]  ( .D(n3977), .CK(n4272), .RN(n3731), .Q(
        \registers[7][24] ) );
  DFFR_X2 \registers_reg[9][24]  ( .D(n3820), .CK(n4272), .RN(n3725), .Q(
        \registers[9][24] ) );
  DFFR_X2 \registers_reg[1][24]  ( .D(n3914), .CK(n4272), .RN(n3748), .Q(
        \registers[1][24] ) );
  DFFR_X2 \registers_reg[4][8]  ( .D(n3198), .CK(n4272), .RN(n3738), .QN(n120)
         );
  DFFR_X2 \registers_reg[25][30]  ( .D(n4169), .CK(n4272), .RN(n3679), .Q(
        \registers[25][30] ) );
  DFFR_X2 \registers_reg[9][30]  ( .D(n3826), .CK(n4272), .RN(n3725), .Q(
        \registers[9][30] ) );
  DFFR_X2 \registers_reg[1][30]  ( .D(n3920), .CK(n4272), .RN(n3749), .Q(
        \registers[1][30] ) );
  DFFR_X2 \registers_reg[28][30]  ( .D(n4200), .CK(n4272), .RN(n3670), .Q(
        \registers[28][30] ) );
  BUF_X1 U2 ( .A(n874), .Z(n411) );
  CLKBUF_X1 U3 ( .A(n874), .Z(n410) );
  INV_X1 U4 ( .A(n786), .ZN(n1) );
  INV_X1 U5 ( .A(net38967), .ZN(n2) );
  BUF_X1 U6 ( .A(n3604), .Z(n3600) );
  BUF_X1 U7 ( .A(n3574), .Z(n3) );
  CLKBUF_X1 U8 ( .A(n3574), .Z(n31) );
  INV_X1 U9 ( .A(n790), .ZN(n4) );
  INV_X1 U10 ( .A(n865), .ZN(n5) );
  BUF_X2 U11 ( .A(DATAIN[8]), .Z(n30) );
  INV_X2 U12 ( .A(n1282), .ZN(n754) );
  BUF_X2 U13 ( .A(n3579), .Z(n3576) );
  INV_X1 U14 ( .A(n881), .ZN(n6) );
  BUF_X1 U15 ( .A(n1489), .Z(n3507) );
  INV_X1 U16 ( .A(n788), .ZN(n7) );
  CLKBUF_X3 U17 ( .A(n176), .Z(n8) );
  INV_X1 U18 ( .A(n792), .ZN(n9) );
  INV_X1 U19 ( .A(n878), .ZN(n10) );
  INV_X1 U20 ( .A(ADD_WR[0]), .ZN(n11) );
  BUF_X1 U21 ( .A(n3317), .Z(n3619) );
  BUF_X1 U22 ( .A(n3317), .Z(n3617) );
  BUF_X1 U23 ( .A(n3317), .Z(n3618) );
  BUF_X1 U24 ( .A(n3317), .Z(n3621) );
  BUF_X2 U25 ( .A(DATAIN[30]), .Z(n394) );
  BUF_X2 U26 ( .A(DATAIN[30]), .Z(n800) );
  BUF_X1 U27 ( .A(n1180), .Z(n3594) );
  BUF_X1 U28 ( .A(n1180), .Z(n3593) );
  BUF_X1 U29 ( .A(n3604), .Z(n3598) );
  INV_X1 U30 ( .A(net38967), .ZN(n12) );
  BUF_X2 U31 ( .A(DATAIN[30]), .Z(n395) );
  BUF_X1 U32 ( .A(n1146), .Z(n13) );
  BUF_X1 U33 ( .A(n1146), .Z(n3604) );
  BUF_X2 U34 ( .A(DATAIN[0]), .Z(n387) );
  INV_X1 U35 ( .A(n3594), .ZN(n14) );
  CLKBUF_X3 U36 ( .A(DATAIN[21]), .Z(n880) );
  BUF_X1 U37 ( .A(n1355), .Z(n3549) );
  INV_X1 U38 ( .A(n897), .ZN(n15) );
  INV_X1 U39 ( .A(n3639), .ZN(n16) );
  BUF_X1 U40 ( .A(DATAIN[29]), .Z(n865) );
  BUF_X1 U41 ( .A(n3550), .Z(n17) );
  BUF_X1 U42 ( .A(n1355), .Z(n3547) );
  BUF_X2 U43 ( .A(DATAIN[18]), .Z(n885) );
  BUF_X1 U44 ( .A(DATAIN[3]), .Z(n791) );
  INV_X1 U45 ( .A(n209), .ZN(n18) );
  BUF_X1 U46 ( .A(DATAIN[22]), .Z(n19) );
  BUF_X1 U47 ( .A(net39096), .Z(n20) );
  INV_X1 U48 ( .A(n165), .ZN(n21) );
  INV_X1 U49 ( .A(n791), .ZN(n22) );
  BUF_X1 U50 ( .A(DATAIN[3]), .Z(n249) );
  BUF_X1 U51 ( .A(ADD_WR[0]), .Z(n393) );
  BUF_X1 U52 ( .A(n1355), .Z(n3548) );
  INV_X1 U53 ( .A(n558), .ZN(n23) );
  INV_X1 U54 ( .A(n558), .ZN(n24) );
  BUF_X1 U55 ( .A(DATAIN[20]), .Z(n882) );
  INV_X1 U56 ( .A(n248), .ZN(n25) );
  BUF_X1 U57 ( .A(DATAIN[31]), .Z(n785) );
  INV_X1 U58 ( .A(n883), .ZN(n26) );
  BUF_X1 U59 ( .A(DATAIN[7]), .Z(n793) );
  BUF_X1 U60 ( .A(DATAIN[4]), .Z(n163) );
  INV_X1 U61 ( .A(n412), .ZN(n27) );
  INV_X1 U62 ( .A(n199), .ZN(n28) );
  INV_X1 U63 ( .A(n868), .ZN(n29) );
  BUF_X1 U64 ( .A(n1388), .Z(n3540) );
  BUF_X1 U65 ( .A(n1388), .Z(n3542) );
  BUF_X1 U66 ( .A(n590), .Z(n3529) );
  BUF_X1 U67 ( .A(n590), .Z(n3531) );
  BUF_X2 U68 ( .A(n1317), .Z(n3565) );
  BUF_X2 U69 ( .A(n1284), .Z(n3572) );
  BUF_X1 U70 ( .A(n1284), .Z(n3575) );
  BUF_X1 U71 ( .A(n3317), .Z(n3620) );
  BUF_X2 U72 ( .A(n1180), .Z(n3592) );
  BUF_X1 U73 ( .A(DATAIN[12]), .Z(n897) );
  BUF_X1 U74 ( .A(n1284), .Z(n3574) );
  BUF_X1 U75 ( .A(ADD_WR[1]), .Z(n726) );
  AND2_X1 U76 ( .A1(n1106), .A2(n1247), .ZN(n175) );
  INV_X1 U77 ( .A(net26597), .ZN(n32) );
  BUF_X1 U78 ( .A(DATAIN[20]), .Z(n161) );
  BUF_X1 U79 ( .A(DATAIN[7]), .Z(n162) );
  BUF_X1 U80 ( .A(DATAIN[4]), .Z(n789) );
  BUF_X2 U81 ( .A(DATAIN[24]), .Z(n874) );
  AND2_X2 U82 ( .A1(n1247), .A2(n1072), .ZN(n247) );
  INV_X1 U83 ( .A(n219), .ZN(n164) );
  BUF_X1 U84 ( .A(DATAIN[12]), .Z(n165) );
  BUF_X1 U85 ( .A(DATAIN[12]), .Z(n166) );
  BUF_X1 U86 ( .A(DATAIN[12]), .Z(n898) );
  BUF_X1 U87 ( .A(DATAIN[3]), .Z(n167) );
  NOR2_X1 U88 ( .A1(n4241), .A2(ADD_RD2[2]), .ZN(n2160) );
  AND2_X1 U89 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n2164) );
  NOR2_X1 U90 ( .A1(n4238), .A2(ADD_RD1[2]), .ZN(n2751) );
  AND2_X1 U91 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n2755) );
  AND2_X1 U92 ( .A1(ADD_RD2[2]), .A2(n4241), .ZN(n2165) );
  AND2_X1 U93 ( .A1(ADD_RD1[2]), .A2(n4238), .ZN(n2756) );
  BUF_X1 U94 ( .A(n1146), .Z(n597) );
  BUF_X1 U95 ( .A(n1317), .Z(n3567) );
  BUF_X1 U96 ( .A(n1355), .Z(n3550) );
  BUF_X1 U97 ( .A(DATAIN[3]), .Z(n790) );
  BUF_X1 U98 ( .A(DATAIN[6]), .Z(n794) );
  BUF_X1 U99 ( .A(DATAIN[14]), .Z(n893) );
  BUF_X1 U100 ( .A(DATAIN[19]), .Z(n884) );
  BUF_X1 U101 ( .A(DATAIN[20]), .Z(n881) );
  BUF_X1 U102 ( .A(DATAIN[7]), .Z(n792) );
  BUF_X1 U103 ( .A(DATAIN[22]), .Z(n878) );
  BUF_X1 U104 ( .A(n3577), .Z(n205) );
  BUF_X1 U105 ( .A(n3579), .Z(n3577) );
  BUF_X1 U106 ( .A(n174), .Z(n3630) );
  BUF_X1 U107 ( .A(DATAIN[17]), .Z(n887) );
  INV_X1 U108 ( .A(n1282), .ZN(n3579) );
  BUF_X1 U109 ( .A(n1074), .Z(n3638) );
  INV_X1 U110 ( .A(n3591), .ZN(n168) );
  BUF_X1 U111 ( .A(n1180), .Z(n3591) );
  BUF_X1 U112 ( .A(n3604), .Z(n234) );
  AND2_X1 U113 ( .A1(n1072), .A2(n1070), .ZN(n169) );
  INV_X1 U114 ( .A(n3594), .ZN(n3589) );
  INV_X1 U115 ( .A(n900), .ZN(n170) );
  BUF_X1 U116 ( .A(DATAIN[2]), .Z(n189) );
  INV_X1 U117 ( .A(n3594), .ZN(n171) );
  INV_X1 U118 ( .A(n3594), .ZN(n3588) );
  BUF_X1 U119 ( .A(n3555), .Z(n3554) );
  BUF_X1 U120 ( .A(n3555), .Z(n3552) );
  BUF_X1 U121 ( .A(n3555), .Z(n3551) );
  BUF_X2 U122 ( .A(n1074), .Z(n3636) );
  BUF_X1 U123 ( .A(n576), .Z(n3522) );
  BUF_X1 U124 ( .A(n576), .Z(n3526) );
  BUF_X1 U125 ( .A(n576), .Z(n3525) );
  INV_X1 U126 ( .A(n784), .ZN(n172) );
  INV_X1 U127 ( .A(n3316), .ZN(n173) );
  BUF_X1 U128 ( .A(DATAIN[11]), .Z(n549) );
  BUF_X1 U129 ( .A(DATAIN[2]), .Z(n190) );
  NAND2_X1 U130 ( .A1(n414), .A2(n1070), .ZN(n174) );
  INV_X1 U131 ( .A(n1556), .ZN(n176) );
  INV_X1 U132 ( .A(n895), .ZN(n177) );
  INV_X1 U133 ( .A(n798), .ZN(n178) );
  INV_X1 U134 ( .A(n779), .ZN(n179) );
  INV_X1 U135 ( .A(n891), .ZN(n180) );
  INV_X1 U136 ( .A(n897), .ZN(n181) );
  BUF_X1 U137 ( .A(DATAIN[11]), .Z(n548) );
  INV_X1 U138 ( .A(n878), .ZN(n182) );
  INV_X1 U139 ( .A(n878), .ZN(n183) );
  INV_X1 U140 ( .A(n872), .ZN(n184) );
  INV_X1 U141 ( .A(n879), .ZN(n185) );
  INV_X1 U142 ( .A(n879), .ZN(n186) );
  BUF_X2 U143 ( .A(DATAIN[21]), .Z(n879) );
  AND2_X1 U144 ( .A1(n1247), .A2(n1178), .ZN(n187) );
  BUF_X1 U145 ( .A(n187), .Z(n3560) );
  BUF_X1 U146 ( .A(DATAIN[19]), .Z(n545) );
  INV_X1 U147 ( .A(n209), .ZN(n188) );
  BUF_X1 U148 ( .A(DATAIN[2]), .Z(n900) );
  BUF_X1 U149 ( .A(n3504), .Z(n3503) );
  BUF_X1 U150 ( .A(n3504), .Z(n3502) );
  INV_X1 U151 ( .A(n901), .ZN(n191) );
  BUF_X1 U152 ( .A(n3604), .Z(n3603) );
  BUF_X1 U153 ( .A(n3604), .Z(n3602) );
  BUF_X2 U154 ( .A(n1047), .Z(n192) );
  INV_X1 U155 ( .A(n788), .ZN(n193) );
  INV_X1 U156 ( .A(n899), .ZN(n194) );
  BUF_X1 U157 ( .A(DATAIN[17]), .Z(n250) );
  BUF_X1 U158 ( .A(n174), .Z(n3628) );
  BUF_X1 U159 ( .A(n174), .Z(n3629) );
  INV_X1 U160 ( .A(n797), .ZN(n195) );
  INV_X1 U161 ( .A(n215), .ZN(n196) );
  INV_X1 U162 ( .A(net28528), .ZN(n197) );
  CLKBUF_X2 U163 ( .A(DATAIN[10]), .Z(n283) );
  BUF_X2 U164 ( .A(n1423), .Z(n3527) );
  BUF_X1 U165 ( .A(DATAIN[17]), .Z(n888) );
  INV_X1 U166 ( .A(n903), .ZN(n198) );
  INV_X1 U167 ( .A(n1556), .ZN(n3504) );
  BUF_X1 U168 ( .A(DATAIN[5]), .Z(n786) );
  BUF_X1 U169 ( .A(DATAIN[11]), .Z(n797) );
  BUF_X1 U170 ( .A(DATAIN[27]), .Z(n867) );
  BUF_X1 U171 ( .A(DATAIN[26]), .Z(n869) );
  BUF_X1 U172 ( .A(DATAIN[25]), .Z(n199) );
  BUF_X1 U173 ( .A(DATAIN[25]), .Z(n200) );
  BUF_X1 U174 ( .A(DATAIN[25]), .Z(n872) );
  INV_X1 U175 ( .A(n781), .ZN(n201) );
  INV_X1 U176 ( .A(DATAIN[8]), .ZN(n4263) );
  BUF_X1 U177 ( .A(DATAIN[21]), .Z(n242) );
  INV_X1 U178 ( .A(n788), .ZN(n4267) );
  INV_X1 U179 ( .A(n899), .ZN(n4269) );
  BUF_X1 U180 ( .A(n1068), .Z(n202) );
  INV_X1 U181 ( .A(n3543), .ZN(n203) );
  INV_X1 U182 ( .A(n3543), .ZN(n204) );
  BUF_X1 U183 ( .A(DATAIN[16]), .Z(n889) );
  INV_X1 U184 ( .A(n163), .ZN(n275) );
  INV_X1 U185 ( .A(n899), .ZN(n268) );
  INV_X1 U186 ( .A(n784), .ZN(n4243) );
  BUF_X1 U187 ( .A(n576), .Z(n3521) );
  BUF_X1 U188 ( .A(n576), .Z(n3524) );
  INV_X1 U189 ( .A(n3587), .ZN(n206) );
  BUF_X1 U190 ( .A(DATAIN[20]), .Z(n207) );
  INV_X1 U191 ( .A(n881), .ZN(n208) );
  BUF_X1 U192 ( .A(DATAIN[15]), .Z(n209) );
  BUF_X1 U193 ( .A(DATAIN[15]), .Z(n210) );
  BUF_X1 U194 ( .A(DATAIN[15]), .Z(n892) );
  BUF_X1 U195 ( .A(DATAIN[7]), .Z(n211) );
  INV_X1 U196 ( .A(n162), .ZN(n212) );
  INV_X1 U197 ( .A(n3511), .ZN(n213) );
  INV_X1 U198 ( .A(n3511), .ZN(n214) );
  BUF_X1 U199 ( .A(n1489), .Z(n3508) );
  BUF_X1 U200 ( .A(n1489), .Z(n3509) );
  BUF_X1 U201 ( .A(n1489), .Z(n3510) );
  BUF_X1 U202 ( .A(DATAIN[2]), .Z(n899) );
  BUF_X1 U203 ( .A(DATAIN[4]), .Z(n788) );
  BUF_X1 U204 ( .A(n3547), .Z(n215) );
  BUF_X1 U205 ( .A(n3547), .Z(n216) );
  BUF_X1 U206 ( .A(n3547), .Z(n217) );
  BUF_X1 U207 ( .A(n3547), .Z(n218) );
  BUF_X1 U208 ( .A(n3548), .Z(n219) );
  BUF_X1 U209 ( .A(n3549), .Z(n220) );
  CLKBUF_X1 U210 ( .A(DATAIN[0]), .Z(n904) );
  CLKBUF_X1 U211 ( .A(DATAIN[0]), .Z(n388) );
  INV_X1 U212 ( .A(n800), .ZN(n221) );
  INV_X1 U213 ( .A(n3517), .ZN(n3512) );
  BUF_X2 U214 ( .A(n3317), .Z(n3622) );
  BUF_X1 U215 ( .A(net39096), .Z(net44604) );
  INV_X1 U216 ( .A(n889), .ZN(n727) );
  BUF_X1 U217 ( .A(n1068), .Z(n222) );
  BUF_X1 U218 ( .A(n1523), .Z(net26589) );
  BUF_X1 U219 ( .A(n3301), .Z(n3534) );
  CLKBUF_X3 U220 ( .A(DATAIN[14]), .Z(n223) );
  INV_X1 U221 ( .A(n875), .ZN(n224) );
  BUF_X2 U222 ( .A(DATAIN[23]), .Z(n875) );
  AND2_X1 U223 ( .A1(n1144), .A2(n1070), .ZN(n783) );
  INV_X1 U224 ( .A(n900), .ZN(n225) );
  INV_X1 U225 ( .A(n899), .ZN(n733) );
  BUF_X1 U226 ( .A(n1074), .Z(n3637) );
  INV_X1 U227 ( .A(n887), .ZN(n739) );
  CLKBUF_X1 U228 ( .A(n874), .Z(n397) );
  OAI22_X1 U229 ( .A1(n280), .A2(n3593), .B1(n3590), .B2(n227), .ZN(n226) );
  BUF_X1 U230 ( .A(n1523), .Z(net26585) );
  BUF_X1 U231 ( .A(net39096), .Z(net26249) );
  BUF_X1 U232 ( .A(n1249), .Z(net38912) );
  INV_X1 U233 ( .A(net26597), .ZN(n228) );
  INV_X1 U234 ( .A(net26593), .ZN(n229) );
  BUF_X1 U235 ( .A(DATAIN[29]), .Z(n230) );
  BUF_X1 U236 ( .A(DATAIN[29]), .Z(n231) );
  BUF_X1 U237 ( .A(DATAIN[29]), .Z(n866) );
  INV_X1 U238 ( .A(n266), .ZN(n232) );
  INV_X1 U239 ( .A(n266), .ZN(n233) );
  BUF_X1 U240 ( .A(n597), .Z(n3599) );
  INV_X1 U241 ( .A(n793), .ZN(n235) );
  OAI22_X1 U242 ( .A1(n705), .A2(n3630), .B1(n768), .B2(n237), .ZN(n236) );
  CLKBUF_X1 U243 ( .A(n174), .Z(n3626) );
  INV_X1 U244 ( .A(n790), .ZN(n238) );
  INV_X1 U245 ( .A(n790), .ZN(n239) );
  INV_X1 U246 ( .A(n267), .ZN(n240) );
  INV_X1 U247 ( .A(n788), .ZN(n731) );
  INV_X1 U248 ( .A(n873), .ZN(n4249) );
  CLKBUF_X1 U249 ( .A(DATAIN[24]), .Z(n873) );
  INV_X1 U250 ( .A(n790), .ZN(n4268) );
  BUF_X1 U251 ( .A(net39096), .Z(n241) );
  INV_X1 U252 ( .A(n3574), .ZN(n243) );
  INV_X1 U253 ( .A(n3573), .ZN(n244) );
  BUF_X1 U254 ( .A(n1249), .Z(net44605) );
  BUF_X1 U255 ( .A(n1249), .Z(net44860) );
  BUF_X1 U256 ( .A(n596), .Z(n3498) );
  BUF_X1 U257 ( .A(n596), .Z(n3495) );
  BUF_X1 U258 ( .A(n596), .Z(n3499) );
  BUF_X1 U259 ( .A(n596), .Z(n3497) );
  BUF_X1 U260 ( .A(n596), .Z(n3496) );
  BUF_X1 U261 ( .A(n596), .Z(n3500) );
  BUF_X1 U262 ( .A(DATAIN[22]), .Z(n245) );
  CLKBUF_X3 U263 ( .A(DATAIN[28]), .Z(n246) );
  BUF_X2 U264 ( .A(DATAIN[28]), .Z(net28528) );
  AOI22_X1 U265 ( .A1(net28529), .A2(net44303), .B1(net44860), .B2(
        \registers[22][28] ), .ZN(n1277) );
  INV_X1 U266 ( .A(n1277), .ZN(net18066) );
  INV_X1 U267 ( .A(n247), .ZN(n1249) );
  INV_X1 U268 ( .A(n1249), .ZN(net26245) );
  INV_X1 U269 ( .A(n248), .ZN(net26243) );
  INV_X1 U270 ( .A(n247), .ZN(n248) );
  INV_X1 U271 ( .A(n248), .ZN(net44303) );
  INV_X1 U272 ( .A(n248), .ZN(net26247) );
  INV_X1 U273 ( .A(n248), .ZN(net44304) );
  CLKBUF_X3 U274 ( .A(DATAIN[28]), .Z(net28529) );
  AOI22_X1 U275 ( .A1(net26747), .A2(\registers[23][28] ), .B1(net26753), .B2(
        \registers[22][28] ), .ZN(n1683) );
  AOI22_X1 U276 ( .A1(net26933), .A2(\registers[23][28] ), .B1(net26939), .B2(
        \registers[22][28] ), .ZN(n2274) );
  INV_X1 U277 ( .A(n247), .ZN(net39096) );
  AND2_X2 U278 ( .A1(n1072), .A2(n1352), .ZN(net33812) );
  NAND2_X1 U279 ( .A1(n1521), .A2(n1072), .ZN(n1523) );
  BUF_X1 U280 ( .A(n874), .Z(n398) );
  OAI22_X1 U281 ( .A1(n741), .A2(net44860), .B1(net26245), .B2(n252), .ZN(n251) );
  OAI22_X1 U282 ( .A1(n183), .A2(net44605), .B1(net26245), .B2(n254), .ZN(n253) );
  OAI22_X1 U283 ( .A1(n709), .A2(n3592), .B1(n171), .B2(n256), .ZN(n255) );
  OAI22_X1 U284 ( .A1(n269), .A2(n3527), .B1(n680), .B2(n258), .ZN(n257) );
  BUF_X1 U285 ( .A(n576), .Z(n3523) );
  CLKBUF_X3 U286 ( .A(DATAIN[18]), .Z(n259) );
  INV_X1 U287 ( .A(n884), .ZN(n260) );
  INV_X1 U288 ( .A(n884), .ZN(n745) );
  BUF_X1 U289 ( .A(DATAIN[16]), .Z(n261) );
  BUF_X1 U290 ( .A(DATAIN[16]), .Z(n262) );
  BUF_X1 U291 ( .A(DATAIN[16]), .Z(n890) );
  BUF_X1 U292 ( .A(n1215), .Z(n3584) );
  BUF_X1 U293 ( .A(n1215), .Z(n3586) );
  BUF_X1 U294 ( .A(n1215), .Z(n3585) );
  INV_X1 U295 ( .A(n893), .ZN(n4257) );
  INV_X1 U296 ( .A(n893), .ZN(n269) );
  INV_X1 U297 ( .A(net28528), .ZN(net17879) );
  INV_X1 U298 ( .A(net28528), .ZN(net44818) );
  INV_X1 U299 ( .A(n784), .ZN(n263) );
  INV_X1 U300 ( .A(n784), .ZN(n605) );
  BUF_X1 U301 ( .A(DATAIN[23]), .Z(n264) );
  BUF_X1 U302 ( .A(DATAIN[23]), .Z(n265) );
  BUF_X1 U303 ( .A(DATAIN[23]), .Z(n876) );
  BUF_X1 U304 ( .A(n1351), .Z(n266) );
  BUF_X1 U305 ( .A(DATAIN[4]), .Z(n267) );
  INV_X1 U306 ( .A(DATAIN[30]), .ZN(n270) );
  INV_X1 U307 ( .A(DATAIN[30]), .ZN(n4244) );
  INV_X1 U308 ( .A(n865), .ZN(n271) );
  OAI22_X1 U309 ( .A1(n280), .A2(n3637), .B1(n3633), .B2(n273), .ZN(n272) );
  INV_X1 U310 ( .A(n166), .ZN(n274) );
  INV_X1 U311 ( .A(n3517), .ZN(n276) );
  INV_X1 U312 ( .A(n3517), .ZN(n277) );
  CLKBUF_X3 U313 ( .A(DATAIN[6]), .Z(n278) );
  BUF_X1 U314 ( .A(n1523), .Z(net26595) );
  BUF_X1 U315 ( .A(n1074), .Z(n3635) );
  CLKBUF_X3 U316 ( .A(DATAIN[1]), .Z(n279) );
  INV_X1 U317 ( .A(n873), .ZN(n280) );
  INV_X1 U318 ( .A(n786), .ZN(n4266) );
  INV_X1 U319 ( .A(n892), .ZN(n281) );
  CLKBUF_X3 U320 ( .A(DATAIN[9]), .Z(n282) );
  CLKBUF_X3 U321 ( .A(DATAIN[13]), .Z(n284) );
  INV_X1 U322 ( .A(n1555), .ZN(n285) );
  INV_X1 U323 ( .A(n1555), .ZN(n286) );
  INV_X1 U324 ( .A(n1555), .ZN(n287) );
  INV_X1 U325 ( .A(n287), .ZN(n288) );
  INV_X1 U326 ( .A(n287), .ZN(n353) );
  INV_X1 U327 ( .A(n287), .ZN(n354) );
  INV_X1 U328 ( .A(n285), .ZN(n355) );
  INV_X1 U329 ( .A(n285), .ZN(n356) );
  INV_X1 U330 ( .A(n355), .ZN(n357) );
  INV_X1 U331 ( .A(n355), .ZN(n358) );
  INV_X1 U332 ( .A(n355), .ZN(n359) );
  INV_X1 U333 ( .A(n356), .ZN(n360) );
  INV_X1 U334 ( .A(n356), .ZN(n361) );
  INV_X1 U335 ( .A(n356), .ZN(n362) );
  INV_X1 U336 ( .A(n286), .ZN(n363) );
  INV_X1 U337 ( .A(n286), .ZN(n364) );
  INV_X1 U338 ( .A(n363), .ZN(n365) );
  INV_X1 U339 ( .A(n363), .ZN(n366) );
  INV_X1 U340 ( .A(n364), .ZN(n367) );
  INV_X1 U341 ( .A(n364), .ZN(n368) );
  INV_X1 U342 ( .A(n364), .ZN(n369) );
  INV_X1 U343 ( .A(n175), .ZN(n370) );
  INV_X1 U344 ( .A(n175), .ZN(n371) );
  INV_X1 U345 ( .A(n175), .ZN(n372) );
  INV_X1 U346 ( .A(n175), .ZN(n373) );
  INV_X1 U347 ( .A(n373), .ZN(n374) );
  INV_X1 U348 ( .A(n373), .ZN(n375) );
  INV_X1 U349 ( .A(n373), .ZN(n376) );
  INV_X1 U350 ( .A(n373), .ZN(n377) );
  INV_X1 U351 ( .A(n379), .ZN(n378) );
  INV_X1 U352 ( .A(n175), .ZN(n379) );
  INV_X1 U353 ( .A(n379), .ZN(n380) );
  INV_X1 U354 ( .A(n373), .ZN(n381) );
  INV_X1 U355 ( .A(n379), .ZN(n382) );
  INV_X1 U356 ( .A(n379), .ZN(n383) );
  INV_X1 U357 ( .A(n379), .ZN(n384) );
  OAI22_X1 U358 ( .A1(n415), .A2(n3514), .B1(n389), .B2(n386), .ZN(n385) );
  CLKBUF_X3 U359 ( .A(DATAIN[18]), .Z(n886) );
  CLKBUF_X1 U360 ( .A(n1456), .Z(n3514) );
  BUF_X2 U361 ( .A(n1456), .Z(n3516) );
  INV_X1 U362 ( .A(n3517), .ZN(n3513) );
  BUF_X1 U363 ( .A(n1284), .Z(n3573) );
  INV_X1 U364 ( .A(n3517), .ZN(n389) );
  INV_X1 U365 ( .A(n3517), .ZN(n390) );
  OAI22_X1 U366 ( .A1(n401), .A2(n217), .B1(n164), .B2(n392), .ZN(n391) );
  INV_X1 U367 ( .A(n865), .ZN(n742) );
  INV_X1 U368 ( .A(DATAIN[29]), .ZN(n743) );
  BUF_X1 U369 ( .A(net39096), .Z(net44322) );
  INV_X1 U370 ( .A(n161), .ZN(n396) );
  INV_X1 U371 ( .A(n395), .ZN(n399) );
  INV_X1 U372 ( .A(n791), .ZN(n400) );
  INV_X1 U373 ( .A(n249), .ZN(n732) );
  INV_X1 U374 ( .A(n891), .ZN(n401) );
  INV_X1 U375 ( .A(n887), .ZN(n402) );
  INV_X1 U376 ( .A(n887), .ZN(n403) );
  INV_X1 U377 ( .A(n887), .ZN(n4255) );
  OAI22_X1 U378 ( .A1(n6), .A2(net44322), .B1(net26243), .B2(n405), .ZN(n404)
         );
  OAI22_X1 U379 ( .A1(n18), .A2(net26595), .B1(n407), .B2(net39089), .ZN(n406)
         );
  BUF_X1 U380 ( .A(DATAIN[25]), .Z(n871) );
  INV_X1 U381 ( .A(n3549), .ZN(n408) );
  BUF_X1 U382 ( .A(n874), .Z(n409) );
  BUF_X1 U383 ( .A(DATAIN[5]), .Z(n412) );
  BUF_X1 U384 ( .A(DATAIN[5]), .Z(n413) );
  BUF_X1 U385 ( .A(DATAIN[5]), .Z(n787) );
  INV_X1 U386 ( .A(net33812), .ZN(net44473) );
  INV_X1 U387 ( .A(net33812), .ZN(net44474) );
  AND3_X1 U388 ( .A1(n681), .A2(n551), .A3(n710), .ZN(n414) );
  INV_X1 U389 ( .A(n885), .ZN(n415) );
  INV_X1 U390 ( .A(n885), .ZN(n4254) );
  BUF_X1 U391 ( .A(DATAIN[15]), .Z(n891) );
  BUF_X1 U392 ( .A(n1074), .Z(n3639) );
  CLKBUF_X1 U393 ( .A(DATAIN[19]), .Z(n416) );
  INV_X1 U394 ( .A(n794), .ZN(n546) );
  INV_X1 U395 ( .A(n794), .ZN(n547) );
  INV_X1 U396 ( .A(n794), .ZN(n4265) );
  BUF_X2 U397 ( .A(DATAIN[31]), .Z(n550) );
  CLKBUF_X1 U398 ( .A(ADD_WR[2]), .Z(n551) );
  INV_X1 U399 ( .A(n889), .ZN(n552) );
  INV_X1 U400 ( .A(n889), .ZN(n553) );
  INV_X1 U401 ( .A(n889), .ZN(n4256) );
  BUF_X1 U402 ( .A(n187), .Z(n3559) );
  BUF_X1 U403 ( .A(n187), .Z(n3561) );
  INV_X1 U404 ( .A(n786), .ZN(n554) );
  INV_X1 U405 ( .A(n786), .ZN(n555) );
  INV_X1 U406 ( .A(n786), .ZN(n738) );
  BUF_X1 U407 ( .A(DATAIN[27]), .Z(n556) );
  BUF_X1 U408 ( .A(DATAIN[27]), .Z(n557) );
  BUF_X1 U409 ( .A(DATAIN[27]), .Z(n868) );
  BUF_X1 U410 ( .A(DATAIN[26]), .Z(n558) );
  BUF_X1 U411 ( .A(DATAIN[26]), .Z(n559) );
  BUF_X1 U412 ( .A(DATAIN[26]), .Z(n870) );
  BUF_X1 U413 ( .A(DATAIN[22]), .Z(n877) );
  INV_X1 U414 ( .A(n884), .ZN(n560) );
  INV_X1 U415 ( .A(n884), .ZN(n4253) );
  INV_X1 U416 ( .A(n3622), .ZN(n561) );
  INV_X1 U417 ( .A(n3622), .ZN(n562) );
  INV_X1 U418 ( .A(n1558), .ZN(n563) );
  INV_X1 U419 ( .A(n1558), .ZN(n564) );
  INV_X2 U420 ( .A(n564), .ZN(n565) );
  INV_X2 U421 ( .A(n564), .ZN(n566) );
  INV_X1 U422 ( .A(n563), .ZN(n567) );
  INV_X1 U423 ( .A(n567), .ZN(n568) );
  INV_X1 U424 ( .A(n567), .ZN(n569) );
  INV_X1 U425 ( .A(n567), .ZN(n570) );
  INV_X1 U426 ( .A(n1558), .ZN(n571) );
  INV_X1 U427 ( .A(n567), .ZN(n572) );
  INV_X1 U428 ( .A(n567), .ZN(n573) );
  INV_X1 U429 ( .A(n797), .ZN(n574) );
  INV_X1 U430 ( .A(n797), .ZN(n575) );
  INV_X1 U431 ( .A(n797), .ZN(n4260) );
  BUF_X1 U432 ( .A(DATAIN[11]), .Z(n796) );
  BUF_X1 U433 ( .A(n1423), .Z(n576) );
  BUF_X1 U434 ( .A(n174), .Z(n3627) );
  INV_X1 U435 ( .A(n3575), .ZN(n577) );
  INV_X1 U436 ( .A(n865), .ZN(n4245) );
  INV_X1 U437 ( .A(n1557), .ZN(n578) );
  INV_X1 U438 ( .A(n1557), .ZN(n579) );
  INV_X2 U439 ( .A(n579), .ZN(n580) );
  INV_X2 U440 ( .A(n579), .ZN(n581) );
  INV_X1 U441 ( .A(n578), .ZN(n582) );
  INV_X1 U442 ( .A(n582), .ZN(n583) );
  INV_X1 U443 ( .A(n582), .ZN(n584) );
  INV_X1 U444 ( .A(n582), .ZN(n585) );
  INV_X1 U445 ( .A(n578), .ZN(n586) );
  INV_X1 U446 ( .A(n586), .ZN(n587) );
  INV_X1 U447 ( .A(n586), .ZN(n588) );
  INV_X1 U448 ( .A(n586), .ZN(n589) );
  AND2_X1 U449 ( .A1(n1144), .A2(n1352), .ZN(n590) );
  INV_X1 U450 ( .A(n869), .ZN(n591) );
  INV_X1 U451 ( .A(n869), .ZN(n592) );
  INV_X1 U452 ( .A(n869), .ZN(n4247) );
  INV_X1 U453 ( .A(n867), .ZN(n593) );
  INV_X1 U454 ( .A(n867), .ZN(n594) );
  INV_X1 U455 ( .A(n867), .ZN(n4246) );
  INV_X1 U456 ( .A(n3567), .ZN(n595) );
  BUF_X1 U457 ( .A(DATAIN[31]), .Z(n784) );
  BUF_X1 U458 ( .A(n1523), .Z(net26591) );
  BUF_X1 U459 ( .A(n1523), .Z(net26593) );
  BUF_X1 U460 ( .A(n1523), .Z(net26597) );
  BUF_X1 U461 ( .A(n1560), .Z(n596) );
  INV_X1 U462 ( .A(n895), .ZN(n598) );
  INV_X1 U463 ( .A(n895), .ZN(n599) );
  INV_X1 U464 ( .A(n895), .ZN(n4258) );
  BUF_X2 U465 ( .A(DATAIN[13]), .Z(n895) );
  INV_X1 U466 ( .A(n779), .ZN(n600) );
  INV_X1 U467 ( .A(n779), .ZN(n601) );
  INV_X1 U468 ( .A(n779), .ZN(n4262) );
  BUF_X2 U469 ( .A(DATAIN[9]), .Z(n779) );
  INV_X1 U470 ( .A(n891), .ZN(n729) );
  INV_X1 U471 ( .A(n165), .ZN(n4259) );
  INV_X1 U472 ( .A(n897), .ZN(n740) );
  INV_X1 U473 ( .A(n891), .ZN(n728) );
  INV_X1 U474 ( .A(net26593), .ZN(net39089) );
  INV_X1 U475 ( .A(net26591), .ZN(net39090) );
  INV_X1 U476 ( .A(n885), .ZN(n602) );
  INV_X1 U477 ( .A(n3594), .ZN(n603) );
  INV_X1 U478 ( .A(n549), .ZN(n604) );
  INV_X1 U479 ( .A(n903), .ZN(n606) );
  INV_X1 U480 ( .A(n903), .ZN(n607) );
  INV_X1 U481 ( .A(n903), .ZN(n4271) );
  BUF_X2 U482 ( .A(DATAIN[0]), .Z(n903) );
  INV_X1 U483 ( .A(net28528), .ZN(net39055) );
  INV_X1 U484 ( .A(n901), .ZN(n608) );
  INV_X1 U485 ( .A(n901), .ZN(n673) );
  INV_X1 U486 ( .A(n901), .ZN(n4270) );
  BUF_X2 U487 ( .A(DATAIN[1]), .Z(n901) );
  INV_X1 U488 ( .A(n798), .ZN(n674) );
  INV_X1 U489 ( .A(n798), .ZN(n675) );
  INV_X1 U490 ( .A(n798), .ZN(n4261) );
  BUF_X2 U491 ( .A(DATAIN[10]), .Z(n798) );
  NOR3_X1 U492 ( .A1(n710), .A2(n4234), .A3(n681), .ZN(n676) );
  NOR3_X1 U493 ( .A1(n710), .A2(n4234), .A3(n681), .ZN(n1069) );
  INV_X1 U494 ( .A(n3501), .ZN(n677) );
  INV_X1 U495 ( .A(n3501), .ZN(n678) );
  INV_X1 U496 ( .A(n3527), .ZN(n679) );
  INV_X1 U497 ( .A(n3527), .ZN(n680) );
  INV_X1 U498 ( .A(net26591), .ZN(net38992) );
  INV_X1 U499 ( .A(net26593), .ZN(net38993) );
  INV_X1 U500 ( .A(n169), .ZN(net38964) );
  INV_X1 U501 ( .A(n169), .ZN(net38965) );
  INV_X1 U502 ( .A(n169), .ZN(net38966) );
  INV_X1 U503 ( .A(n169), .ZN(net38967) );
  INV_X1 U504 ( .A(net38967), .ZN(net38968) );
  INV_X1 U505 ( .A(net38967), .ZN(net38969) );
  INV_X1 U506 ( .A(net38967), .ZN(net38970) );
  INV_X1 U507 ( .A(n169), .ZN(net38971) );
  INV_X1 U508 ( .A(net38971), .ZN(net38972) );
  INV_X1 U509 ( .A(net38971), .ZN(net38973) );
  INV_X1 U510 ( .A(net38971), .ZN(net38974) );
  AND3_X1 U511 ( .A1(ADD_WR[3]), .A2(n1213), .A3(ADD_WR[4]), .ZN(n1070) );
  INV_X1 U512 ( .A(ADD_WR[1]), .ZN(n681) );
  INV_X1 U513 ( .A(n3511), .ZN(n682) );
  INV_X1 U514 ( .A(n3511), .ZN(n683) );
  INV_X1 U515 ( .A(n3587), .ZN(n684) );
  OAI22_X1 U516 ( .A1(n4), .A2(n3585), .B1(n765), .B2(n686), .ZN(n685) );
  INV_X1 U517 ( .A(n3550), .ZN(n687) );
  INV_X1 U518 ( .A(n3631), .ZN(n688) );
  INV_X1 U519 ( .A(n3631), .ZN(n689) );
  INV_X1 U520 ( .A(n3639), .ZN(n690) );
  INV_X1 U521 ( .A(n3635), .ZN(n691) );
  INV_X1 U522 ( .A(n3543), .ZN(n692) );
  INV_X1 U523 ( .A(n3543), .ZN(n693) );
  OAI22_X1 U524 ( .A1(n15), .A2(n3542), .B1(n203), .B2(n695), .ZN(n694) );
  INV_X1 U525 ( .A(n897), .ZN(n741) );
  AND3_X1 U526 ( .A1(n681), .A2(n551), .A3(n710), .ZN(n1140) );
  INV_X1 U527 ( .A(ADD_WR[1]), .ZN(n4235) );
  INV_X1 U528 ( .A(DATAIN[14]), .ZN(n696) );
  INV_X1 U529 ( .A(n875), .ZN(n697) );
  INV_X1 U530 ( .A(n875), .ZN(n698) );
  INV_X1 U532 ( .A(n875), .ZN(n4250) );
  INV_X1 U533 ( .A(n19), .ZN(n699) );
  INV_X1 U534 ( .A(n877), .ZN(n700) );
  INV_X1 U535 ( .A(n878), .ZN(n4251) );
  INV_X1 U536 ( .A(n881), .ZN(n701) );
  INV_X1 U537 ( .A(n881), .ZN(n702) );
  INV_X1 U538 ( .A(n882), .ZN(n4252) );
  CLKBUF_X3 U539 ( .A(DATAIN[14]), .Z(n894) );
  INV_X1 U540 ( .A(n549), .ZN(n703) );
  CLKBUF_X3 U541 ( .A(DATAIN[10]), .Z(n799) );
  INV_X1 U542 ( .A(n792), .ZN(n704) );
  INV_X1 U543 ( .A(n792), .ZN(n705) );
  INV_X1 U544 ( .A(n792), .ZN(n4264) );
  CLKBUF_X3 U545 ( .A(DATAIN[6]), .Z(n795) );
  INV_X1 U546 ( .A(n871), .ZN(n706) );
  INV_X1 U547 ( .A(n871), .ZN(n707) );
  INV_X1 U548 ( .A(n871), .ZN(n4248) );
  INV_X1 U549 ( .A(n879), .ZN(n708) );
  INV_X1 U550 ( .A(n879), .ZN(n709) );
  BUF_X2 U551 ( .A(n1456), .Z(n3517) );
  INV_X1 U552 ( .A(ADD_WR[0]), .ZN(n710) );
  BUF_X1 U553 ( .A(n1212), .Z(n711) );
  INV_X1 U554 ( .A(n1068), .ZN(n712) );
  INV_X1 U555 ( .A(n712), .ZN(n713) );
  INV_X1 U556 ( .A(n712), .ZN(n714) );
  INV_X1 U557 ( .A(n712), .ZN(n715) );
  INV_X1 U558 ( .A(n712), .ZN(n716) );
  INV_X1 U559 ( .A(n712), .ZN(n717) );
  INV_X1 U560 ( .A(n202), .ZN(n718) );
  INV_X1 U561 ( .A(n202), .ZN(n719) );
  INV_X1 U562 ( .A(n202), .ZN(n720) );
  INV_X1 U563 ( .A(n222), .ZN(n721) );
  INV_X1 U564 ( .A(n222), .ZN(n722) );
  INV_X1 U565 ( .A(n222), .ZN(n723) );
  INV_X1 U566 ( .A(n202), .ZN(n724) );
  INV_X1 U567 ( .A(n222), .ZN(n725) );
  INV_X1 U568 ( .A(n781), .ZN(n730) );
  BUF_X1 U569 ( .A(DATAIN[8]), .Z(n781) );
  INV_X1 U570 ( .A(n867), .ZN(n734) );
  INV_X1 U571 ( .A(n869), .ZN(n735) );
  INV_X1 U572 ( .A(n13), .ZN(n736) );
  INV_X1 U573 ( .A(n597), .ZN(n737) );
  CLKBUF_X3 U574 ( .A(DATAIN[13]), .Z(n896) );
  CLKBUF_X3 U575 ( .A(DATAIN[9]), .Z(n780) );
  INV_X1 U576 ( .A(n873), .ZN(n744) );
  BUF_X1 U577 ( .A(DATAIN[19]), .Z(n883) );
  CLKBUF_X3 U578 ( .A(DATAIN[1]), .Z(n902) );
  INV_X1 U579 ( .A(n747), .ZN(n746) );
  INV_X1 U580 ( .A(n3504), .ZN(n747) );
  INV_X1 U581 ( .A(n747), .ZN(n748) );
  INV_X1 U582 ( .A(n176), .ZN(n749) );
  INV_X1 U583 ( .A(n176), .ZN(n750) );
  INV_X1 U584 ( .A(n176), .ZN(n751) );
  INV_X1 U585 ( .A(n3579), .ZN(n752) );
  INV_X1 U586 ( .A(n752), .ZN(n753) );
  INV_X1 U587 ( .A(n754), .ZN(n755) );
  INV_X1 U588 ( .A(n754), .ZN(n756) );
  INV_X1 U589 ( .A(n754), .ZN(n757) );
  CLKBUF_X1 U590 ( .A(n3579), .Z(n3578) );
  INV_X1 U591 ( .A(n3567), .ZN(n758) );
  INV_X1 U592 ( .A(n3567), .ZN(n759) );
  INV_X1 U593 ( .A(n3575), .ZN(n760) );
  INV_X1 U594 ( .A(n3575), .ZN(n761) );
  INV_X1 U595 ( .A(n3639), .ZN(n762) );
  INV_X1 U596 ( .A(n3639), .ZN(n763) );
  INV_X1 U597 ( .A(n3511), .ZN(n764) );
  BUF_X2 U598 ( .A(n1489), .Z(n3511) );
  INV_X1 U599 ( .A(n3587), .ZN(n765) );
  INV_X1 U600 ( .A(n3587), .ZN(n766) );
  BUF_X2 U601 ( .A(n1215), .Z(n3587) );
  INV_X1 U602 ( .A(n3631), .ZN(n767) );
  INV_X1 U603 ( .A(n3631), .ZN(n768) );
  BUF_X2 U604 ( .A(n1108), .Z(n3631) );
  INV_X1 U605 ( .A(n3543), .ZN(n769) );
  INV_X1 U606 ( .A(n3543), .ZN(n770) );
  BUF_X2 U607 ( .A(n1388), .Z(n3543) );
  INV_X1 U608 ( .A(n3501), .ZN(n771) );
  INV_X1 U609 ( .A(n3501), .ZN(n772) );
  BUF_X2 U610 ( .A(n1560), .Z(n3501) );
  INV_X1 U611 ( .A(n3527), .ZN(n773) );
  INV_X1 U612 ( .A(n3527), .ZN(n774) );
  INV_X1 U613 ( .A(n3548), .ZN(n775) );
  INV_X1 U614 ( .A(n3548), .ZN(n776) );
  INV_X1 U615 ( .A(n597), .ZN(n777) );
  INV_X1 U616 ( .A(n13), .ZN(n778) );
  AND3_X1 U617 ( .A1(n681), .A2(n551), .A3(n393), .ZN(n1106) );
  BUF_X2 U618 ( .A(DATAIN[8]), .Z(n782) );
  CLKBUF_X1 U619 ( .A(net33812), .Z(net26419) );
  CLKBUF_X1 U620 ( .A(net33812), .Z(net26421) );
  CLKBUF_X1 U621 ( .A(net33812), .Z(net26423) );
  CLKBUF_X1 U622 ( .A(net33812), .Z(net26425) );
  CLKBUF_X1 U623 ( .A(net33812), .Z(net26427) );
  CLKBUF_X1 U624 ( .A(net33812), .Z(net26429) );
  CLKBUF_X1 U625 ( .A(n783), .Z(n3610) );
  CLKBUF_X1 U626 ( .A(n783), .Z(n3611) );
  CLKBUF_X1 U627 ( .A(n783), .Z(n3609) );
  CLKBUF_X1 U628 ( .A(n783), .Z(n3608) );
  CLKBUF_X1 U629 ( .A(n1388), .Z(n3541) );
  CLKBUF_X1 U630 ( .A(n1388), .Z(n3539) );
  CLKBUF_X1 U631 ( .A(n1284), .Z(n3571) );
  CLKBUF_X1 U632 ( .A(n1456), .Z(n3515) );
  NOR3_X2 U633 ( .A1(n726), .A2(n11), .A3(ADD_WR[2]), .ZN(n1178) );
  INV_X1 U634 ( .A(n3567), .ZN(n3563) );
  INV_X1 U635 ( .A(n3575), .ZN(n3569) );
  INV_X1 U636 ( .A(n13), .ZN(n3596) );
  INV_X1 U637 ( .A(n3550), .ZN(n3545) );
  INV_X1 U638 ( .A(n3543), .ZN(n3537) );
  INV_X1 U639 ( .A(n3635), .ZN(n3633) );
  INV_X1 U640 ( .A(n3631), .ZN(n3624) );
  INV_X1 U641 ( .A(n3567), .ZN(n3562) );
  INV_X1 U642 ( .A(n3575), .ZN(n3568) );
  INV_X1 U643 ( .A(n13), .ZN(n3595) );
  INV_X1 U644 ( .A(n3587), .ZN(n3581) );
  INV_X1 U645 ( .A(n3511), .ZN(n3506) );
  INV_X1 U646 ( .A(n3527), .ZN(n3519) );
  INV_X1 U647 ( .A(n3501), .ZN(n3493) );
  INV_X1 U648 ( .A(n3549), .ZN(n3544) );
  INV_X1 U649 ( .A(n3635), .ZN(n3632) );
  INV_X1 U650 ( .A(n3631), .ZN(n3623) );
  INV_X1 U651 ( .A(n3587), .ZN(n3580) );
  INV_X1 U652 ( .A(n3507), .ZN(n3505) );
  INV_X1 U653 ( .A(n3527), .ZN(n3518) );
  INV_X1 U654 ( .A(n3501), .ZN(n3492) );
  INV_X1 U655 ( .A(net26597), .ZN(net26581) );
  INV_X1 U656 ( .A(net26593), .ZN(net26579) );
  INV_X1 U657 ( .A(n3622), .ZN(n3615) );
  INV_X1 U658 ( .A(n3622), .ZN(n3614) );
  INV_X1 U659 ( .A(n783), .ZN(n3606) );
  INV_X1 U660 ( .A(net33812), .ZN(net26415) );
  INV_X1 U661 ( .A(net33812), .ZN(net26413) );
  INV_X1 U662 ( .A(n783), .ZN(n3605) );
  INV_X1 U663 ( .A(n1351), .ZN(n3555) );
  INV_X1 U664 ( .A(n1350), .ZN(n3556) );
  CLKBUF_X1 U665 ( .A(n1317), .Z(n3566) );
  CLKBUF_X1 U666 ( .A(n13), .Z(n3601) );
  CLKBUF_X1 U667 ( .A(n1215), .Z(n3583) );
  BUF_X1 U668 ( .A(n3655), .Z(n3765) );
  BUF_X1 U669 ( .A(n3655), .Z(n3764) );
  BUF_X1 U670 ( .A(n3654), .Z(n3763) );
  BUF_X1 U671 ( .A(n3654), .Z(n3762) );
  BUF_X1 U672 ( .A(n3653), .Z(n3761) );
  BUF_X1 U673 ( .A(n3653), .Z(n3760) );
  BUF_X1 U674 ( .A(n3652), .Z(n3759) );
  BUF_X1 U675 ( .A(n3652), .Z(n3758) );
  BUF_X1 U676 ( .A(n3651), .Z(n3757) );
  BUF_X1 U677 ( .A(n3651), .Z(n3756) );
  BUF_X1 U678 ( .A(n3650), .Z(n3755) );
  BUF_X1 U679 ( .A(n3650), .Z(n3754) );
  BUF_X1 U680 ( .A(n3649), .Z(n3753) );
  BUF_X1 U681 ( .A(n3649), .Z(n3752) );
  BUF_X1 U682 ( .A(n3648), .Z(n3751) );
  BUF_X1 U683 ( .A(n3648), .Z(n3750) );
  BUF_X1 U684 ( .A(n1630), .Z(n3426) );
  BUF_X1 U685 ( .A(n1630), .Z(n3427) );
  BUF_X1 U686 ( .A(n1635), .Z(n3414) );
  BUF_X1 U687 ( .A(n1635), .Z(n3415) );
  BUF_X1 U688 ( .A(n2221), .Z(n3339) );
  BUF_X1 U689 ( .A(n2226), .Z(n3327) );
  BUF_X1 U690 ( .A(n2221), .Z(n3340) );
  BUF_X1 U691 ( .A(n2226), .Z(n3328) );
  BUF_X1 U692 ( .A(n1620), .Z(n3447) );
  BUF_X1 U693 ( .A(n1620), .Z(n3448) );
  BUF_X1 U694 ( .A(n2211), .Z(n3360) );
  BUF_X1 U695 ( .A(n2211), .Z(n3361) );
  BUF_X1 U696 ( .A(n1603), .Z(n3483) );
  BUF_X1 U697 ( .A(n1608), .Z(net26743) );
  BUF_X1 U698 ( .A(n1613), .Z(n3465) );
  BUF_X1 U699 ( .A(n1618), .Z(n3453) );
  BUF_X1 U700 ( .A(n1628), .Z(n3432) );
  BUF_X1 U701 ( .A(n1603), .Z(n3484) );
  BUF_X1 U702 ( .A(n1608), .Z(net26745) );
  BUF_X1 U703 ( .A(n1613), .Z(n3466) );
  BUF_X1 U704 ( .A(n1618), .Z(n3454) );
  BUF_X1 U705 ( .A(n1628), .Z(n3433) );
  BUF_X1 U706 ( .A(n2194), .Z(n3396) );
  BUF_X1 U707 ( .A(n2199), .Z(net26929) );
  BUF_X1 U708 ( .A(n2204), .Z(n3378) );
  BUF_X1 U709 ( .A(n2209), .Z(n3366) );
  BUF_X1 U710 ( .A(n2219), .Z(n3345) );
  BUF_X1 U711 ( .A(n2194), .Z(n3397) );
  BUF_X1 U712 ( .A(n2199), .Z(net26931) );
  BUF_X1 U713 ( .A(n2204), .Z(n3379) );
  BUF_X1 U714 ( .A(n2209), .Z(n3367) );
  BUF_X1 U715 ( .A(n2219), .Z(n3346) );
  BUF_X1 U716 ( .A(n1631), .Z(n3423) );
  BUF_X1 U717 ( .A(n1636), .Z(n3411) );
  BUF_X1 U718 ( .A(n1631), .Z(n3424) );
  BUF_X1 U719 ( .A(n1636), .Z(n3412) );
  BUF_X1 U720 ( .A(n2222), .Z(n3336) );
  BUF_X1 U721 ( .A(n2227), .Z(n3324) );
  BUF_X1 U722 ( .A(n2222), .Z(n3337) );
  BUF_X1 U723 ( .A(n2227), .Z(n3325) );
  BUF_X1 U724 ( .A(n1600), .Z(n3489) );
  BUF_X1 U725 ( .A(n1605), .Z(n3477) );
  BUF_X1 U726 ( .A(n1610), .Z(n3471) );
  BUF_X1 U727 ( .A(n1615), .Z(n3459) );
  BUF_X1 U728 ( .A(n1625), .Z(n3438) );
  BUF_X1 U729 ( .A(n2191), .Z(n3402) );
  BUF_X1 U730 ( .A(n2196), .Z(n3390) );
  BUF_X1 U731 ( .A(n2201), .Z(n3384) );
  BUF_X1 U732 ( .A(n2206), .Z(n3372) );
  BUF_X1 U733 ( .A(n2216), .Z(n3351) );
  BUF_X1 U734 ( .A(n1604), .Z(n3480) );
  BUF_X1 U735 ( .A(n1609), .Z(net26749) );
  BUF_X1 U736 ( .A(n1614), .Z(n3462) );
  BUF_X1 U737 ( .A(n1619), .Z(n3450) );
  BUF_X1 U738 ( .A(n1629), .Z(n3429) );
  BUF_X1 U739 ( .A(n1604), .Z(n3481) );
  BUF_X1 U740 ( .A(n1609), .Z(net26751) );
  BUF_X1 U741 ( .A(n1614), .Z(n3463) );
  BUF_X1 U742 ( .A(n1619), .Z(n3451) );
  BUF_X1 U743 ( .A(n1629), .Z(n3430) );
  BUF_X1 U744 ( .A(n2195), .Z(n3393) );
  BUF_X1 U745 ( .A(n2200), .Z(net26935) );
  BUF_X1 U746 ( .A(n2205), .Z(n3375) );
  BUF_X1 U747 ( .A(n2210), .Z(n3363) );
  BUF_X1 U748 ( .A(n2220), .Z(n3342) );
  BUF_X1 U749 ( .A(n2195), .Z(n3394) );
  BUF_X1 U750 ( .A(n2200), .Z(net26937) );
  BUF_X1 U751 ( .A(n2205), .Z(n3376) );
  BUF_X1 U752 ( .A(n2210), .Z(n3364) );
  BUF_X1 U753 ( .A(n2220), .Z(n3343) );
  BUF_X1 U754 ( .A(n1601), .Z(n3488) );
  BUF_X1 U755 ( .A(n1606), .Z(n3476) );
  BUF_X1 U756 ( .A(n1611), .Z(n3470) );
  BUF_X1 U757 ( .A(n1616), .Z(n3458) );
  BUF_X1 U758 ( .A(n1626), .Z(n3437) );
  BUF_X1 U759 ( .A(n2192), .Z(n3401) );
  BUF_X1 U760 ( .A(n2197), .Z(n3389) );
  BUF_X1 U761 ( .A(n2202), .Z(n3383) );
  BUF_X1 U762 ( .A(n2207), .Z(n3371) );
  BUF_X1 U763 ( .A(n2217), .Z(n3350) );
  BUF_X1 U764 ( .A(n1630), .Z(n3428) );
  BUF_X1 U765 ( .A(n1635), .Z(n3416) );
  BUF_X1 U766 ( .A(n2221), .Z(n3341) );
  BUF_X1 U767 ( .A(n2226), .Z(n3329) );
  BUF_X1 U768 ( .A(n1620), .Z(n3449) );
  BUF_X1 U769 ( .A(n2211), .Z(n3362) );
  BUF_X1 U770 ( .A(n1603), .Z(n3485) );
  BUF_X1 U771 ( .A(n1608), .Z(net26747) );
  BUF_X1 U772 ( .A(n1613), .Z(n3467) );
  BUF_X1 U773 ( .A(n1618), .Z(n3455) );
  BUF_X1 U774 ( .A(n1628), .Z(n3434) );
  BUF_X1 U775 ( .A(n2194), .Z(n3398) );
  BUF_X1 U776 ( .A(n2199), .Z(net26933) );
  BUF_X1 U777 ( .A(n2204), .Z(n3380) );
  BUF_X1 U778 ( .A(n2209), .Z(n3368) );
  BUF_X1 U779 ( .A(n2219), .Z(n3347) );
  BUF_X1 U780 ( .A(n1631), .Z(n3425) );
  BUF_X1 U781 ( .A(n1636), .Z(n3413) );
  BUF_X1 U782 ( .A(n2222), .Z(n3338) );
  BUF_X1 U783 ( .A(n2227), .Z(n3326) );
  BUF_X1 U784 ( .A(n1600), .Z(n3491) );
  BUF_X1 U785 ( .A(n1605), .Z(n3479) );
  BUF_X1 U786 ( .A(n1610), .Z(n3473) );
  BUF_X1 U787 ( .A(n1615), .Z(n3461) );
  BUF_X1 U788 ( .A(n1625), .Z(n3440) );
  BUF_X1 U789 ( .A(n2191), .Z(n3404) );
  BUF_X1 U790 ( .A(n2196), .Z(n3392) );
  BUF_X1 U791 ( .A(n2201), .Z(n3386) );
  BUF_X1 U792 ( .A(n2206), .Z(n3374) );
  BUF_X1 U793 ( .A(n2216), .Z(n3353) );
  BUF_X1 U794 ( .A(n1604), .Z(n3482) );
  BUF_X1 U795 ( .A(n1609), .Z(net26753) );
  BUF_X1 U797 ( .A(n1614), .Z(n3464) );
  BUF_X1 U798 ( .A(n1619), .Z(n3452) );
  BUF_X1 U799 ( .A(n1629), .Z(n3431) );
  BUF_X1 U800 ( .A(n2195), .Z(n3395) );
  BUF_X1 U801 ( .A(n2200), .Z(net26939) );
  BUF_X1 U802 ( .A(n2205), .Z(n3377) );
  BUF_X1 U803 ( .A(n2210), .Z(n3365) );
  BUF_X1 U804 ( .A(n2220), .Z(n3344) );
  BUF_X1 U805 ( .A(n1623), .Z(n3444) );
  BUF_X1 U806 ( .A(n1638), .Z(n3408) );
  BUF_X1 U807 ( .A(n1623), .Z(n3445) );
  BUF_X1 U808 ( .A(n1638), .Z(n3409) );
  BUF_X1 U809 ( .A(n2214), .Z(n3357) );
  BUF_X1 U810 ( .A(n2229), .Z(n3321) );
  BUF_X1 U811 ( .A(n2214), .Z(n3358) );
  BUF_X1 U812 ( .A(n2229), .Z(n3322) );
  BUF_X1 U813 ( .A(n1633), .Z(n3420) );
  BUF_X1 U814 ( .A(n1633), .Z(n3421) );
  BUF_X1 U815 ( .A(n2224), .Z(n3333) );
  BUF_X1 U816 ( .A(n2224), .Z(n3334) );
  BUF_X1 U817 ( .A(n1624), .Z(n3441) );
  BUF_X1 U818 ( .A(n1639), .Z(n3405) );
  BUF_X1 U819 ( .A(n1624), .Z(n3442) );
  BUF_X1 U820 ( .A(n1639), .Z(n3406) );
  BUF_X1 U821 ( .A(n2215), .Z(n3354) );
  BUF_X1 U822 ( .A(n2230), .Z(n3318) );
  BUF_X1 U823 ( .A(n2215), .Z(n3355) );
  BUF_X1 U824 ( .A(n2230), .Z(n3319) );
  BUF_X1 U825 ( .A(n1634), .Z(n3417) );
  BUF_X1 U826 ( .A(n1634), .Z(n3418) );
  BUF_X1 U827 ( .A(n2225), .Z(n3330) );
  BUF_X1 U828 ( .A(n2225), .Z(n3331) );
  BUF_X1 U829 ( .A(n1623), .Z(n3446) );
  BUF_X1 U830 ( .A(n1638), .Z(n3410) );
  BUF_X1 U831 ( .A(n2214), .Z(n3359) );
  BUF_X1 U832 ( .A(n2229), .Z(n3323) );
  BUF_X1 U833 ( .A(n1633), .Z(n3422) );
  BUF_X1 U834 ( .A(n2224), .Z(n3335) );
  BUF_X1 U835 ( .A(n1624), .Z(n3443) );
  BUF_X1 U836 ( .A(n1639), .Z(n3407) );
  BUF_X1 U837 ( .A(n2215), .Z(n3356) );
  BUF_X1 U838 ( .A(n2230), .Z(n3320) );
  BUF_X1 U839 ( .A(n1634), .Z(n3419) );
  BUF_X1 U840 ( .A(n2225), .Z(n3332) );
  BUF_X1 U841 ( .A(n1601), .Z(n3486) );
  BUF_X1 U842 ( .A(n1606), .Z(n3474) );
  BUF_X1 U843 ( .A(n1611), .Z(n3468) );
  BUF_X1 U844 ( .A(n1616), .Z(n3456) );
  BUF_X1 U845 ( .A(n1626), .Z(n3435) );
  BUF_X1 U846 ( .A(n1601), .Z(n3487) );
  BUF_X1 U847 ( .A(n1606), .Z(n3475) );
  BUF_X1 U848 ( .A(n1611), .Z(n3469) );
  BUF_X1 U849 ( .A(n1616), .Z(n3457) );
  BUF_X1 U850 ( .A(n1626), .Z(n3436) );
  BUF_X1 U851 ( .A(n2192), .Z(n3399) );
  BUF_X1 U852 ( .A(n2197), .Z(n3387) );
  BUF_X1 U853 ( .A(n2202), .Z(n3381) );
  BUF_X1 U854 ( .A(n2207), .Z(n3369) );
  BUF_X1 U855 ( .A(n2217), .Z(n3348) );
  BUF_X1 U856 ( .A(n2192), .Z(n3400) );
  BUF_X1 U857 ( .A(n2197), .Z(n3388) );
  BUF_X1 U858 ( .A(n2202), .Z(n3382) );
  BUF_X1 U859 ( .A(n2207), .Z(n3370) );
  BUF_X1 U860 ( .A(n2217), .Z(n3349) );
  BUF_X1 U861 ( .A(n1600), .Z(n3490) );
  BUF_X1 U862 ( .A(n1605), .Z(n3478) );
  BUF_X1 U863 ( .A(n1610), .Z(n3472) );
  BUF_X1 U865 ( .A(n1615), .Z(n3460) );
  BUF_X1 U866 ( .A(n1625), .Z(n3439) );
  BUF_X1 U867 ( .A(n2191), .Z(n3403) );
  BUF_X1 U868 ( .A(n2196), .Z(n3391) );
  BUF_X1 U869 ( .A(n2201), .Z(n3385) );
  BUF_X1 U870 ( .A(n2216), .Z(n3352) );
  BUF_X1 U871 ( .A(n2206), .Z(n3373) );
  NAND2_X1 U872 ( .A1(n1106), .A2(n1070), .ZN(n1074) );
  NAND2_X1 U873 ( .A1(n414), .A2(n1070), .ZN(n1108) );
  NAND2_X1 U874 ( .A1(n711), .A2(n1070), .ZN(n1180) );
  NAND2_X1 U875 ( .A1(n1069), .A2(n1352), .ZN(n1351) );
  NAND2_X1 U876 ( .A1(n1247), .A2(n1142), .ZN(n1284) );
  NAND2_X1 U877 ( .A1(n711), .A2(n1352), .ZN(n1456) );
  NAND2_X1 U878 ( .A1(n1106), .A2(n1352), .ZN(n1355) );
  NAND2_X1 U879 ( .A1(n1352), .A2(n1140), .ZN(n1388) );
  NAND2_X1 U880 ( .A1(n1144), .A2(n1521), .ZN(n1558) );
  NAND2_X1 U881 ( .A1(n711), .A2(n1247), .ZN(n1350) );
  NAND2_X1 U882 ( .A1(n1352), .A2(n1142), .ZN(n1420) );
  NAND2_X1 U883 ( .A1(n1142), .A2(n1521), .ZN(n1557) );
  BUF_X1 U884 ( .A(n3656), .Z(n3655) );
  BUF_X1 U885 ( .A(n3656), .Z(n3654) );
  BUF_X1 U886 ( .A(n3656), .Z(n3653) );
  BUF_X1 U887 ( .A(n3657), .Z(n3652) );
  BUF_X1 U888 ( .A(n3657), .Z(n3651) );
  BUF_X1 U889 ( .A(n3657), .Z(n3650) );
  BUF_X1 U890 ( .A(n3658), .Z(n3649) );
  BUF_X1 U891 ( .A(n3658), .Z(n3648) );
  NOR3_X1 U892 ( .A1(n726), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n1212) );
  NAND2_X1 U893 ( .A1(n2160), .A2(n2168), .ZN(n1611) );
  NAND2_X1 U894 ( .A1(n2751), .A2(n2759), .ZN(n2202) );
  NAND2_X1 U895 ( .A1(n2160), .A2(n2169), .ZN(n1610) );
  NAND2_X1 U896 ( .A1(n2751), .A2(n2760), .ZN(n2201) );
  INV_X1 U897 ( .A(ADD_WR[2]), .ZN(n4234) );
  INV_X1 U898 ( .A(ADD_WR[0]), .ZN(n4236) );
  NAND2_X1 U899 ( .A1(n2174), .A2(n2160), .ZN(n1624) );
  NAND2_X1 U900 ( .A1(n2175), .A2(n2160), .ZN(n1623) );
  NAND2_X1 U901 ( .A1(n2179), .A2(n2160), .ZN(n1639) );
  NAND2_X1 U902 ( .A1(n2180), .A2(n2160), .ZN(n1638) );
  NAND2_X1 U903 ( .A1(n2765), .A2(n2751), .ZN(n2215) );
  NAND2_X1 U904 ( .A1(n2766), .A2(n2751), .ZN(n2214) );
  NAND2_X1 U905 ( .A1(n2770), .A2(n2751), .ZN(n2230) );
  NAND2_X1 U906 ( .A1(n2771), .A2(n2751), .ZN(n2229) );
  AND2_X1 U907 ( .A1(n2171), .A2(n4242), .ZN(n2168) );
  AND2_X1 U908 ( .A1(n2762), .A2(n4239), .ZN(n2759) );
  NAND2_X1 U909 ( .A1(n2159), .A2(n2162), .ZN(n1601) );
  AND2_X1 U910 ( .A1(n2182), .A2(n4242), .ZN(n2180) );
  AND2_X1 U911 ( .A1(n2773), .A2(n4239), .ZN(n2771) );
  AND2_X1 U912 ( .A1(n2166), .A2(n4242), .ZN(n2159) );
  AND2_X1 U913 ( .A1(n2757), .A2(n4239), .ZN(n2750) );
  NAND2_X1 U914 ( .A1(n2750), .A2(n2753), .ZN(n2192) );
  NAND2_X1 U915 ( .A1(n2159), .A2(n2165), .ZN(n1606) );
  NAND2_X1 U916 ( .A1(n2175), .A2(n2165), .ZN(n1626) );
  NAND2_X1 U917 ( .A1(n2750), .A2(n2756), .ZN(n2197) );
  NAND2_X1 U918 ( .A1(n2766), .A2(n2756), .ZN(n2217) );
  NAND2_X1 U919 ( .A1(n2168), .A2(n2164), .ZN(n1616) );
  NAND2_X1 U920 ( .A1(n2180), .A2(n2164), .ZN(n1633) );
  NAND2_X1 U921 ( .A1(n2179), .A2(n2164), .ZN(n1634) );
  NAND2_X1 U922 ( .A1(n2759), .A2(n2755), .ZN(n2207) );
  NAND2_X1 U923 ( .A1(n2771), .A2(n2755), .ZN(n2224) );
  NAND2_X1 U924 ( .A1(n2770), .A2(n2755), .ZN(n2225) );
  NAND2_X1 U925 ( .A1(n2161), .A2(n2162), .ZN(n1600) );
  NAND2_X1 U926 ( .A1(n2752), .A2(n2753), .ZN(n2191) );
  NAND2_X1 U927 ( .A1(n2164), .A2(n2169), .ZN(n1615) );
  NAND2_X1 U928 ( .A1(n2755), .A2(n2760), .ZN(n2206) );
  AND2_X1 U929 ( .A1(n2177), .A2(n4242), .ZN(n2175) );
  AND2_X1 U930 ( .A1(n2768), .A2(n4239), .ZN(n2766) );
  NAND2_X1 U931 ( .A1(n2161), .A2(n2165), .ZN(n1605) );
  NAND2_X1 U932 ( .A1(n2174), .A2(n2165), .ZN(n1625) );
  NAND2_X1 U933 ( .A1(n2752), .A2(n2756), .ZN(n2196) );
  NAND2_X1 U934 ( .A1(n2765), .A2(n2756), .ZN(n2216) );
  AND2_X1 U935 ( .A1(n2159), .A2(n2160), .ZN(n1604) );
  AND2_X1 U936 ( .A1(n2161), .A2(n2160), .ZN(n1603) );
  AND2_X1 U937 ( .A1(n2750), .A2(n2751), .ZN(n2195) );
  AND2_X1 U938 ( .A1(n2752), .A2(n2751), .ZN(n2194) );
  AND2_X1 U939 ( .A1(n2162), .A2(n2168), .ZN(n1614) );
  AND2_X1 U940 ( .A1(n2162), .A2(n2169), .ZN(n1613) );
  AND2_X1 U941 ( .A1(n2753), .A2(n2759), .ZN(n2205) );
  AND2_X1 U942 ( .A1(n2753), .A2(n2760), .ZN(n2204) );
  AND2_X1 U943 ( .A1(n2174), .A2(n2162), .ZN(n1620) );
  AND2_X1 U944 ( .A1(n2179), .A2(n2162), .ZN(n1635) );
  AND2_X1 U945 ( .A1(n2180), .A2(n2162), .ZN(n1636) );
  AND2_X1 U946 ( .A1(n2765), .A2(n2753), .ZN(n2211) );
  AND2_X1 U947 ( .A1(n2770), .A2(n2753), .ZN(n2226) );
  AND2_X1 U948 ( .A1(n2771), .A2(n2753), .ZN(n2227) );
  AND2_X1 U949 ( .A1(n2165), .A2(n2168), .ZN(n1619) );
  AND2_X1 U950 ( .A1(n2165), .A2(n2169), .ZN(n1618) );
  AND2_X1 U951 ( .A1(n2756), .A2(n2759), .ZN(n2210) );
  AND2_X1 U952 ( .A1(n2756), .A2(n2760), .ZN(n2209) );
  AND2_X1 U953 ( .A1(n2179), .A2(n2165), .ZN(n1630) );
  AND2_X1 U954 ( .A1(n2180), .A2(n2165), .ZN(n1631) );
  AND2_X1 U955 ( .A1(n2770), .A2(n2756), .ZN(n2221) );
  AND2_X1 U956 ( .A1(n2771), .A2(n2756), .ZN(n2222) );
  AND2_X1 U957 ( .A1(n2159), .A2(n2164), .ZN(n1609) );
  AND2_X1 U958 ( .A1(n2161), .A2(n2164), .ZN(n1608) );
  AND2_X1 U959 ( .A1(n2175), .A2(n2164), .ZN(n1629) );
  AND2_X1 U960 ( .A1(n2174), .A2(n2164), .ZN(n1628) );
  AND2_X1 U961 ( .A1(n2750), .A2(n2755), .ZN(n2200) );
  AND2_X1 U962 ( .A1(n2752), .A2(n2755), .ZN(n2199) );
  AND2_X1 U963 ( .A1(n2766), .A2(n2755), .ZN(n2220) );
  AND2_X1 U964 ( .A1(n2765), .A2(n2755), .ZN(n2219) );
  INV_X1 U965 ( .A(ADD_WR[4]), .ZN(n3985) );
  INV_X1 U967 ( .A(ADD_WR[3]), .ZN(n4233) );
  BUF_X1 U968 ( .A(RST_AN), .Z(n3656) );
  BUF_X1 U969 ( .A(RST_AN), .Z(n3657) );
  BUF_X1 U970 ( .A(RST_AN), .Z(n3658) );
  NOR2_X1 U971 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n2162) );
  NOR2_X1 U972 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2753) );
  NOR4_X1 U973 ( .A1(n1780), .A2(n1781), .A3(n1782), .A4(n1783), .ZN(n1779) );
  OAI221_X1 U974 ( .B1(n970), .B2(n3461), .C1(n938), .C2(n3458), .A(n1787), 
        .ZN(n1780) );
  OAI221_X1 U975 ( .B1(n842), .B2(n3473), .C1(n810), .C2(n3470), .A(n1786), 
        .ZN(n1781) );
  OAI221_X1 U976 ( .B1(n650), .B2(n3479), .C1(n618), .C2(n3476), .A(n1785), 
        .ZN(n1782) );
  NOR4_X1 U977 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .ZN(n1762) );
  OAI221_X1 U978 ( .B1(n969), .B2(n3461), .C1(n937), .C2(n3458), .A(n1770), 
        .ZN(n1763) );
  OAI221_X1 U979 ( .B1(n841), .B2(n3473), .C1(n809), .C2(n3470), .A(n1769), 
        .ZN(n1764) );
  OAI221_X1 U980 ( .B1(n649), .B2(n3479), .C1(n617), .C2(n3476), .A(n1768), 
        .ZN(n1765) );
  NOR4_X1 U981 ( .A1(n1746), .A2(n1747), .A3(n1748), .A4(n1749), .ZN(n1745) );
  OAI221_X1 U982 ( .B1(n968), .B2(n3461), .C1(n936), .C2(n3458), .A(n1753), 
        .ZN(n1746) );
  OAI221_X1 U983 ( .B1(n840), .B2(n3473), .C1(n808), .C2(n3470), .A(n1752), 
        .ZN(n1747) );
  OAI221_X1 U984 ( .B1(n648), .B2(n3479), .C1(n616), .C2(n3476), .A(n1751), 
        .ZN(n1748) );
  NOR4_X1 U985 ( .A1(n1729), .A2(n1730), .A3(n1731), .A4(n1732), .ZN(n1728) );
  OAI221_X1 U986 ( .B1(n967), .B2(n3461), .C1(n935), .C2(n3458), .A(n1736), 
        .ZN(n1729) );
  OAI221_X1 U987 ( .B1(n839), .B2(n3473), .C1(n807), .C2(n3470), .A(n1735), 
        .ZN(n1730) );
  OAI221_X1 U988 ( .B1(n647), .B2(n3479), .C1(n615), .C2(n3476), .A(n1734), 
        .ZN(n1731) );
  NOR4_X1 U989 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711) );
  OAI221_X1 U990 ( .B1(n966), .B2(n3461), .C1(n934), .C2(n3458), .A(n1719), 
        .ZN(n1712) );
  OAI221_X1 U991 ( .B1(n838), .B2(n3473), .C1(n806), .C2(n3470), .A(n1718), 
        .ZN(n1713) );
  OAI221_X1 U992 ( .B1(n646), .B2(n3479), .C1(n614), .C2(n3476), .A(n1717), 
        .ZN(n1714) );
  NOR4_X1 U993 ( .A1(n1695), .A2(n1696), .A3(n1697), .A4(n1698), .ZN(n1694) );
  OAI221_X1 U994 ( .B1(n965), .B2(n3461), .C1(n933), .C2(n3458), .A(n1702), 
        .ZN(n1695) );
  OAI221_X1 U995 ( .B1(n837), .B2(n3473), .C1(n805), .C2(n3470), .A(n1701), 
        .ZN(n1696) );
  OAI221_X1 U996 ( .B1(n645), .B2(n3479), .C1(n613), .C2(n3476), .A(n1700), 
        .ZN(n1697) );
  NOR4_X1 U997 ( .A1(n1678), .A2(n1679), .A3(n1680), .A4(n1681), .ZN(n1677) );
  OAI221_X1 U998 ( .B1(n964), .B2(n3461), .C1(n932), .C2(n3458), .A(n1685), 
        .ZN(n1678) );
  OAI221_X1 U999 ( .B1(n836), .B2(n3473), .C1(n804), .C2(n3470), .A(n1684), 
        .ZN(n1679) );
  OAI221_X1 U1001 ( .B1(n644), .B2(n3479), .C1(n612), .C2(n3476), .A(n1683), 
        .ZN(n1680) );
  NOR4_X1 U1002 ( .A1(n1661), .A2(n1662), .A3(n1663), .A4(n1664), .ZN(n1660)
         );
  OAI221_X1 U1003 ( .B1(n963), .B2(n3461), .C1(n931), .C2(n3458), .A(n1668), 
        .ZN(n1661) );
  OAI221_X1 U1004 ( .B1(n835), .B2(n3473), .C1(n803), .C2(n3470), .A(n1667), 
        .ZN(n1662) );
  OAI221_X1 U1005 ( .B1(n643), .B2(n3479), .C1(n611), .C2(n3476), .A(n1666), 
        .ZN(n1663) );
  NOR4_X1 U1006 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .ZN(n1643)
         );
  OAI221_X1 U1007 ( .B1(n962), .B2(n3461), .C1(n930), .C2(n3458), .A(n1651), 
        .ZN(n1644) );
  OAI221_X1 U1008 ( .B1(n834), .B2(n3473), .C1(n802), .C2(n3470), .A(n1650), 
        .ZN(n1645) );
  OAI221_X1 U1009 ( .B1(n642), .B2(n3479), .C1(n610), .C2(n3476), .A(n1649), 
        .ZN(n1646) );
  NOR4_X1 U1010 ( .A1(n1596), .A2(n1597), .A3(n1598), .A4(n1599), .ZN(n1595)
         );
  OAI221_X1 U1011 ( .B1(n961), .B2(n3461), .C1(n929), .C2(n3458), .A(n1617), 
        .ZN(n1596) );
  OAI221_X1 U1012 ( .B1(n833), .B2(n3473), .C1(n801), .C2(n3470), .A(n1612), 
        .ZN(n1597) );
  OAI221_X1 U1013 ( .B1(n641), .B2(n3479), .C1(n609), .C2(n3476), .A(n1607), 
        .ZN(n1598) );
  NOR4_X1 U1014 ( .A1(n2371), .A2(n2372), .A3(n2373), .A4(n2374), .ZN(n2370)
         );
  OAI221_X1 U1015 ( .B1(n970), .B2(n3374), .C1(n938), .C2(n3371), .A(n2378), 
        .ZN(n2371) );
  OAI221_X1 U1016 ( .B1(n842), .B2(n3386), .C1(n810), .C2(n3383), .A(n2377), 
        .ZN(n2372) );
  OAI221_X1 U1017 ( .B1(n650), .B2(n3392), .C1(n618), .C2(n3389), .A(n2376), 
        .ZN(n2373) );
  NOR4_X1 U1018 ( .A1(n2354), .A2(n2355), .A3(n2356), .A4(n2357), .ZN(n2353)
         );
  OAI221_X1 U1019 ( .B1(n969), .B2(n3374), .C1(n937), .C2(n3371), .A(n2361), 
        .ZN(n2354) );
  OAI221_X1 U1020 ( .B1(n841), .B2(n3386), .C1(n809), .C2(n3383), .A(n2360), 
        .ZN(n2355) );
  OAI221_X1 U1021 ( .B1(n649), .B2(n3392), .C1(n617), .C2(n3389), .A(n2359), 
        .ZN(n2356) );
  NOR4_X1 U1022 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n2336)
         );
  OAI221_X1 U1023 ( .B1(n968), .B2(n3374), .C1(n936), .C2(n3371), .A(n2344), 
        .ZN(n2337) );
  OAI221_X1 U1024 ( .B1(n840), .B2(n3386), .C1(n808), .C2(n3383), .A(n2343), 
        .ZN(n2338) );
  OAI221_X1 U1025 ( .B1(n648), .B2(n3392), .C1(n616), .C2(n3389), .A(n2342), 
        .ZN(n2339) );
  NOR4_X1 U1026 ( .A1(n2320), .A2(n2321), .A3(n2322), .A4(n2323), .ZN(n2319)
         );
  OAI221_X1 U1027 ( .B1(n967), .B2(n3374), .C1(n935), .C2(n3371), .A(n2327), 
        .ZN(n2320) );
  OAI221_X1 U1028 ( .B1(n839), .B2(n3386), .C1(n807), .C2(n3383), .A(n2326), 
        .ZN(n2321) );
  OAI221_X1 U1029 ( .B1(n647), .B2(n3392), .C1(n615), .C2(n3389), .A(n2325), 
        .ZN(n2322) );
  NOR4_X1 U1030 ( .A1(n2303), .A2(n2304), .A3(n2305), .A4(n2306), .ZN(n2302)
         );
  OAI221_X1 U1031 ( .B1(n966), .B2(n3374), .C1(n934), .C2(n3371), .A(n2310), 
        .ZN(n2303) );
  OAI221_X1 U1032 ( .B1(n838), .B2(n3386), .C1(n806), .C2(n3383), .A(n2309), 
        .ZN(n2304) );
  OAI221_X1 U1033 ( .B1(n646), .B2(n3392), .C1(n614), .C2(n3389), .A(n2308), 
        .ZN(n2305) );
  NOR4_X1 U1034 ( .A1(n2286), .A2(n2287), .A3(n2288), .A4(n2289), .ZN(n2285)
         );
  OAI221_X1 U1035 ( .B1(n965), .B2(n3374), .C1(n933), .C2(n3371), .A(n2293), 
        .ZN(n2286) );
  OAI221_X1 U1038 ( .B1(n837), .B2(n3386), .C1(n805), .C2(n3383), .A(n2292), 
        .ZN(n2287) );
  OAI221_X1 U1039 ( .B1(n645), .B2(n3392), .C1(n613), .C2(n3389), .A(n2291), 
        .ZN(n2288) );
  NOR4_X1 U1040 ( .A1(n2269), .A2(n2270), .A3(n2271), .A4(n2272), .ZN(n2268)
         );
  OAI221_X1 U1041 ( .B1(n964), .B2(n3374), .C1(n932), .C2(n3371), .A(n2276), 
        .ZN(n2269) );
  OAI221_X1 U1042 ( .B1(n836), .B2(n3386), .C1(n804), .C2(n3383), .A(n2275), 
        .ZN(n2270) );
  OAI221_X1 U1043 ( .B1(n644), .B2(n3392), .C1(n612), .C2(n3389), .A(n2274), 
        .ZN(n2271) );
  NOR4_X1 U1044 ( .A1(n2252), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2251)
         );
  OAI221_X1 U1045 ( .B1(n963), .B2(n3374), .C1(n931), .C2(n3371), .A(n2259), 
        .ZN(n2252) );
  OAI221_X1 U1046 ( .B1(n835), .B2(n3386), .C1(n803), .C2(n3383), .A(n2258), 
        .ZN(n2253) );
  OAI221_X1 U1047 ( .B1(n643), .B2(n3392), .C1(n611), .C2(n3389), .A(n2257), 
        .ZN(n2254) );
  NOR4_X1 U1048 ( .A1(n2235), .A2(n2236), .A3(n2237), .A4(n2238), .ZN(n2234)
         );
  OAI221_X1 U1049 ( .B1(n962), .B2(n3374), .C1(n930), .C2(n3371), .A(n2242), 
        .ZN(n2235) );
  OAI221_X1 U1050 ( .B1(n834), .B2(n3386), .C1(n802), .C2(n3383), .A(n2241), 
        .ZN(n2236) );
  OAI221_X1 U1051 ( .B1(n642), .B2(n3392), .C1(n610), .C2(n3389), .A(n2240), 
        .ZN(n2237) );
  NOR4_X1 U1052 ( .A1(n2187), .A2(n2188), .A3(n2189), .A4(n2190), .ZN(n2186)
         );
  OAI221_X1 U1053 ( .B1(n961), .B2(n3374), .C1(n929), .C2(n3371), .A(n2208), 
        .ZN(n2187) );
  OAI221_X1 U1054 ( .B1(n833), .B2(n3386), .C1(n801), .C2(n3383), .A(n2203), 
        .ZN(n2188) );
  OAI221_X1 U1055 ( .B1(n641), .B2(n3392), .C1(n609), .C2(n3389), .A(n2198), 
        .ZN(n2189) );
  NOR4_X1 U1056 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2153)
         );
  OAI221_X1 U1057 ( .B1(n992), .B2(n3459), .C1(n960), .C2(n3456), .A(n2170), 
        .ZN(n2154) );
  OAI221_X1 U1058 ( .B1(n864), .B2(n3471), .C1(n832), .C2(n3468), .A(n2167), 
        .ZN(n2155) );
  OAI221_X1 U1059 ( .B1(n672), .B2(n3477), .C1(n640), .C2(n3474), .A(n2163), 
        .ZN(n2156) );
  NOR4_X1 U1060 ( .A1(n2137), .A2(n2138), .A3(n2139), .A4(n2140), .ZN(n2136)
         );
  OAI221_X1 U1061 ( .B1(n991), .B2(n3459), .C1(n959), .C2(n3456), .A(n2144), 
        .ZN(n2137) );
  OAI221_X1 U1062 ( .B1(n863), .B2(n3471), .C1(n831), .C2(n3468), .A(n2143), 
        .ZN(n2138) );
  OAI221_X1 U1063 ( .B1(n671), .B2(n3477), .C1(n639), .C2(n3474), .A(n2142), 
        .ZN(n2139) );
  NOR4_X1 U1064 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2119)
         );
  OAI221_X1 U1065 ( .B1(n990), .B2(n3459), .C1(n958), .C2(n3456), .A(n2127), 
        .ZN(n2120) );
  OAI221_X1 U1066 ( .B1(n862), .B2(n3471), .C1(n830), .C2(n3468), .A(n2126), 
        .ZN(n2121) );
  OAI221_X1 U1067 ( .B1(n670), .B2(n3477), .C1(n638), .C2(n3474), .A(n2125), 
        .ZN(n2122) );
  NOR4_X1 U1068 ( .A1(n2103), .A2(n2104), .A3(n2105), .A4(n2106), .ZN(n2102)
         );
  OAI221_X1 U1069 ( .B1(n989), .B2(n3459), .C1(n957), .C2(n3456), .A(n2110), 
        .ZN(n2103) );
  OAI221_X1 U1070 ( .B1(n861), .B2(n3471), .C1(n829), .C2(n3468), .A(n2109), 
        .ZN(n2104) );
  OAI221_X1 U1071 ( .B1(n669), .B2(n3477), .C1(n637), .C2(n3474), .A(n2108), 
        .ZN(n2105) );
  NOR4_X1 U1072 ( .A1(n2086), .A2(n2087), .A3(n2088), .A4(n2089), .ZN(n2085)
         );
  OAI221_X1 U1073 ( .B1(n988), .B2(n3459), .C1(n956), .C2(n3456), .A(n2093), 
        .ZN(n2086) );
  OAI221_X1 U1074 ( .B1(n860), .B2(n3471), .C1(n828), .C2(n3468), .A(n2092), 
        .ZN(n2087) );
  OAI221_X1 U1075 ( .B1(n668), .B2(n3477), .C1(n636), .C2(n3474), .A(n2091), 
        .ZN(n2088) );
  NOR4_X1 U1076 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2068)
         );
  OAI221_X1 U1077 ( .B1(n987), .B2(n3459), .C1(n955), .C2(n3456), .A(n2076), 
        .ZN(n2069) );
  OAI221_X1 U1078 ( .B1(n859), .B2(n3471), .C1(n827), .C2(n3468), .A(n2075), 
        .ZN(n2070) );
  OAI221_X1 U1079 ( .B1(n667), .B2(n3477), .C1(n635), .C2(n3474), .A(n2074), 
        .ZN(n2071) );
  NOR4_X1 U1080 ( .A1(n2052), .A2(n2053), .A3(n2054), .A4(n2055), .ZN(n2051)
         );
  OAI221_X1 U1081 ( .B1(n986), .B2(n3459), .C1(n954), .C2(n3456), .A(n2059), 
        .ZN(n2052) );
  OAI221_X1 U1082 ( .B1(n858), .B2(n3471), .C1(n826), .C2(n3468), .A(n2058), 
        .ZN(n2053) );
  OAI221_X1 U1083 ( .B1(n666), .B2(n3477), .C1(n634), .C2(n3474), .A(n2057), 
        .ZN(n2054) );
  NOR4_X1 U1084 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .ZN(n2034)
         );
  OAI221_X1 U1085 ( .B1(n985), .B2(n3459), .C1(n953), .C2(n3456), .A(n2042), 
        .ZN(n2035) );
  OAI221_X1 U1086 ( .B1(n857), .B2(n3471), .C1(n825), .C2(n3468), .A(n2041), 
        .ZN(n2036) );
  OAI221_X1 U1087 ( .B1(n665), .B2(n3477), .C1(n633), .C2(n3474), .A(n2040), 
        .ZN(n2037) );
  NOR4_X1 U1088 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2017)
         );
  OAI221_X1 U1089 ( .B1(n984), .B2(n3459), .C1(n952), .C2(n3456), .A(n2025), 
        .ZN(n2018) );
  OAI221_X1 U1090 ( .B1(n856), .B2(n3471), .C1(n824), .C2(n3468), .A(n2024), 
        .ZN(n2019) );
  OAI221_X1 U1091 ( .B1(n664), .B2(n3477), .C1(n632), .C2(n3474), .A(n2023), 
        .ZN(n2020) );
  NOR4_X1 U1092 ( .A1(n2001), .A2(n2002), .A3(n2003), .A4(n2004), .ZN(n2000)
         );
  OAI221_X1 U1093 ( .B1(n983), .B2(n3459), .C1(n951), .C2(n3456), .A(n2008), 
        .ZN(n2001) );
  OAI221_X1 U1094 ( .B1(n855), .B2(n3471), .C1(n823), .C2(n3468), .A(n2007), 
        .ZN(n2002) );
  OAI221_X1 U1095 ( .B1(n663), .B2(n3477), .C1(n631), .C2(n3474), .A(n2006), 
        .ZN(n2003) );
  NOR4_X1 U1096 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(n1983)
         );
  OAI221_X1 U1097 ( .B1(n982), .B2(n3459), .C1(n950), .C2(n3456), .A(n1991), 
        .ZN(n1984) );
  OAI221_X1 U1098 ( .B1(n854), .B2(n3471), .C1(n822), .C2(n3468), .A(n1990), 
        .ZN(n1985) );
  OAI221_X1 U1099 ( .B1(n662), .B2(n3477), .C1(n630), .C2(n3474), .A(n1989), 
        .ZN(n1986) );
  NOR4_X1 U1100 ( .A1(n1967), .A2(n1968), .A3(n1969), .A4(n1970), .ZN(n1966)
         );
  OAI221_X1 U1101 ( .B1(n981), .B2(n3460), .C1(n949), .C2(n3457), .A(n1974), 
        .ZN(n1967) );
  OAI221_X1 U1102 ( .B1(n853), .B2(n3472), .C1(n821), .C2(n3469), .A(n1973), 
        .ZN(n1968) );
  OAI221_X1 U1103 ( .B1(n661), .B2(n3478), .C1(n629), .C2(n3475), .A(n1972), 
        .ZN(n1969) );
  NOR4_X1 U1104 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1949)
         );
  OAI221_X1 U1105 ( .B1(n980), .B2(n3460), .C1(n948), .C2(n3457), .A(n1957), 
        .ZN(n1950) );
  OAI221_X1 U1106 ( .B1(n852), .B2(n3472), .C1(n820), .C2(n3469), .A(n1956), 
        .ZN(n1951) );
  OAI221_X1 U1107 ( .B1(n660), .B2(n3478), .C1(n628), .C2(n3475), .A(n1955), 
        .ZN(n1952) );
  NOR4_X1 U1108 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(n1932)
         );
  OAI221_X1 U1109 ( .B1(n979), .B2(n3460), .C1(n947), .C2(n3457), .A(n1940), 
        .ZN(n1933) );
  OAI221_X1 U1110 ( .B1(n851), .B2(n3472), .C1(n819), .C2(n3469), .A(n1939), 
        .ZN(n1934) );
  OAI221_X1 U1111 ( .B1(n659), .B2(n3478), .C1(n627), .C2(n3475), .A(n1938), 
        .ZN(n1935) );
  NOR4_X1 U1112 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(n1915)
         );
  OAI221_X1 U1113 ( .B1(n978), .B2(n3460), .C1(n946), .C2(n3457), .A(n1923), 
        .ZN(n1916) );
  OAI221_X1 U1114 ( .B1(n850), .B2(n3472), .C1(n818), .C2(n3469), .A(n1922), 
        .ZN(n1917) );
  OAI221_X1 U1115 ( .B1(n658), .B2(n3478), .C1(n626), .C2(n3475), .A(n1921), 
        .ZN(n1918) );
  NOR4_X1 U1116 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898)
         );
  OAI221_X1 U1117 ( .B1(n977), .B2(n3460), .C1(n945), .C2(n3457), .A(n1906), 
        .ZN(n1899) );
  OAI221_X1 U1118 ( .B1(n849), .B2(n3472), .C1(n817), .C2(n3469), .A(n1905), 
        .ZN(n1900) );
  OAI221_X1 U1119 ( .B1(n657), .B2(n3478), .C1(n625), .C2(n3475), .A(n1904), 
        .ZN(n1901) );
  NOR4_X1 U1120 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .ZN(n1881)
         );
  OAI221_X1 U1121 ( .B1(n976), .B2(n3460), .C1(n944), .C2(n3457), .A(n1889), 
        .ZN(n1882) );
  OAI221_X1 U1122 ( .B1(n848), .B2(n3472), .C1(n816), .C2(n3469), .A(n1888), 
        .ZN(n1883) );
  OAI221_X1 U1123 ( .B1(n656), .B2(n3478), .C1(n624), .C2(n3475), .A(n1887), 
        .ZN(n1884) );
  NOR4_X1 U1124 ( .A1(n1865), .A2(n1866), .A3(n1867), .A4(n1868), .ZN(n1864)
         );
  OAI221_X1 U1125 ( .B1(n975), .B2(n3460), .C1(n943), .C2(n3457), .A(n1872), 
        .ZN(n1865) );
  OAI221_X1 U1126 ( .B1(n847), .B2(n3472), .C1(n815), .C2(n3469), .A(n1871), 
        .ZN(n1866) );
  OAI221_X1 U1127 ( .B1(n655), .B2(n3478), .C1(n623), .C2(n3475), .A(n1870), 
        .ZN(n1867) );
  NOR4_X1 U1128 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1847)
         );
  OAI221_X1 U1129 ( .B1(n974), .B2(n3460), .C1(n942), .C2(n3457), .A(n1855), 
        .ZN(n1848) );
  OAI221_X1 U1130 ( .B1(n846), .B2(n3472), .C1(n814), .C2(n3469), .A(n1854), 
        .ZN(n1849) );
  OAI221_X1 U1131 ( .B1(n654), .B2(n3478), .C1(n622), .C2(n3475), .A(n1853), 
        .ZN(n1850) );
  NOR4_X1 U1132 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(n1830)
         );
  OAI221_X1 U1133 ( .B1(n973), .B2(n3460), .C1(n941), .C2(n3457), .A(n1838), 
        .ZN(n1831) );
  OAI221_X1 U1134 ( .B1(n845), .B2(n3472), .C1(n813), .C2(n3469), .A(n1837), 
        .ZN(n1832) );
  OAI221_X1 U1135 ( .B1(n653), .B2(n3478), .C1(n621), .C2(n3475), .A(n1836), 
        .ZN(n1833) );
  NOR4_X1 U1136 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .ZN(n1813)
         );
  OAI221_X1 U1137 ( .B1(n972), .B2(n3460), .C1(n940), .C2(n3457), .A(n1821), 
        .ZN(n1814) );
  OAI221_X1 U1138 ( .B1(n844), .B2(n3472), .C1(n812), .C2(n3469), .A(n1820), 
        .ZN(n1815) );
  OAI221_X1 U1139 ( .B1(n652), .B2(n3478), .C1(n620), .C2(n3475), .A(n1819), 
        .ZN(n1816) );
  NOR4_X1 U1140 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1796)
         );
  OAI221_X1 U1141 ( .B1(n971), .B2(n3460), .C1(n939), .C2(n3457), .A(n1804), 
        .ZN(n1797) );
  OAI221_X1 U1142 ( .B1(n843), .B2(n3472), .C1(n811), .C2(n3469), .A(n1803), 
        .ZN(n1798) );
  OAI221_X1 U1143 ( .B1(n651), .B2(n3478), .C1(n619), .C2(n3475), .A(n1802), 
        .ZN(n1799) );
  NOR4_X1 U1144 ( .A1(n2745), .A2(n2746), .A3(n2747), .A4(n2748), .ZN(n2744)
         );
  OAI221_X1 U1145 ( .B1(n992), .B2(n3372), .C1(n960), .C2(n3369), .A(n2761), 
        .ZN(n2745) );
  OAI221_X1 U1146 ( .B1(n864), .B2(n3384), .C1(n832), .C2(n3381), .A(n2758), 
        .ZN(n2746) );
  OAI221_X1 U1147 ( .B1(n672), .B2(n3390), .C1(n640), .C2(n3387), .A(n2754), 
        .ZN(n2747) );
  NOR4_X1 U1148 ( .A1(n2728), .A2(n2729), .A3(n2730), .A4(n2731), .ZN(n2727)
         );
  OAI221_X1 U1149 ( .B1(n991), .B2(n3372), .C1(n959), .C2(n3369), .A(n2735), 
        .ZN(n2728) );
  OAI221_X1 U1150 ( .B1(n863), .B2(n3384), .C1(n831), .C2(n3381), .A(n2734), 
        .ZN(n2729) );
  OAI221_X1 U1151 ( .B1(n671), .B2(n3390), .C1(n639), .C2(n3387), .A(n2733), 
        .ZN(n2730) );
  NOR4_X1 U1152 ( .A1(n2711), .A2(n2712), .A3(n2713), .A4(n2714), .ZN(n2710)
         );
  OAI221_X1 U1153 ( .B1(n990), .B2(n3372), .C1(n958), .C2(n3369), .A(n2718), 
        .ZN(n2711) );
  OAI221_X1 U1154 ( .B1(n862), .B2(n3384), .C1(n830), .C2(n3381), .A(n2717), 
        .ZN(n2712) );
  OAI221_X1 U1155 ( .B1(n670), .B2(n3390), .C1(n638), .C2(n3387), .A(n2716), 
        .ZN(n2713) );
  NOR4_X1 U1156 ( .A1(n2694), .A2(n2695), .A3(n2696), .A4(n2697), .ZN(n2693)
         );
  OAI221_X1 U1157 ( .B1(n989), .B2(n3372), .C1(n957), .C2(n3369), .A(n2701), 
        .ZN(n2694) );
  OAI221_X1 U1158 ( .B1(n861), .B2(n3384), .C1(n829), .C2(n3381), .A(n2700), 
        .ZN(n2695) );
  OAI221_X1 U1159 ( .B1(n669), .B2(n3390), .C1(n637), .C2(n3387), .A(n2699), 
        .ZN(n2696) );
  NOR4_X1 U1160 ( .A1(n2677), .A2(n2678), .A3(n2679), .A4(n2680), .ZN(n2676)
         );
  OAI221_X1 U1161 ( .B1(n988), .B2(n3372), .C1(n956), .C2(n3369), .A(n2684), 
        .ZN(n2677) );
  OAI221_X1 U1162 ( .B1(n860), .B2(n3384), .C1(n828), .C2(n3381), .A(n2683), 
        .ZN(n2678) );
  OAI221_X1 U1163 ( .B1(n668), .B2(n3390), .C1(n636), .C2(n3387), .A(n2682), 
        .ZN(n2679) );
  NOR4_X1 U1164 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(n2659)
         );
  OAI221_X1 U1165 ( .B1(n987), .B2(n3372), .C1(n955), .C2(n3369), .A(n2667), 
        .ZN(n2660) );
  OAI221_X1 U1166 ( .B1(n859), .B2(n3384), .C1(n827), .C2(n3381), .A(n2666), 
        .ZN(n2661) );
  OAI221_X1 U1167 ( .B1(n667), .B2(n3390), .C1(n635), .C2(n3387), .A(n2665), 
        .ZN(n2662) );
  NOR4_X1 U1168 ( .A1(n2643), .A2(n2644), .A3(n2645), .A4(n2646), .ZN(n2642)
         );
  OAI221_X1 U1169 ( .B1(n986), .B2(n3372), .C1(n954), .C2(n3369), .A(n2650), 
        .ZN(n2643) );
  OAI221_X1 U1170 ( .B1(n858), .B2(n3384), .C1(n826), .C2(n3381), .A(n2649), 
        .ZN(n2644) );
  OAI221_X1 U1171 ( .B1(n666), .B2(n3390), .C1(n634), .C2(n3387), .A(n2648), 
        .ZN(n2645) );
  NOR4_X1 U1172 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(n2625)
         );
  OAI221_X1 U1173 ( .B1(n985), .B2(n3372), .C1(n953), .C2(n3369), .A(n2633), 
        .ZN(n2626) );
  OAI221_X1 U1174 ( .B1(n857), .B2(n3384), .C1(n825), .C2(n3381), .A(n2632), 
        .ZN(n2627) );
  OAI221_X1 U1175 ( .B1(n665), .B2(n3390), .C1(n633), .C2(n3387), .A(n2631), 
        .ZN(n2628) );
  NOR4_X1 U1176 ( .A1(n2609), .A2(n2610), .A3(n2611), .A4(n2612), .ZN(n2608)
         );
  OAI221_X1 U1177 ( .B1(n984), .B2(n3372), .C1(n952), .C2(n3369), .A(n2616), 
        .ZN(n2609) );
  OAI221_X1 U1178 ( .B1(n856), .B2(n3384), .C1(n824), .C2(n3381), .A(n2615), 
        .ZN(n2610) );
  OAI221_X1 U1179 ( .B1(n664), .B2(n3390), .C1(n632), .C2(n3387), .A(n2614), 
        .ZN(n2611) );
  NOR4_X1 U1180 ( .A1(n2592), .A2(n2593), .A3(n2594), .A4(n2595), .ZN(n2591)
         );
  OAI221_X1 U1181 ( .B1(n983), .B2(n3372), .C1(n951), .C2(n3369), .A(n2599), 
        .ZN(n2592) );
  OAI221_X1 U1182 ( .B1(n855), .B2(n3384), .C1(n823), .C2(n3381), .A(n2598), 
        .ZN(n2593) );
  OAI221_X1 U1183 ( .B1(n663), .B2(n3390), .C1(n631), .C2(n3387), .A(n2597), 
        .ZN(n2594) );
  NOR4_X1 U1184 ( .A1(n2575), .A2(n2576), .A3(n2577), .A4(n2578), .ZN(n2574)
         );
  OAI221_X1 U1185 ( .B1(n982), .B2(n3372), .C1(n950), .C2(n3369), .A(n2582), 
        .ZN(n2575) );
  OAI221_X1 U1186 ( .B1(n854), .B2(n3384), .C1(n822), .C2(n3381), .A(n2581), 
        .ZN(n2576) );
  OAI221_X1 U1187 ( .B1(n662), .B2(n3390), .C1(n630), .C2(n3387), .A(n2580), 
        .ZN(n2577) );
  NOR4_X1 U1188 ( .A1(n2558), .A2(n2559), .A3(n2560), .A4(n2561), .ZN(n2557)
         );
  OAI221_X1 U1189 ( .B1(n981), .B2(n3373), .C1(n949), .C2(n3370), .A(n2565), 
        .ZN(n2558) );
  OAI221_X1 U1190 ( .B1(n853), .B2(n3385), .C1(n821), .C2(n3382), .A(n2564), 
        .ZN(n2559) );
  OAI221_X1 U1191 ( .B1(n661), .B2(n3391), .C1(n629), .C2(n3388), .A(n2563), 
        .ZN(n2560) );
  NOR4_X1 U1192 ( .A1(n2541), .A2(n2542), .A3(n2543), .A4(n2544), .ZN(n2540)
         );
  OAI221_X1 U1193 ( .B1(n980), .B2(n3373), .C1(n948), .C2(n3370), .A(n2548), 
        .ZN(n2541) );
  OAI221_X1 U1194 ( .B1(n852), .B2(n3385), .C1(n820), .C2(n3382), .A(n2547), 
        .ZN(n2542) );
  OAI221_X1 U1195 ( .B1(n660), .B2(n3391), .C1(n628), .C2(n3388), .A(n2546), 
        .ZN(n2543) );
  NOR4_X1 U1196 ( .A1(n2524), .A2(n2525), .A3(n2526), .A4(n2527), .ZN(n2523)
         );
  OAI221_X1 U1197 ( .B1(n979), .B2(n3373), .C1(n947), .C2(n3370), .A(n2531), 
        .ZN(n2524) );
  OAI221_X1 U1198 ( .B1(n851), .B2(n3385), .C1(n819), .C2(n3382), .A(n2530), 
        .ZN(n2525) );
  OAI221_X1 U1199 ( .B1(n659), .B2(n3391), .C1(n627), .C2(n3388), .A(n2529), 
        .ZN(n2526) );
  NOR4_X1 U1200 ( .A1(n2507), .A2(n2508), .A3(n2509), .A4(n2510), .ZN(n2506)
         );
  OAI221_X1 U1201 ( .B1(n978), .B2(n3373), .C1(n946), .C2(n3370), .A(n2514), 
        .ZN(n2507) );
  OAI221_X1 U1202 ( .B1(n850), .B2(n3385), .C1(n818), .C2(n3382), .A(n2513), 
        .ZN(n2508) );
  OAI221_X1 U1203 ( .B1(n658), .B2(n3391), .C1(n626), .C2(n3388), .A(n2512), 
        .ZN(n2509) );
  NOR4_X1 U1204 ( .A1(n2490), .A2(n2491), .A3(n2492), .A4(n2493), .ZN(n2489)
         );
  OAI221_X1 U1205 ( .B1(n977), .B2(n3373), .C1(n945), .C2(n3370), .A(n2497), 
        .ZN(n2490) );
  OAI221_X1 U1206 ( .B1(n849), .B2(n3385), .C1(n817), .C2(n3382), .A(n2496), 
        .ZN(n2491) );
  OAI221_X1 U1207 ( .B1(n657), .B2(n3391), .C1(n625), .C2(n3388), .A(n2495), 
        .ZN(n2492) );
  NOR4_X1 U1208 ( .A1(n2473), .A2(n2474), .A3(n2475), .A4(n2476), .ZN(n2472)
         );
  OAI221_X1 U1209 ( .B1(n976), .B2(n3373), .C1(n944), .C2(n3370), .A(n2480), 
        .ZN(n2473) );
  OAI221_X1 U1210 ( .B1(n848), .B2(n3385), .C1(n816), .C2(n3382), .A(n2479), 
        .ZN(n2474) );
  OAI221_X1 U1211 ( .B1(n656), .B2(n3391), .C1(n624), .C2(n3388), .A(n2478), 
        .ZN(n2475) );
  NOR4_X1 U1212 ( .A1(n2456), .A2(n2457), .A3(n2458), .A4(n2459), .ZN(n2455)
         );
  OAI221_X1 U1213 ( .B1(n975), .B2(n3373), .C1(n943), .C2(n3370), .A(n2463), 
        .ZN(n2456) );
  OAI221_X1 U1214 ( .B1(n847), .B2(n3385), .C1(n815), .C2(n3382), .A(n2462), 
        .ZN(n2457) );
  OAI221_X1 U1215 ( .B1(n655), .B2(n3391), .C1(n623), .C2(n3388), .A(n2461), 
        .ZN(n2458) );
  NOR4_X1 U1216 ( .A1(n2439), .A2(n2440), .A3(n2441), .A4(n2442), .ZN(n2438)
         );
  OAI221_X1 U1217 ( .B1(n974), .B2(n3373), .C1(n942), .C2(n3370), .A(n2446), 
        .ZN(n2439) );
  OAI221_X1 U1218 ( .B1(n846), .B2(n3385), .C1(n814), .C2(n3382), .A(n2445), 
        .ZN(n2440) );
  OAI221_X1 U1219 ( .B1(n654), .B2(n3391), .C1(n622), .C2(n3388), .A(n2444), 
        .ZN(n2441) );
  NOR4_X1 U1220 ( .A1(n2422), .A2(n2423), .A3(n2424), .A4(n2425), .ZN(n2421)
         );
  OAI221_X1 U1221 ( .B1(n973), .B2(n3373), .C1(n941), .C2(n3370), .A(n2429), 
        .ZN(n2422) );
  OAI221_X1 U1222 ( .B1(n845), .B2(n3385), .C1(n813), .C2(n3382), .A(n2428), 
        .ZN(n2423) );
  OAI221_X1 U1223 ( .B1(n653), .B2(n3391), .C1(n621), .C2(n3388), .A(n2427), 
        .ZN(n2424) );
  NOR4_X1 U1224 ( .A1(n2405), .A2(n2406), .A3(n2407), .A4(n2408), .ZN(n2404)
         );
  OAI221_X1 U1225 ( .B1(n972), .B2(n3373), .C1(n940), .C2(n3370), .A(n2412), 
        .ZN(n2405) );
  OAI221_X1 U1226 ( .B1(n844), .B2(n3385), .C1(n812), .C2(n3382), .A(n2411), 
        .ZN(n2406) );
  OAI221_X1 U1227 ( .B1(n652), .B2(n3391), .C1(n620), .C2(n3388), .A(n2410), 
        .ZN(n2407) );
  NOR4_X1 U1228 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2387)
         );
  OAI221_X1 U1229 ( .B1(n971), .B2(n3373), .C1(n939), .C2(n3370), .A(n2395), 
        .ZN(n2388) );
  OAI221_X1 U1230 ( .B1(n843), .B2(n3385), .C1(n811), .C2(n3382), .A(n2394), 
        .ZN(n2389) );
  OAI221_X1 U1231 ( .B1(n651), .B2(n3391), .C1(n619), .C2(n3388), .A(n2393), 
        .ZN(n2390) );
  OAI221_X1 U1232 ( .B1(n544), .B2(n3489), .C1(n512), .C2(n3486), .A(n2158), 
        .ZN(n2157) );
  AOI22_X1 U1233 ( .A1(n3483), .A2(\registers[19][0] ), .B1(n3480), .B2(
        \registers[18][0] ), .ZN(n2158) );
  OAI221_X1 U1234 ( .B1(n543), .B2(n3489), .C1(n511), .C2(n3486), .A(n2141), 
        .ZN(n2140) );
  AOI22_X1 U1235 ( .A1(n3483), .A2(\registers[19][1] ), .B1(n3480), .B2(
        \registers[18][1] ), .ZN(n2141) );
  OAI221_X1 U1236 ( .B1(n542), .B2(n3489), .C1(n510), .C2(n3486), .A(n2124), 
        .ZN(n2123) );
  AOI22_X1 U1237 ( .A1(n3483), .A2(\registers[19][2] ), .B1(n3480), .B2(
        \registers[18][2] ), .ZN(n2124) );
  OAI221_X1 U1238 ( .B1(n541), .B2(n3489), .C1(n509), .C2(n3486), .A(n2107), 
        .ZN(n2106) );
  AOI22_X1 U1239 ( .A1(n3483), .A2(\registers[19][3] ), .B1(n3480), .B2(
        \registers[18][3] ), .ZN(n2107) );
  OAI221_X1 U1240 ( .B1(n540), .B2(n3489), .C1(n508), .C2(n3486), .A(n2090), 
        .ZN(n2089) );
  AOI22_X1 U1241 ( .A1(n3483), .A2(\registers[19][4] ), .B1(n3480), .B2(
        \registers[18][4] ), .ZN(n2090) );
  OAI221_X1 U1242 ( .B1(n539), .B2(n3489), .C1(n507), .C2(n3486), .A(n2073), 
        .ZN(n2072) );
  AOI22_X1 U1243 ( .A1(n3483), .A2(\registers[19][5] ), .B1(n3480), .B2(
        \registers[18][5] ), .ZN(n2073) );
  OAI221_X1 U1244 ( .B1(n538), .B2(n3489), .C1(n506), .C2(n3486), .A(n2056), 
        .ZN(n2055) );
  AOI22_X1 U1245 ( .A1(n3483), .A2(\registers[19][6] ), .B1(n3480), .B2(
        \registers[18][6] ), .ZN(n2056) );
  OAI221_X1 U1246 ( .B1(n537), .B2(n3489), .C1(n505), .C2(n3486), .A(n2039), 
        .ZN(n2038) );
  AOI22_X1 U1247 ( .A1(n3483), .A2(\registers[19][7] ), .B1(n3480), .B2(
        \registers[18][7] ), .ZN(n2039) );
  OAI221_X1 U1248 ( .B1(n536), .B2(n3489), .C1(n504), .C2(n3486), .A(n2022), 
        .ZN(n2021) );
  AOI22_X1 U1249 ( .A1(n3483), .A2(\registers[19][8] ), .B1(n3480), .B2(
        \registers[18][8] ), .ZN(n2022) );
  OAI221_X1 U1250 ( .B1(n535), .B2(n3489), .C1(n503), .C2(n3486), .A(n2005), 
        .ZN(n2004) );
  AOI22_X1 U1251 ( .A1(n3483), .A2(\registers[19][9] ), .B1(n3480), .B2(
        \registers[18][9] ), .ZN(n2005) );
  OAI221_X1 U1252 ( .B1(n534), .B2(n3489), .C1(n502), .C2(n3486), .A(n1988), 
        .ZN(n1987) );
  AOI22_X1 U1253 ( .A1(n3483), .A2(\registers[19][10] ), .B1(n3480), .B2(
        \registers[18][10] ), .ZN(n1988) );
  OAI221_X1 U1254 ( .B1(n544), .B2(n3402), .C1(n512), .C2(n3399), .A(n2749), 
        .ZN(n2748) );
  AOI22_X1 U1255 ( .A1(n3396), .A2(\registers[19][0] ), .B1(n3393), .B2(
        \registers[18][0] ), .ZN(n2749) );
  OAI221_X1 U1256 ( .B1(n543), .B2(n3402), .C1(n511), .C2(n3399), .A(n2732), 
        .ZN(n2731) );
  AOI22_X1 U1257 ( .A1(n3396), .A2(\registers[19][1] ), .B1(n3393), .B2(
        \registers[18][1] ), .ZN(n2732) );
  OAI221_X1 U1258 ( .B1(n542), .B2(n3402), .C1(n510), .C2(n3399), .A(n2715), 
        .ZN(n2714) );
  AOI22_X1 U1259 ( .A1(n3396), .A2(\registers[19][2] ), .B1(n3393), .B2(
        \registers[18][2] ), .ZN(n2715) );
  OAI221_X1 U1260 ( .B1(n541), .B2(n3402), .C1(n509), .C2(n3399), .A(n2698), 
        .ZN(n2697) );
  AOI22_X1 U1261 ( .A1(n3396), .A2(\registers[19][3] ), .B1(n3393), .B2(
        \registers[18][3] ), .ZN(n2698) );
  OAI221_X1 U1262 ( .B1(n540), .B2(n3402), .C1(n508), .C2(n3399), .A(n2681), 
        .ZN(n2680) );
  AOI22_X1 U1263 ( .A1(n3396), .A2(\registers[19][4] ), .B1(n3393), .B2(
        \registers[18][4] ), .ZN(n2681) );
  OAI221_X1 U1264 ( .B1(n539), .B2(n3402), .C1(n507), .C2(n3399), .A(n2664), 
        .ZN(n2663) );
  AOI22_X1 U1265 ( .A1(n3396), .A2(\registers[19][5] ), .B1(n3393), .B2(
        \registers[18][5] ), .ZN(n2664) );
  OAI221_X1 U1266 ( .B1(n538), .B2(n3402), .C1(n506), .C2(n3399), .A(n2647), 
        .ZN(n2646) );
  AOI22_X1 U1267 ( .A1(n3396), .A2(\registers[19][6] ), .B1(n3393), .B2(
        \registers[18][6] ), .ZN(n2647) );
  OAI221_X1 U1268 ( .B1(n537), .B2(n3402), .C1(n505), .C2(n3399), .A(n2630), 
        .ZN(n2629) );
  AOI22_X1 U1269 ( .A1(n3396), .A2(\registers[19][7] ), .B1(n3393), .B2(
        \registers[18][7] ), .ZN(n2630) );
  OAI221_X1 U1270 ( .B1(n536), .B2(n3402), .C1(n504), .C2(n3399), .A(n2613), 
        .ZN(n2612) );
  AOI22_X1 U1271 ( .A1(n3396), .A2(\registers[19][8] ), .B1(n3393), .B2(
        \registers[18][8] ), .ZN(n2613) );
  OAI221_X1 U1272 ( .B1(n535), .B2(n3402), .C1(n503), .C2(n3399), .A(n2596), 
        .ZN(n2595) );
  AOI22_X1 U1273 ( .A1(n3396), .A2(\registers[19][9] ), .B1(n3393), .B2(
        \registers[18][9] ), .ZN(n2596) );
  OAI221_X1 U1274 ( .B1(n534), .B2(n3402), .C1(n502), .C2(n3399), .A(n2579), 
        .ZN(n2578) );
  AOI22_X1 U1275 ( .A1(n3396), .A2(\registers[19][10] ), .B1(n3393), .B2(
        \registers[18][10] ), .ZN(n2579) );
  OAI221_X1 U1276 ( .B1(n522), .B2(n3491), .C1(n490), .C2(n3488), .A(n1784), 
        .ZN(n1783) );
  AOI22_X1 U1277 ( .A1(n3485), .A2(\registers[19][22] ), .B1(n3482), .B2(
        \registers[18][22] ), .ZN(n1784) );
  OAI221_X1 U1278 ( .B1(n521), .B2(n3491), .C1(n489), .C2(n3488), .A(n1767), 
        .ZN(n1766) );
  AOI22_X1 U1279 ( .A1(n3485), .A2(\registers[19][23] ), .B1(n3482), .B2(
        \registers[18][23] ), .ZN(n1767) );
  OAI221_X1 U1280 ( .B1(n520), .B2(n3491), .C1(n488), .C2(n3488), .A(n1750), 
        .ZN(n1749) );
  AOI22_X1 U1281 ( .A1(n3485), .A2(\registers[19][24] ), .B1(n3482), .B2(
        \registers[18][24] ), .ZN(n1750) );
  OAI221_X1 U1282 ( .B1(n519), .B2(n3491), .C1(n487), .C2(n3488), .A(n1733), 
        .ZN(n1732) );
  AOI22_X1 U1283 ( .A1(n3485), .A2(\registers[19][25] ), .B1(n3482), .B2(
        \registers[18][25] ), .ZN(n1733) );
  OAI221_X1 U1284 ( .B1(n518), .B2(n3491), .C1(n486), .C2(n3488), .A(n1716), 
        .ZN(n1715) );
  AOI22_X1 U1285 ( .A1(n3485), .A2(\registers[19][26] ), .B1(n3482), .B2(
        \registers[18][26] ), .ZN(n1716) );
  OAI221_X1 U1286 ( .B1(n517), .B2(n3491), .C1(n485), .C2(n3488), .A(n1699), 
        .ZN(n1698) );
  AOI22_X1 U1287 ( .A1(n3485), .A2(\registers[19][27] ), .B1(n3482), .B2(
        \registers[18][27] ), .ZN(n1699) );
  OAI221_X1 U1288 ( .B1(n516), .B2(n3491), .C1(n484), .C2(n3488), .A(n1682), 
        .ZN(n1681) );
  AOI22_X1 U1289 ( .A1(n3485), .A2(\registers[19][28] ), .B1(n3482), .B2(
        \registers[18][28] ), .ZN(n1682) );
  OAI221_X1 U1290 ( .B1(n515), .B2(n3491), .C1(n483), .C2(n3488), .A(n1665), 
        .ZN(n1664) );
  AOI22_X1 U1291 ( .A1(n3485), .A2(\registers[19][29] ), .B1(n3482), .B2(
        \registers[18][29] ), .ZN(n1665) );
  OAI221_X1 U1292 ( .B1(n514), .B2(n3491), .C1(n482), .C2(n3488), .A(n1648), 
        .ZN(n1647) );
  AOI22_X1 U1293 ( .A1(n3485), .A2(\registers[19][30] ), .B1(n3482), .B2(
        \registers[18][30] ), .ZN(n1648) );
  OAI221_X1 U1294 ( .B1(n513), .B2(n3491), .C1(n481), .C2(n3488), .A(n1602), 
        .ZN(n1599) );
  AOI22_X1 U1295 ( .A1(n3485), .A2(\registers[19][31] ), .B1(n3482), .B2(
        \registers[18][31] ), .ZN(n1602) );
  OAI221_X1 U1296 ( .B1(n522), .B2(n3404), .C1(n490), .C2(n3401), .A(n2375), 
        .ZN(n2374) );
  AOI22_X1 U1297 ( .A1(n3398), .A2(\registers[19][22] ), .B1(n3395), .B2(
        \registers[18][22] ), .ZN(n2375) );
  OAI221_X1 U1298 ( .B1(n521), .B2(n3404), .C1(n489), .C2(n3401), .A(n2358), 
        .ZN(n2357) );
  AOI22_X1 U1299 ( .A1(n3398), .A2(\registers[19][23] ), .B1(n3395), .B2(
        \registers[18][23] ), .ZN(n2358) );
  OAI221_X1 U1300 ( .B1(n520), .B2(n3404), .C1(n488), .C2(n3401), .A(n2341), 
        .ZN(n2340) );
  AOI22_X1 U1301 ( .A1(n3398), .A2(\registers[19][24] ), .B1(n3395), .B2(
        \registers[18][24] ), .ZN(n2341) );
  OAI221_X1 U1302 ( .B1(n519), .B2(n3404), .C1(n487), .C2(n3401), .A(n2324), 
        .ZN(n2323) );
  AOI22_X1 U1303 ( .A1(n3398), .A2(\registers[19][25] ), .B1(n3395), .B2(
        \registers[18][25] ), .ZN(n2324) );
  OAI221_X1 U1304 ( .B1(n518), .B2(n3404), .C1(n486), .C2(n3401), .A(n2307), 
        .ZN(n2306) );
  AOI22_X1 U1305 ( .A1(n3398), .A2(\registers[19][26] ), .B1(n3395), .B2(
        \registers[18][26] ), .ZN(n2307) );
  OAI221_X1 U1306 ( .B1(n517), .B2(n3404), .C1(n485), .C2(n3401), .A(n2290), 
        .ZN(n2289) );
  AOI22_X1 U1307 ( .A1(n3398), .A2(\registers[19][27] ), .B1(n3395), .B2(
        \registers[18][27] ), .ZN(n2290) );
  OAI221_X1 U1308 ( .B1(n516), .B2(n3404), .C1(n484), .C2(n3401), .A(n2273), 
        .ZN(n2272) );
  AOI22_X1 U1309 ( .A1(n3398), .A2(\registers[19][28] ), .B1(n3395), .B2(
        \registers[18][28] ), .ZN(n2273) );
  OAI221_X1 U1310 ( .B1(n515), .B2(n3404), .C1(n483), .C2(n3401), .A(n2256), 
        .ZN(n2255) );
  AOI22_X1 U1311 ( .A1(n3398), .A2(\registers[19][29] ), .B1(n3395), .B2(
        \registers[18][29] ), .ZN(n2256) );
  OAI221_X1 U1312 ( .B1(n514), .B2(n3404), .C1(n482), .C2(n3401), .A(n2239), 
        .ZN(n2238) );
  AOI22_X1 U1313 ( .A1(n3398), .A2(\registers[19][30] ), .B1(n3395), .B2(
        \registers[18][30] ), .ZN(n2239) );
  OAI221_X1 U1314 ( .B1(n513), .B2(n3404), .C1(n481), .C2(n3401), .A(n2193), 
        .ZN(n2190) );
  AOI22_X1 U1315 ( .A1(n3398), .A2(\registers[19][31] ), .B1(n3395), .B2(
        \registers[18][31] ), .ZN(n2193) );
  OAI221_X1 U1316 ( .B1(n524), .B2(n3490), .C1(n492), .C2(n3487), .A(n1818), 
        .ZN(n1817) );
  AOI22_X1 U1317 ( .A1(n3484), .A2(\registers[19][20] ), .B1(n3481), .B2(
        \registers[18][20] ), .ZN(n1818) );
  OAI221_X1 U1318 ( .B1(n523), .B2(n3490), .C1(n491), .C2(n3487), .A(n1801), 
        .ZN(n1800) );
  AOI22_X1 U1319 ( .A1(n3484), .A2(\registers[19][21] ), .B1(n3481), .B2(
        \registers[18][21] ), .ZN(n1801) );
  OAI221_X1 U1320 ( .B1(n524), .B2(n3403), .C1(n492), .C2(n3400), .A(n2409), 
        .ZN(n2408) );
  AOI22_X1 U1321 ( .A1(n3397), .A2(\registers[19][20] ), .B1(n3394), .B2(
        \registers[18][20] ), .ZN(n2409) );
  OAI221_X1 U1322 ( .B1(n523), .B2(n3403), .C1(n491), .C2(n3400), .A(n2392), 
        .ZN(n2391) );
  AOI22_X1 U1323 ( .A1(n3397), .A2(\registers[19][21] ), .B1(n3394), .B2(
        \registers[18][21] ), .ZN(n2392) );
  OAI221_X1 U1324 ( .B1(n533), .B2(n3490), .C1(n501), .C2(n3487), .A(n1971), 
        .ZN(n1970) );
  AOI22_X1 U1325 ( .A1(n3484), .A2(\registers[19][11] ), .B1(n3481), .B2(
        \registers[18][11] ), .ZN(n1971) );
  OAI221_X1 U1326 ( .B1(n532), .B2(n3490), .C1(n500), .C2(n3487), .A(n1954), 
        .ZN(n1953) );
  AOI22_X1 U1327 ( .A1(n3484), .A2(\registers[19][12] ), .B1(n3481), .B2(
        \registers[18][12] ), .ZN(n1954) );
  OAI221_X1 U1328 ( .B1(n531), .B2(n3490), .C1(n499), .C2(n3487), .A(n1937), 
        .ZN(n1936) );
  AOI22_X1 U1329 ( .A1(n3484), .A2(\registers[19][13] ), .B1(n3481), .B2(
        \registers[18][13] ), .ZN(n1937) );
  OAI221_X1 U1330 ( .B1(n530), .B2(n3490), .C1(n498), .C2(n3487), .A(n1920), 
        .ZN(n1919) );
  AOI22_X1 U1331 ( .A1(n3484), .A2(\registers[19][14] ), .B1(n3481), .B2(
        \registers[18][14] ), .ZN(n1920) );
  OAI221_X1 U1332 ( .B1(n529), .B2(n3490), .C1(n497), .C2(n3487), .A(n1903), 
        .ZN(n1902) );
  AOI22_X1 U1333 ( .A1(n3484), .A2(\registers[19][15] ), .B1(n3481), .B2(
        \registers[18][15] ), .ZN(n1903) );
  OAI221_X1 U1334 ( .B1(n528), .B2(n3490), .C1(n496), .C2(n3487), .A(n1886), 
        .ZN(n1885) );
  AOI22_X1 U1335 ( .A1(n3484), .A2(\registers[19][16] ), .B1(n3481), .B2(
        \registers[18][16] ), .ZN(n1886) );
  OAI221_X1 U1336 ( .B1(n527), .B2(n3490), .C1(n495), .C2(n3487), .A(n1869), 
        .ZN(n1868) );
  AOI22_X1 U1337 ( .A1(n3484), .A2(\registers[19][17] ), .B1(n3481), .B2(
        \registers[18][17] ), .ZN(n1869) );
  OAI221_X1 U1338 ( .B1(n526), .B2(n3490), .C1(n494), .C2(n3487), .A(n1852), 
        .ZN(n1851) );
  AOI22_X1 U1339 ( .A1(n3484), .A2(\registers[19][18] ), .B1(n3481), .B2(
        \registers[18][18] ), .ZN(n1852) );
  OAI221_X1 U1340 ( .B1(n525), .B2(n3490), .C1(n493), .C2(n3487), .A(n1835), 
        .ZN(n1834) );
  AOI22_X1 U1341 ( .A1(n3484), .A2(\registers[19][19] ), .B1(n3481), .B2(
        \registers[18][19] ), .ZN(n1835) );
  OAI221_X1 U1342 ( .B1(n533), .B2(n3403), .C1(n501), .C2(n3400), .A(n2562), 
        .ZN(n2561) );
  AOI22_X1 U1343 ( .A1(n3397), .A2(\registers[19][11] ), .B1(n3394), .B2(
        \registers[18][11] ), .ZN(n2562) );
  OAI221_X1 U1344 ( .B1(n532), .B2(n3403), .C1(n500), .C2(n3400), .A(n2545), 
        .ZN(n2544) );
  AOI22_X1 U1345 ( .A1(n3397), .A2(\registers[19][12] ), .B1(n3394), .B2(
        \registers[18][12] ), .ZN(n2545) );
  OAI221_X1 U1346 ( .B1(n531), .B2(n3403), .C1(n499), .C2(n3400), .A(n2528), 
        .ZN(n2527) );
  AOI22_X1 U1347 ( .A1(n3397), .A2(\registers[19][13] ), .B1(n3394), .B2(
        \registers[18][13] ), .ZN(n2528) );
  OAI221_X1 U1348 ( .B1(n530), .B2(n3403), .C1(n498), .C2(n3400), .A(n2511), 
        .ZN(n2510) );
  AOI22_X1 U1349 ( .A1(n3397), .A2(\registers[19][14] ), .B1(n3394), .B2(
        \registers[18][14] ), .ZN(n2511) );
  OAI221_X1 U1350 ( .B1(n529), .B2(n3403), .C1(n497), .C2(n3400), .A(n2494), 
        .ZN(n2493) );
  AOI22_X1 U1351 ( .A1(n3397), .A2(\registers[19][15] ), .B1(n3394), .B2(
        \registers[18][15] ), .ZN(n2494) );
  OAI221_X1 U1352 ( .B1(n528), .B2(n3403), .C1(n496), .C2(n3400), .A(n2477), 
        .ZN(n2476) );
  AOI22_X1 U1353 ( .A1(n3397), .A2(\registers[19][16] ), .B1(n3394), .B2(
        \registers[18][16] ), .ZN(n2477) );
  OAI221_X1 U1354 ( .B1(n527), .B2(n3403), .C1(n495), .C2(n3400), .A(n2460), 
        .ZN(n2459) );
  AOI22_X1 U1355 ( .A1(n3397), .A2(\registers[19][17] ), .B1(n3394), .B2(
        \registers[18][17] ), .ZN(n2460) );
  OAI221_X1 U1356 ( .B1(n526), .B2(n3403), .C1(n494), .C2(n3400), .A(n2443), 
        .ZN(n2442) );
  AOI22_X1 U1357 ( .A1(n3397), .A2(\registers[19][18] ), .B1(n3394), .B2(
        \registers[18][18] ), .ZN(n2443) );
  OAI221_X1 U1358 ( .B1(n525), .B2(n3403), .C1(n493), .C2(n3400), .A(n2426), 
        .ZN(n2425) );
  AOI22_X1 U1359 ( .A1(n3397), .A2(\registers[19][19] ), .B1(n3394), .B2(
        \registers[18][19] ), .ZN(n2426) );
  OAI221_X1 U1360 ( .B1(n160), .B2(n3438), .C1(n128), .C2(n3435), .A(n2176), 
        .ZN(n2172) );
  AOI22_X1 U1361 ( .A1(n3432), .A2(\registers[7][0] ), .B1(n3429), .B2(
        \registers[6][0] ), .ZN(n2176) );
  OAI221_X1 U1362 ( .B1(n159), .B2(n3438), .C1(n127), .C2(n3435), .A(n2147), 
        .ZN(n2145) );
  AOI22_X1 U1363 ( .A1(n3432), .A2(\registers[7][1] ), .B1(n3429), .B2(
        \registers[6][1] ), .ZN(n2147) );
  OAI221_X1 U1364 ( .B1(n158), .B2(n3438), .C1(n126), .C2(n3435), .A(n2130), 
        .ZN(n2128) );
  AOI22_X1 U1365 ( .A1(n3432), .A2(\registers[7][2] ), .B1(n3429), .B2(
        \registers[6][2] ), .ZN(n2130) );
  OAI221_X1 U1366 ( .B1(n157), .B2(n3438), .C1(n125), .C2(n3435), .A(n2113), 
        .ZN(n2111) );
  AOI22_X1 U1367 ( .A1(n3432), .A2(\registers[7][3] ), .B1(n3429), .B2(
        \registers[6][3] ), .ZN(n2113) );
  OAI221_X1 U1368 ( .B1(n156), .B2(n3438), .C1(n124), .C2(n3435), .A(n2096), 
        .ZN(n2094) );
  AOI22_X1 U1369 ( .A1(n3432), .A2(\registers[7][4] ), .B1(n3429), .B2(
        \registers[6][4] ), .ZN(n2096) );
  OAI221_X1 U1370 ( .B1(n155), .B2(n3438), .C1(n123), .C2(n3435), .A(n2079), 
        .ZN(n2077) );
  AOI22_X1 U1371 ( .A1(n3432), .A2(\registers[7][5] ), .B1(n3429), .B2(
        \registers[6][5] ), .ZN(n2079) );
  OAI221_X1 U1372 ( .B1(n154), .B2(n3438), .C1(n122), .C2(n3435), .A(n2062), 
        .ZN(n2060) );
  AOI22_X1 U1373 ( .A1(n3432), .A2(\registers[7][6] ), .B1(n3429), .B2(
        \registers[6][6] ), .ZN(n2062) );
  OAI221_X1 U1374 ( .B1(n153), .B2(n3438), .C1(n121), .C2(n3435), .A(n2045), 
        .ZN(n2043) );
  AOI22_X1 U1375 ( .A1(n3432), .A2(\registers[7][7] ), .B1(n3429), .B2(
        \registers[6][7] ), .ZN(n2045) );
  OAI221_X1 U1376 ( .B1(n152), .B2(n3438), .C1(n120), .C2(n3435), .A(n2028), 
        .ZN(n2026) );
  AOI22_X1 U1377 ( .A1(n3432), .A2(\registers[7][8] ), .B1(n3429), .B2(
        \registers[6][8] ), .ZN(n2028) );
  OAI221_X1 U1378 ( .B1(n151), .B2(n3438), .C1(n119), .C2(n3435), .A(n2011), 
        .ZN(n2009) );
  AOI22_X1 U1379 ( .A1(n3432), .A2(\registers[7][9] ), .B1(n3429), .B2(
        \registers[6][9] ), .ZN(n2011) );
  OAI221_X1 U1380 ( .B1(n150), .B2(n3438), .C1(n118), .C2(n3435), .A(n1994), 
        .ZN(n1992) );
  AOI22_X1 U1381 ( .A1(n3432), .A2(\registers[7][10] ), .B1(n3429), .B2(
        \registers[6][10] ), .ZN(n1994) );
  OAI221_X1 U1382 ( .B1(n160), .B2(n3351), .C1(n128), .C2(n3348), .A(n2767), 
        .ZN(n2763) );
  AOI22_X1 U1383 ( .A1(n3345), .A2(\registers[7][0] ), .B1(n3342), .B2(
        \registers[6][0] ), .ZN(n2767) );
  OAI221_X1 U1384 ( .B1(n159), .B2(n3351), .C1(n127), .C2(n3348), .A(n2738), 
        .ZN(n2736) );
  AOI22_X1 U1385 ( .A1(n3345), .A2(\registers[7][1] ), .B1(n3342), .B2(
        \registers[6][1] ), .ZN(n2738) );
  OAI221_X1 U1386 ( .B1(n158), .B2(n3351), .C1(n126), .C2(n3348), .A(n2721), 
        .ZN(n2719) );
  AOI22_X1 U1387 ( .A1(n3345), .A2(\registers[7][2] ), .B1(n3342), .B2(
        \registers[6][2] ), .ZN(n2721) );
  OAI221_X1 U1388 ( .B1(n157), .B2(n3351), .C1(n125), .C2(n3348), .A(n2704), 
        .ZN(n2702) );
  AOI22_X1 U1389 ( .A1(n3345), .A2(\registers[7][3] ), .B1(n3342), .B2(
        \registers[6][3] ), .ZN(n2704) );
  OAI221_X1 U1390 ( .B1(n156), .B2(n3351), .C1(n124), .C2(n3348), .A(n2687), 
        .ZN(n2685) );
  AOI22_X1 U1391 ( .A1(n3345), .A2(\registers[7][4] ), .B1(n3342), .B2(
        \registers[6][4] ), .ZN(n2687) );
  OAI221_X1 U1392 ( .B1(n155), .B2(n3351), .C1(n123), .C2(n3348), .A(n2670), 
        .ZN(n2668) );
  AOI22_X1 U1393 ( .A1(n3345), .A2(\registers[7][5] ), .B1(n3342), .B2(
        \registers[6][5] ), .ZN(n2670) );
  OAI221_X1 U1394 ( .B1(n154), .B2(n3351), .C1(n122), .C2(n3348), .A(n2653), 
        .ZN(n2651) );
  AOI22_X1 U1395 ( .A1(n3345), .A2(\registers[7][6] ), .B1(n3342), .B2(
        \registers[6][6] ), .ZN(n2653) );
  OAI221_X1 U1396 ( .B1(n153), .B2(n3351), .C1(n121), .C2(n3348), .A(n2636), 
        .ZN(n2634) );
  AOI22_X1 U1397 ( .A1(n3345), .A2(\registers[7][7] ), .B1(n3342), .B2(
        \registers[6][7] ), .ZN(n2636) );
  OAI221_X1 U1398 ( .B1(n152), .B2(n3351), .C1(n120), .C2(n3348), .A(n2619), 
        .ZN(n2617) );
  AOI22_X1 U1399 ( .A1(n3345), .A2(\registers[7][8] ), .B1(n3342), .B2(
        \registers[6][8] ), .ZN(n2619) );
  OAI221_X1 U1400 ( .B1(n151), .B2(n3351), .C1(n119), .C2(n3348), .A(n2602), 
        .ZN(n2600) );
  AOI22_X1 U1401 ( .A1(n3345), .A2(\registers[7][9] ), .B1(n3342), .B2(
        \registers[6][9] ), .ZN(n2602) );
  OAI221_X1 U1402 ( .B1(n150), .B2(n3351), .C1(n118), .C2(n3348), .A(n2585), 
        .ZN(n2583) );
  AOI22_X1 U1403 ( .A1(n3345), .A2(\registers[7][10] ), .B1(n3342), .B2(
        \registers[6][10] ), .ZN(n2585) );
  OAI221_X1 U1404 ( .B1(n138), .B2(n3440), .C1(n106), .C2(n3437), .A(n1790), 
        .ZN(n1788) );
  AOI22_X1 U1405 ( .A1(n3434), .A2(\registers[7][22] ), .B1(n3431), .B2(
        \registers[6][22] ), .ZN(n1790) );
  OAI221_X1 U1406 ( .B1(n137), .B2(n3440), .C1(n105), .C2(n3437), .A(n1773), 
        .ZN(n1771) );
  AOI22_X1 U1407 ( .A1(n3434), .A2(\registers[7][23] ), .B1(n3431), .B2(
        \registers[6][23] ), .ZN(n1773) );
  OAI221_X1 U1408 ( .B1(n136), .B2(n3440), .C1(n104), .C2(n3437), .A(n1756), 
        .ZN(n1754) );
  AOI22_X1 U1409 ( .A1(n3434), .A2(\registers[7][24] ), .B1(n3431), .B2(
        \registers[6][24] ), .ZN(n1756) );
  OAI221_X1 U1410 ( .B1(n135), .B2(n3440), .C1(n103), .C2(n3437), .A(n1739), 
        .ZN(n1737) );
  AOI22_X1 U1411 ( .A1(n3434), .A2(\registers[7][25] ), .B1(n3431), .B2(
        \registers[6][25] ), .ZN(n1739) );
  OAI221_X1 U1412 ( .B1(n134), .B2(n3440), .C1(n102), .C2(n3437), .A(n1722), 
        .ZN(n1720) );
  AOI22_X1 U1413 ( .A1(n3434), .A2(\registers[7][26] ), .B1(n3431), .B2(
        \registers[6][26] ), .ZN(n1722) );
  OAI221_X1 U1414 ( .B1(n133), .B2(n3440), .C1(n101), .C2(n3437), .A(n1705), 
        .ZN(n1703) );
  AOI22_X1 U1415 ( .A1(n3434), .A2(\registers[7][27] ), .B1(n3431), .B2(
        \registers[6][27] ), .ZN(n1705) );
  OAI221_X1 U1416 ( .B1(n132), .B2(n3440), .C1(n100), .C2(n3437), .A(n1688), 
        .ZN(n1686) );
  AOI22_X1 U1417 ( .A1(n3434), .A2(\registers[7][28] ), .B1(n3431), .B2(
        \registers[6][28] ), .ZN(n1688) );
  OAI221_X1 U1418 ( .B1(n131), .B2(n3440), .C1(n99), .C2(n3437), .A(n1671), 
        .ZN(n1669) );
  AOI22_X1 U1419 ( .A1(n3434), .A2(\registers[7][29] ), .B1(n3431), .B2(
        \registers[6][29] ), .ZN(n1671) );
  OAI221_X1 U1420 ( .B1(n130), .B2(n3440), .C1(n98), .C2(n3437), .A(n1654), 
        .ZN(n1652) );
  AOI22_X1 U1421 ( .A1(n3434), .A2(\registers[7][30] ), .B1(n3431), .B2(
        \registers[6][30] ), .ZN(n1654) );
  OAI221_X1 U1422 ( .B1(n129), .B2(n3440), .C1(n97), .C2(n3437), .A(n1627), 
        .ZN(n1621) );
  AOI22_X1 U1423 ( .A1(n3434), .A2(\registers[7][31] ), .B1(n3431), .B2(
        \registers[6][31] ), .ZN(n1627) );
  OAI221_X1 U1424 ( .B1(n138), .B2(n3353), .C1(n106), .C2(n3350), .A(n2381), 
        .ZN(n2379) );
  AOI22_X1 U1425 ( .A1(n3347), .A2(\registers[7][22] ), .B1(n3344), .B2(
        \registers[6][22] ), .ZN(n2381) );
  OAI221_X1 U1426 ( .B1(n137), .B2(n3353), .C1(n105), .C2(n3350), .A(n2364), 
        .ZN(n2362) );
  AOI22_X1 U1427 ( .A1(n3347), .A2(\registers[7][23] ), .B1(n3344), .B2(
        \registers[6][23] ), .ZN(n2364) );
  OAI221_X1 U1428 ( .B1(n136), .B2(n3353), .C1(n104), .C2(n3350), .A(n2347), 
        .ZN(n2345) );
  AOI22_X1 U1429 ( .A1(n3347), .A2(\registers[7][24] ), .B1(n3344), .B2(
        \registers[6][24] ), .ZN(n2347) );
  OAI221_X1 U1430 ( .B1(n135), .B2(n3353), .C1(n103), .C2(n3350), .A(n2330), 
        .ZN(n2328) );
  AOI22_X1 U1431 ( .A1(n3347), .A2(\registers[7][25] ), .B1(n3344), .B2(
        \registers[6][25] ), .ZN(n2330) );
  OAI221_X1 U1432 ( .B1(n134), .B2(n3353), .C1(n102), .C2(n3350), .A(n2313), 
        .ZN(n2311) );
  AOI22_X1 U1433 ( .A1(n3347), .A2(\registers[7][26] ), .B1(n3344), .B2(
        \registers[6][26] ), .ZN(n2313) );
  OAI221_X1 U1434 ( .B1(n133), .B2(n3353), .C1(n101), .C2(n3350), .A(n2296), 
        .ZN(n2294) );
  AOI22_X1 U1435 ( .A1(n3347), .A2(\registers[7][27] ), .B1(n3344), .B2(
        \registers[6][27] ), .ZN(n2296) );
  OAI221_X1 U1436 ( .B1(n132), .B2(n3353), .C1(n100), .C2(n3350), .A(n2279), 
        .ZN(n2277) );
  AOI22_X1 U1437 ( .A1(n3347), .A2(\registers[7][28] ), .B1(n3344), .B2(
        \registers[6][28] ), .ZN(n2279) );
  OAI221_X1 U1438 ( .B1(n131), .B2(n3353), .C1(n99), .C2(n3350), .A(n2262), 
        .ZN(n2260) );
  AOI22_X1 U1439 ( .A1(n3347), .A2(\registers[7][29] ), .B1(n3344), .B2(
        \registers[6][29] ), .ZN(n2262) );
  OAI221_X1 U1440 ( .B1(n130), .B2(n3353), .C1(n98), .C2(n3350), .A(n2245), 
        .ZN(n2243) );
  AOI22_X1 U1441 ( .A1(n3347), .A2(\registers[7][30] ), .B1(n3344), .B2(
        \registers[6][30] ), .ZN(n2245) );
  OAI221_X1 U1442 ( .B1(n129), .B2(n3353), .C1(n97), .C2(n3350), .A(n2218), 
        .ZN(n2212) );
  AOI22_X1 U1443 ( .A1(n3347), .A2(\registers[7][31] ), .B1(n3344), .B2(
        \registers[6][31] ), .ZN(n2218) );
  OAI221_X1 U1444 ( .B1(n148), .B2(n3439), .C1(n116), .C2(n3436), .A(n1960), 
        .ZN(n1958) );
  AOI22_X1 U1445 ( .A1(n3433), .A2(\registers[7][12] ), .B1(n3430), .B2(
        \registers[6][12] ), .ZN(n1960) );
  OAI221_X1 U1446 ( .B1(n147), .B2(n3439), .C1(n115), .C2(n3436), .A(n1943), 
        .ZN(n1941) );
  AOI22_X1 U1447 ( .A1(n3433), .A2(\registers[7][13] ), .B1(n3430), .B2(
        \registers[6][13] ), .ZN(n1943) );
  OAI221_X1 U1448 ( .B1(n146), .B2(n3439), .C1(n114), .C2(n3436), .A(n1926), 
        .ZN(n1924) );
  AOI22_X1 U1449 ( .A1(n3433), .A2(\registers[7][14] ), .B1(n3430), .B2(
        \registers[6][14] ), .ZN(n1926) );
  OAI221_X1 U1450 ( .B1(n145), .B2(n3439), .C1(n113), .C2(n3436), .A(n1909), 
        .ZN(n1907) );
  AOI22_X1 U1451 ( .A1(n3433), .A2(\registers[7][15] ), .B1(n3430), .B2(
        \registers[6][15] ), .ZN(n1909) );
  OAI221_X1 U1452 ( .B1(n144), .B2(n3439), .C1(n112), .C2(n3436), .A(n1892), 
        .ZN(n1890) );
  AOI22_X1 U1453 ( .A1(n3433), .A2(\registers[7][16] ), .B1(n3430), .B2(
        \registers[6][16] ), .ZN(n1892) );
  OAI221_X1 U1454 ( .B1(n143), .B2(n3439), .C1(n111), .C2(n3436), .A(n1875), 
        .ZN(n1873) );
  AOI22_X1 U1455 ( .A1(n3433), .A2(\registers[7][17] ), .B1(n3430), .B2(
        \registers[6][17] ), .ZN(n1875) );
  OAI221_X1 U1456 ( .B1(n142), .B2(n3439), .C1(n110), .C2(n3436), .A(n1858), 
        .ZN(n1856) );
  AOI22_X1 U1457 ( .A1(n3433), .A2(\registers[7][18] ), .B1(n3430), .B2(
        \registers[6][18] ), .ZN(n1858) );
  OAI221_X1 U1458 ( .B1(n141), .B2(n3439), .C1(n109), .C2(n3436), .A(n1841), 
        .ZN(n1839) );
  AOI22_X1 U1459 ( .A1(n3433), .A2(\registers[7][19] ), .B1(n3430), .B2(
        \registers[6][19] ), .ZN(n1841) );
  OAI221_X1 U1460 ( .B1(n140), .B2(n3439), .C1(n108), .C2(n3436), .A(n1824), 
        .ZN(n1822) );
  AOI22_X1 U1461 ( .A1(n3433), .A2(\registers[7][20] ), .B1(n3430), .B2(
        \registers[6][20] ), .ZN(n1824) );
  OAI221_X1 U1462 ( .B1(n139), .B2(n3439), .C1(n107), .C2(n3436), .A(n1807), 
        .ZN(n1805) );
  AOI22_X1 U1463 ( .A1(n3433), .A2(\registers[7][21] ), .B1(n3430), .B2(
        \registers[6][21] ), .ZN(n1807) );
  OAI221_X1 U1464 ( .B1(n148), .B2(n3352), .C1(n116), .C2(n3349), .A(n2551), 
        .ZN(n2549) );
  AOI22_X1 U1465 ( .A1(n3346), .A2(\registers[7][12] ), .B1(n3343), .B2(
        \registers[6][12] ), .ZN(n2551) );
  OAI221_X1 U1466 ( .B1(n147), .B2(n3352), .C1(n115), .C2(n3349), .A(n2534), 
        .ZN(n2532) );
  AOI22_X1 U1467 ( .A1(n3346), .A2(\registers[7][13] ), .B1(n3343), .B2(
        \registers[6][13] ), .ZN(n2534) );
  OAI221_X1 U1468 ( .B1(n146), .B2(n3352), .C1(n114), .C2(n3349), .A(n2517), 
        .ZN(n2515) );
  AOI22_X1 U1469 ( .A1(n3346), .A2(\registers[7][14] ), .B1(n3343), .B2(
        \registers[6][14] ), .ZN(n2517) );
  OAI221_X1 U1470 ( .B1(n145), .B2(n3352), .C1(n113), .C2(n3349), .A(n2500), 
        .ZN(n2498) );
  AOI22_X1 U1471 ( .A1(n3346), .A2(\registers[7][15] ), .B1(n3343), .B2(
        \registers[6][15] ), .ZN(n2500) );
  OAI221_X1 U1472 ( .B1(n144), .B2(n3352), .C1(n112), .C2(n3349), .A(n2483), 
        .ZN(n2481) );
  AOI22_X1 U1473 ( .A1(n3346), .A2(\registers[7][16] ), .B1(n3343), .B2(
        \registers[6][16] ), .ZN(n2483) );
  OAI221_X1 U1474 ( .B1(n143), .B2(n3352), .C1(n111), .C2(n3349), .A(n2466), 
        .ZN(n2464) );
  AOI22_X1 U1475 ( .A1(n3346), .A2(\registers[7][17] ), .B1(n3343), .B2(
        \registers[6][17] ), .ZN(n2466) );
  OAI221_X1 U1476 ( .B1(n142), .B2(n3352), .C1(n110), .C2(n3349), .A(n2449), 
        .ZN(n2447) );
  AOI22_X1 U1477 ( .A1(n3346), .A2(\registers[7][18] ), .B1(n3343), .B2(
        \registers[6][18] ), .ZN(n2449) );
  OAI221_X1 U1478 ( .B1(n141), .B2(n3352), .C1(n109), .C2(n3349), .A(n2432), 
        .ZN(n2430) );
  AOI22_X1 U1479 ( .A1(n3346), .A2(\registers[7][19] ), .B1(n3343), .B2(
        \registers[6][19] ), .ZN(n2432) );
  OAI221_X1 U1480 ( .B1(n140), .B2(n3352), .C1(n108), .C2(n3349), .A(n2415), 
        .ZN(n2413) );
  AOI22_X1 U1481 ( .A1(n3346), .A2(\registers[7][20] ), .B1(n3343), .B2(
        \registers[6][20] ), .ZN(n2415) );
  OAI221_X1 U1482 ( .B1(n139), .B2(n3352), .C1(n107), .C2(n3349), .A(n2398), 
        .ZN(n2396) );
  AOI22_X1 U1483 ( .A1(n3346), .A2(\registers[7][21] ), .B1(n3343), .B2(
        \registers[6][21] ), .ZN(n2398) );
  OAI221_X1 U1484 ( .B1(n149), .B2(n3439), .C1(n117), .C2(n3436), .A(n1977), 
        .ZN(n1975) );
  AOI22_X1 U1485 ( .A1(n3433), .A2(\registers[7][11] ), .B1(n3430), .B2(
        \registers[6][11] ), .ZN(n1977) );
  OAI221_X1 U1486 ( .B1(n149), .B2(n3352), .C1(n117), .C2(n3349), .A(n2568), 
        .ZN(n2566) );
  AOI22_X1 U1487 ( .A1(n3346), .A2(\registers[7][11] ), .B1(n3343), .B2(
        \registers[6][11] ), .ZN(n2568) );
  OAI22_X1 U1488 ( .A1(n296), .A2(n3410), .B1(n328), .B2(n3407), .ZN(n1758) );
  OAI22_X1 U1489 ( .A1(n295), .A2(n3410), .B1(n327), .B2(n3407), .ZN(n1741) );
  OAI22_X1 U1490 ( .A1(n294), .A2(n3410), .B1(n326), .B2(n3407), .ZN(n1724) );
  OAI22_X1 U1491 ( .A1(n293), .A2(n3410), .B1(n325), .B2(n3407), .ZN(n1707) );
  OAI22_X1 U1492 ( .A1(n292), .A2(n3410), .B1(n324), .B2(n3407), .ZN(n1690) );
  OAI22_X1 U1493 ( .A1(n291), .A2(n3410), .B1(n323), .B2(n3407), .ZN(n1673) );
  OAI22_X1 U1494 ( .A1(n290), .A2(n3410), .B1(n322), .B2(n3407), .ZN(n1656) );
  OAI22_X1 U1495 ( .A1(n289), .A2(n3410), .B1(n321), .B2(n3407), .ZN(n1637) );
  OAI22_X1 U1496 ( .A1(n296), .A2(n3323), .B1(n328), .B2(n3320), .ZN(n2349) );
  OAI22_X1 U1497 ( .A1(n295), .A2(n3323), .B1(n327), .B2(n3320), .ZN(n2332) );
  OAI22_X1 U1498 ( .A1(n294), .A2(n3323), .B1(n326), .B2(n3320), .ZN(n2315) );
  OAI22_X1 U1499 ( .A1(n293), .A2(n3323), .B1(n325), .B2(n3320), .ZN(n2298) );
  OAI22_X1 U1500 ( .A1(n292), .A2(n3323), .B1(n324), .B2(n3320), .ZN(n2281) );
  OAI22_X1 U1501 ( .A1(n291), .A2(n3323), .B1(n323), .B2(n3320), .ZN(n2264) );
  OAI22_X1 U1502 ( .A1(n290), .A2(n3323), .B1(n322), .B2(n3320), .ZN(n2247) );
  OAI22_X1 U1503 ( .A1(n289), .A2(n3323), .B1(n321), .B2(n3320), .ZN(n2228) );
  OAI22_X1 U1504 ( .A1(n424), .A2(n3422), .B1(n456), .B2(n3419), .ZN(n1757) );
  OAI22_X1 U1505 ( .A1(n423), .A2(n3422), .B1(n455), .B2(n3419), .ZN(n1740) );
  OAI22_X1 U1506 ( .A1(n422), .A2(n3422), .B1(n454), .B2(n3419), .ZN(n1723) );
  OAI22_X1 U1507 ( .A1(n421), .A2(n3422), .B1(n453), .B2(n3419), .ZN(n1706) );
  OAI22_X1 U1508 ( .A1(n420), .A2(n3422), .B1(n452), .B2(n3419), .ZN(n1689) );
  OAI22_X1 U1509 ( .A1(n419), .A2(n3422), .B1(n451), .B2(n3419), .ZN(n1672) );
  OAI22_X1 U1510 ( .A1(n418), .A2(n3422), .B1(n450), .B2(n3419), .ZN(n1655) );
  OAI22_X1 U1511 ( .A1(n417), .A2(n3422), .B1(n449), .B2(n3419), .ZN(n1632) );
  OAI22_X1 U1512 ( .A1(n424), .A2(n3335), .B1(n456), .B2(n3332), .ZN(n2348) );
  OAI22_X1 U1513 ( .A1(n423), .A2(n3335), .B1(n455), .B2(n3332), .ZN(n2331) );
  OAI22_X1 U1514 ( .A1(n422), .A2(n3335), .B1(n454), .B2(n3332), .ZN(n2314) );
  OAI22_X1 U1515 ( .A1(n421), .A2(n3335), .B1(n453), .B2(n3332), .ZN(n2297) );
  OAI22_X1 U1516 ( .A1(n420), .A2(n3335), .B1(n452), .B2(n3332), .ZN(n2280) );
  OAI22_X1 U1517 ( .A1(n419), .A2(n3335), .B1(n451), .B2(n3332), .ZN(n2263) );
  OAI22_X1 U1518 ( .A1(n418), .A2(n3335), .B1(n450), .B2(n3332), .ZN(n2246) );
  OAI22_X1 U1519 ( .A1(n417), .A2(n3335), .B1(n449), .B2(n3332), .ZN(n2223) );
  OAI22_X1 U1520 ( .A1(n448), .A2(n3420), .B1(n480), .B2(n3417), .ZN(n2178) );
  OAI22_X1 U1521 ( .A1(n447), .A2(n3420), .B1(n479), .B2(n3417), .ZN(n2148) );
  OAI22_X1 U1522 ( .A1(n446), .A2(n3420), .B1(n478), .B2(n3417), .ZN(n2131) );
  OAI22_X1 U1523 ( .A1(n445), .A2(n3420), .B1(n477), .B2(n3417), .ZN(n2114) );
  OAI22_X1 U1524 ( .A1(n444), .A2(n3420), .B1(n476), .B2(n3417), .ZN(n2097) );
  OAI22_X1 U1525 ( .A1(n443), .A2(n3420), .B1(n475), .B2(n3417), .ZN(n2080) );
  OAI22_X1 U1526 ( .A1(n442), .A2(n3420), .B1(n474), .B2(n3417), .ZN(n2063) );
  OAI22_X1 U1527 ( .A1(n441), .A2(n3420), .B1(n473), .B2(n3417), .ZN(n2046) );
  OAI22_X1 U1528 ( .A1(n440), .A2(n3420), .B1(n472), .B2(n3417), .ZN(n2029) );
  OAI22_X1 U1529 ( .A1(n439), .A2(n3420), .B1(n471), .B2(n3417), .ZN(n2012) );
  OAI22_X1 U1530 ( .A1(n438), .A2(n3420), .B1(n470), .B2(n3417), .ZN(n1995) );
  OAI22_X1 U1531 ( .A1(n437), .A2(n3420), .B1(n469), .B2(n3417), .ZN(n1978) );
  OAI22_X1 U1532 ( .A1(n436), .A2(n3421), .B1(n468), .B2(n3418), .ZN(n1961) );
  OAI22_X1 U1533 ( .A1(n435), .A2(n3421), .B1(n467), .B2(n3418), .ZN(n1944) );
  OAI22_X1 U1534 ( .A1(n434), .A2(n3421), .B1(n466), .B2(n3418), .ZN(n1927) );
  OAI22_X1 U1535 ( .A1(n433), .A2(n3421), .B1(n465), .B2(n3418), .ZN(n1910) );
  OAI22_X1 U1536 ( .A1(n432), .A2(n3421), .B1(n464), .B2(n3418), .ZN(n1893) );
  OAI22_X1 U1537 ( .A1(n431), .A2(n3421), .B1(n463), .B2(n3418), .ZN(n1876) );
  OAI22_X1 U1538 ( .A1(n430), .A2(n3421), .B1(n462), .B2(n3418), .ZN(n1859) );
  OAI22_X1 U1539 ( .A1(n429), .A2(n3421), .B1(n461), .B2(n3418), .ZN(n1842) );
  OAI22_X1 U1540 ( .A1(n448), .A2(n3333), .B1(n480), .B2(n3330), .ZN(n2769) );
  OAI22_X1 U1541 ( .A1(n447), .A2(n3333), .B1(n479), .B2(n3330), .ZN(n2739) );
  OAI22_X1 U1542 ( .A1(n446), .A2(n3333), .B1(n478), .B2(n3330), .ZN(n2722) );
  OAI22_X1 U1543 ( .A1(n445), .A2(n3333), .B1(n477), .B2(n3330), .ZN(n2705) );
  OAI22_X1 U1544 ( .A1(n444), .A2(n3333), .B1(n476), .B2(n3330), .ZN(n2688) );
  OAI22_X1 U1545 ( .A1(n443), .A2(n3333), .B1(n475), .B2(n3330), .ZN(n2671) );
  OAI22_X1 U1546 ( .A1(n442), .A2(n3333), .B1(n474), .B2(n3330), .ZN(n2654) );
  OAI22_X1 U1547 ( .A1(n441), .A2(n3333), .B1(n473), .B2(n3330), .ZN(n2637) );
  OAI22_X1 U1548 ( .A1(n440), .A2(n3333), .B1(n472), .B2(n3330), .ZN(n2620) );
  OAI22_X1 U1549 ( .A1(n439), .A2(n3333), .B1(n471), .B2(n3330), .ZN(n2603) );
  OAI22_X1 U1550 ( .A1(n438), .A2(n3333), .B1(n470), .B2(n3330), .ZN(n2586) );
  OAI22_X1 U1551 ( .A1(n437), .A2(n3333), .B1(n469), .B2(n3330), .ZN(n2569) );
  OAI22_X1 U1552 ( .A1(n436), .A2(n3334), .B1(n468), .B2(n3331), .ZN(n2552) );
  OAI22_X1 U1553 ( .A1(n435), .A2(n3334), .B1(n467), .B2(n3331), .ZN(n2535) );
  OAI22_X1 U1554 ( .A1(n434), .A2(n3334), .B1(n466), .B2(n3331), .ZN(n2518) );
  OAI22_X1 U1555 ( .A1(n433), .A2(n3334), .B1(n465), .B2(n3331), .ZN(n2501) );
  OAI22_X1 U1556 ( .A1(n432), .A2(n3334), .B1(n464), .B2(n3331), .ZN(n2484) );
  OAI22_X1 U1557 ( .A1(n431), .A2(n3334), .B1(n463), .B2(n3331), .ZN(n2467) );
  OAI22_X1 U1558 ( .A1(n430), .A2(n3334), .B1(n462), .B2(n3331), .ZN(n2450) );
  OAI22_X1 U1559 ( .A1(n429), .A2(n3334), .B1(n461), .B2(n3331), .ZN(n2433) );
  OAI22_X1 U1560 ( .A1(n298), .A2(n3409), .B1(n330), .B2(n3406), .ZN(n1792) );
  OAI22_X1 U1561 ( .A1(n297), .A2(n3409), .B1(n329), .B2(n3406), .ZN(n1775) );
  OAI22_X1 U1562 ( .A1(n298), .A2(n3322), .B1(n330), .B2(n3319), .ZN(n2383) );
  OAI22_X1 U1563 ( .A1(n297), .A2(n3322), .B1(n329), .B2(n3319), .ZN(n2366) );
  OAI22_X1 U1564 ( .A1(n320), .A2(n3408), .B1(n352), .B2(n3405), .ZN(n2181) );
  OAI22_X1 U1565 ( .A1(n319), .A2(n3408), .B1(n351), .B2(n3405), .ZN(n2149) );
  OAI22_X1 U1566 ( .A1(n318), .A2(n3408), .B1(n350), .B2(n3405), .ZN(n2132) );
  OAI22_X1 U1567 ( .A1(n317), .A2(n3408), .B1(n349), .B2(n3405), .ZN(n2115) );
  OAI22_X1 U1568 ( .A1(n316), .A2(n3408), .B1(n348), .B2(n3405), .ZN(n2098) );
  OAI22_X1 U1569 ( .A1(n315), .A2(n3408), .B1(n347), .B2(n3405), .ZN(n2081) );
  OAI22_X1 U1570 ( .A1(n314), .A2(n3408), .B1(n346), .B2(n3405), .ZN(n2064) );
  OAI22_X1 U1571 ( .A1(n313), .A2(n3408), .B1(n345), .B2(n3405), .ZN(n2047) );
  OAI22_X1 U1572 ( .A1(n312), .A2(n3408), .B1(n344), .B2(n3405), .ZN(n2030) );
  OAI22_X1 U1573 ( .A1(n311), .A2(n3408), .B1(n343), .B2(n3405), .ZN(n2013) );
  OAI22_X1 U1574 ( .A1(n310), .A2(n3408), .B1(n342), .B2(n3405), .ZN(n1996) );
  OAI22_X1 U1575 ( .A1(n309), .A2(n3408), .B1(n341), .B2(n3405), .ZN(n1979) );
  OAI22_X1 U1576 ( .A1(n308), .A2(n3409), .B1(n340), .B2(n3406), .ZN(n1962) );
  OAI22_X1 U1577 ( .A1(n307), .A2(n3409), .B1(n339), .B2(n3406), .ZN(n1945) );
  OAI22_X1 U1578 ( .A1(n306), .A2(n3409), .B1(n338), .B2(n3406), .ZN(n1928) );
  OAI22_X1 U1579 ( .A1(n305), .A2(n3409), .B1(n337), .B2(n3406), .ZN(n1911) );
  OAI22_X1 U1580 ( .A1(n304), .A2(n3409), .B1(n336), .B2(n3406), .ZN(n1894) );
  OAI22_X1 U1581 ( .A1(n303), .A2(n3409), .B1(n335), .B2(n3406), .ZN(n1877) );
  OAI22_X1 U1582 ( .A1(n302), .A2(n3409), .B1(n334), .B2(n3406), .ZN(n1860) );
  OAI22_X1 U1583 ( .A1(n301), .A2(n3409), .B1(n333), .B2(n3406), .ZN(n1843) );
  OAI22_X1 U1584 ( .A1(n300), .A2(n3409), .B1(n332), .B2(n3406), .ZN(n1826) );
  OAI22_X1 U1585 ( .A1(n299), .A2(n3409), .B1(n331), .B2(n3406), .ZN(n1809) );
  OAI22_X1 U1586 ( .A1(n320), .A2(n3321), .B1(n352), .B2(n3318), .ZN(n2772) );
  OAI22_X1 U1587 ( .A1(n319), .A2(n3321), .B1(n351), .B2(n3318), .ZN(n2740) );
  OAI22_X1 U1588 ( .A1(n318), .A2(n3321), .B1(n350), .B2(n3318), .ZN(n2723) );
  OAI22_X1 U1589 ( .A1(n317), .A2(n3321), .B1(n349), .B2(n3318), .ZN(n2706) );
  OAI22_X1 U1590 ( .A1(n316), .A2(n3321), .B1(n348), .B2(n3318), .ZN(n2689) );
  OAI22_X1 U1591 ( .A1(n315), .A2(n3321), .B1(n347), .B2(n3318), .ZN(n2672) );
  OAI22_X1 U1592 ( .A1(n314), .A2(n3321), .B1(n346), .B2(n3318), .ZN(n2655) );
  OAI22_X1 U1593 ( .A1(n313), .A2(n3321), .B1(n345), .B2(n3318), .ZN(n2638) );
  OAI22_X1 U1594 ( .A1(n312), .A2(n3321), .B1(n344), .B2(n3318), .ZN(n2621) );
  OAI22_X1 U1595 ( .A1(n311), .A2(n3321), .B1(n343), .B2(n3318), .ZN(n2604) );
  OAI22_X1 U1596 ( .A1(n310), .A2(n3321), .B1(n342), .B2(n3318), .ZN(n2587) );
  OAI22_X1 U1597 ( .A1(n309), .A2(n3321), .B1(n341), .B2(n3318), .ZN(n2570) );
  OAI22_X1 U1598 ( .A1(n308), .A2(n3322), .B1(n340), .B2(n3319), .ZN(n2553) );
  OAI22_X1 U1599 ( .A1(n307), .A2(n3322), .B1(n339), .B2(n3319), .ZN(n2536) );
  OAI22_X1 U1600 ( .A1(n306), .A2(n3322), .B1(n338), .B2(n3319), .ZN(n2519) );
  OAI22_X1 U1601 ( .A1(n305), .A2(n3322), .B1(n337), .B2(n3319), .ZN(n2502) );
  OAI22_X1 U1602 ( .A1(n304), .A2(n3322), .B1(n336), .B2(n3319), .ZN(n2485) );
  OAI22_X1 U1603 ( .A1(n303), .A2(n3322), .B1(n335), .B2(n3319), .ZN(n2468) );
  OAI22_X1 U1604 ( .A1(n302), .A2(n3322), .B1(n334), .B2(n3319), .ZN(n2451) );
  OAI22_X1 U1605 ( .A1(n301), .A2(n3322), .B1(n333), .B2(n3319), .ZN(n2434) );
  OAI22_X1 U1606 ( .A1(n300), .A2(n3322), .B1(n332), .B2(n3319), .ZN(n2417) );
  OAI22_X1 U1607 ( .A1(n299), .A2(n3322), .B1(n331), .B2(n3319), .ZN(n2400) );
  OAI22_X1 U1608 ( .A1(n40), .A2(n3446), .B1(n72), .B2(n3443), .ZN(n1755) );
  OAI22_X1 U1609 ( .A1(n39), .A2(n3446), .B1(n71), .B2(n3443), .ZN(n1738) );
  OAI22_X1 U1610 ( .A1(n38), .A2(n3446), .B1(n70), .B2(n3443), .ZN(n1721) );
  OAI22_X1 U1611 ( .A1(n37), .A2(n3446), .B1(n69), .B2(n3443), .ZN(n1704) );
  OAI22_X1 U1612 ( .A1(n36), .A2(n3446), .B1(n68), .B2(n3443), .ZN(n1687) );
  OAI22_X1 U1613 ( .A1(n35), .A2(n3446), .B1(n67), .B2(n3443), .ZN(n1670) );
  OAI22_X1 U1614 ( .A1(n34), .A2(n3446), .B1(n66), .B2(n3443), .ZN(n1653) );
  OAI22_X1 U1615 ( .A1(n33), .A2(n3446), .B1(n65), .B2(n3443), .ZN(n1622) );
  OAI22_X1 U1616 ( .A1(n40), .A2(n3359), .B1(n72), .B2(n3356), .ZN(n2346) );
  OAI22_X1 U1617 ( .A1(n39), .A2(n3359), .B1(n71), .B2(n3356), .ZN(n2329) );
  OAI22_X1 U1618 ( .A1(n38), .A2(n3359), .B1(n70), .B2(n3356), .ZN(n2312) );
  OAI22_X1 U1619 ( .A1(n37), .A2(n3359), .B1(n69), .B2(n3356), .ZN(n2295) );
  OAI22_X1 U1620 ( .A1(n36), .A2(n3359), .B1(n68), .B2(n3356), .ZN(n2278) );
  OAI22_X1 U1621 ( .A1(n35), .A2(n3359), .B1(n67), .B2(n3356), .ZN(n2261) );
  OAI22_X1 U1622 ( .A1(n34), .A2(n3359), .B1(n66), .B2(n3356), .ZN(n2244) );
  OAI22_X1 U1623 ( .A1(n33), .A2(n3359), .B1(n65), .B2(n3356), .ZN(n2213) );
  OAI22_X1 U1624 ( .A1(n426), .A2(n3421), .B1(n458), .B2(n3418), .ZN(n1791) );
  OAI22_X1 U1625 ( .A1(n425), .A2(n3421), .B1(n457), .B2(n3418), .ZN(n1774) );
  OAI22_X1 U1626 ( .A1(n426), .A2(n3334), .B1(n458), .B2(n3331), .ZN(n2382) );
  OAI22_X1 U1627 ( .A1(n425), .A2(n3334), .B1(n457), .B2(n3331), .ZN(n2365) );
  OAI22_X1 U1628 ( .A1(n428), .A2(n3421), .B1(n460), .B2(n3418), .ZN(n1825) );
  OAI22_X1 U1629 ( .A1(n427), .A2(n3421), .B1(n459), .B2(n3418), .ZN(n1808) );
  OAI22_X1 U1630 ( .A1(n428), .A2(n3334), .B1(n460), .B2(n3331), .ZN(n2416) );
  OAI22_X1 U1631 ( .A1(n427), .A2(n3334), .B1(n459), .B2(n3331), .ZN(n2399) );
  OAI22_X1 U1632 ( .A1(n42), .A2(n3445), .B1(n74), .B2(n3442), .ZN(n1789) );
  OAI22_X1 U1633 ( .A1(n41), .A2(n3445), .B1(n73), .B2(n3442), .ZN(n1772) );
  OAI22_X1 U1634 ( .A1(n42), .A2(n3358), .B1(n74), .B2(n3355), .ZN(n2380) );
  OAI22_X1 U1635 ( .A1(n41), .A2(n3358), .B1(n73), .B2(n3355), .ZN(n2363) );
  OAI22_X1 U1636 ( .A1(n64), .A2(n3444), .B1(n96), .B2(n3441), .ZN(n2173) );
  OAI22_X1 U1637 ( .A1(n63), .A2(n3444), .B1(n95), .B2(n3441), .ZN(n2146) );
  OAI22_X1 U1638 ( .A1(n62), .A2(n3444), .B1(n94), .B2(n3441), .ZN(n2129) );
  OAI22_X1 U1639 ( .A1(n61), .A2(n3444), .B1(n93), .B2(n3441), .ZN(n2112) );
  OAI22_X1 U1640 ( .A1(n60), .A2(n3444), .B1(n92), .B2(n3441), .ZN(n2095) );
  OAI22_X1 U1641 ( .A1(n59), .A2(n3444), .B1(n91), .B2(n3441), .ZN(n2078) );
  OAI22_X1 U1642 ( .A1(n58), .A2(n3444), .B1(n90), .B2(n3441), .ZN(n2061) );
  OAI22_X1 U1643 ( .A1(n57), .A2(n3444), .B1(n89), .B2(n3441), .ZN(n2044) );
  OAI22_X1 U1644 ( .A1(n56), .A2(n3444), .B1(n88), .B2(n3441), .ZN(n2027) );
  OAI22_X1 U1645 ( .A1(n55), .A2(n3444), .B1(n87), .B2(n3441), .ZN(n2010) );
  OAI22_X1 U1646 ( .A1(n54), .A2(n3444), .B1(n86), .B2(n3441), .ZN(n1993) );
  OAI22_X1 U1647 ( .A1(n53), .A2(n3444), .B1(n85), .B2(n3441), .ZN(n1976) );
  OAI22_X1 U1648 ( .A1(n52), .A2(n3445), .B1(n84), .B2(n3442), .ZN(n1959) );
  OAI22_X1 U1649 ( .A1(n51), .A2(n3445), .B1(n83), .B2(n3442), .ZN(n1942) );
  OAI22_X1 U1650 ( .A1(n50), .A2(n3445), .B1(n82), .B2(n3442), .ZN(n1925) );
  OAI22_X1 U1651 ( .A1(n49), .A2(n3445), .B1(n81), .B2(n3442), .ZN(n1908) );
  OAI22_X1 U1652 ( .A1(n48), .A2(n3445), .B1(n80), .B2(n3442), .ZN(n1891) );
  OAI22_X1 U1653 ( .A1(n47), .A2(n3445), .B1(n79), .B2(n3442), .ZN(n1874) );
  OAI22_X1 U1654 ( .A1(n46), .A2(n3445), .B1(n78), .B2(n3442), .ZN(n1857) );
  OAI22_X1 U1655 ( .A1(n45), .A2(n3445), .B1(n77), .B2(n3442), .ZN(n1840) );
  OAI22_X1 U1656 ( .A1(n44), .A2(n3445), .B1(n76), .B2(n3442), .ZN(n1823) );
  OAI22_X1 U1657 ( .A1(n43), .A2(n3445), .B1(n75), .B2(n3442), .ZN(n1806) );
  OAI22_X1 U1658 ( .A1(n64), .A2(n3357), .B1(n96), .B2(n3354), .ZN(n2764) );
  OAI22_X1 U1659 ( .A1(n63), .A2(n3357), .B1(n95), .B2(n3354), .ZN(n2737) );
  OAI22_X1 U1660 ( .A1(n62), .A2(n3357), .B1(n94), .B2(n3354), .ZN(n2720) );
  OAI22_X1 U1661 ( .A1(n61), .A2(n3357), .B1(n93), .B2(n3354), .ZN(n2703) );
  OAI22_X1 U1662 ( .A1(n60), .A2(n3357), .B1(n92), .B2(n3354), .ZN(n2686) );
  OAI22_X1 U1663 ( .A1(n59), .A2(n3357), .B1(n91), .B2(n3354), .ZN(n2669) );
  OAI22_X1 U1664 ( .A1(n58), .A2(n3357), .B1(n90), .B2(n3354), .ZN(n2652) );
  OAI22_X1 U1665 ( .A1(n57), .A2(n3357), .B1(n89), .B2(n3354), .ZN(n2635) );
  OAI22_X1 U1666 ( .A1(n56), .A2(n3357), .B1(n88), .B2(n3354), .ZN(n2618) );
  OAI22_X1 U1667 ( .A1(n55), .A2(n3357), .B1(n87), .B2(n3354), .ZN(n2601) );
  OAI22_X1 U1668 ( .A1(n54), .A2(n3357), .B1(n86), .B2(n3354), .ZN(n2584) );
  OAI22_X1 U1669 ( .A1(n53), .A2(n3357), .B1(n85), .B2(n3354), .ZN(n2567) );
  OAI22_X1 U1670 ( .A1(n52), .A2(n3358), .B1(n84), .B2(n3355), .ZN(n2550) );
  OAI22_X1 U1671 ( .A1(n51), .A2(n3358), .B1(n83), .B2(n3355), .ZN(n2533) );
  OAI22_X1 U1672 ( .A1(n50), .A2(n3358), .B1(n82), .B2(n3355), .ZN(n2516) );
  OAI22_X1 U1673 ( .A1(n49), .A2(n3358), .B1(n81), .B2(n3355), .ZN(n2499) );
  OAI22_X1 U1674 ( .A1(n48), .A2(n3358), .B1(n80), .B2(n3355), .ZN(n2482) );
  OAI22_X1 U1675 ( .A1(n47), .A2(n3358), .B1(n79), .B2(n3355), .ZN(n2465) );
  OAI22_X1 U1676 ( .A1(n46), .A2(n3358), .B1(n78), .B2(n3355), .ZN(n2448) );
  OAI22_X1 U1677 ( .A1(n45), .A2(n3358), .B1(n77), .B2(n3355), .ZN(n2431) );
  OAI22_X1 U1678 ( .A1(n44), .A2(n3358), .B1(n76), .B2(n3355), .ZN(n2414) );
  OAI22_X1 U1679 ( .A1(n43), .A2(n3358), .B1(n75), .B2(n3355), .ZN(n2397) );
  OAI22_X1 U1680 ( .A1(n606), .A2(n1031), .B1(n1044), .B2(n480), .ZN(n3030) );
  OAI22_X1 U1681 ( .A1(n673), .A2(n1032), .B1(n1046), .B2(n479), .ZN(n3031) );
  OAI22_X1 U1682 ( .A1(n225), .A2(n1033), .B1(n233), .B2(n478), .ZN(n3032) );
  OAI22_X1 U1683 ( .A1(n4259), .A2(n1038), .B1(n1044), .B2(n468), .ZN(n3042)
         );
  OAI22_X1 U1684 ( .A1(n696), .A2(n1040), .B1(n1046), .B2(n466), .ZN(n3044) );
  OAI22_X1 U1685 ( .A1(n1034), .A2(n552), .B1(n232), .B2(n464), .ZN(n3046) );
  OAI22_X1 U1686 ( .A1(n4254), .A2(n1036), .B1(n233), .B2(n462), .ZN(n3048) );
  OAI22_X1 U1687 ( .A1(n4264), .A2(n1033), .B1(n1045), .B2(n473), .ZN(n3037)
         );
  AOI22_X1 U1688 ( .A1(net26747), .A2(\registers[23][22] ), .B1(net26753), 
        .B2(\registers[22][22] ), .ZN(n1785) );
  AOI22_X1 U1689 ( .A1(net26747), .A2(\registers[23][23] ), .B1(net26753), 
        .B2(\registers[22][23] ), .ZN(n1768) );
  AOI22_X1 U1690 ( .A1(net26747), .A2(\registers[23][24] ), .B1(net26753), 
        .B2(\registers[22][24] ), .ZN(n1751) );
  AOI22_X1 U1691 ( .A1(net26747), .A2(\registers[23][25] ), .B1(net26753), 
        .B2(\registers[22][25] ), .ZN(n1734) );
  AOI22_X1 U1692 ( .A1(net26747), .A2(\registers[23][26] ), .B1(net26753), 
        .B2(\registers[22][26] ), .ZN(n1717) );
  AOI22_X1 U1693 ( .A1(net26747), .A2(\registers[23][27] ), .B1(net26753), 
        .B2(\registers[22][27] ), .ZN(n1700) );
  AOI22_X1 U1694 ( .A1(net26747), .A2(\registers[23][29] ), .B1(net26753), 
        .B2(\registers[22][29] ), .ZN(n1666) );
  AOI22_X1 U1695 ( .A1(net26747), .A2(\registers[23][30] ), .B1(net26753), 
        .B2(\registers[22][30] ), .ZN(n1649) );
  AOI22_X1 U1696 ( .A1(net26747), .A2(\registers[23][31] ), .B1(net26753), 
        .B2(\registers[22][31] ), .ZN(n1607) );
  AOI22_X1 U1697 ( .A1(net26933), .A2(\registers[23][22] ), .B1(net26939), 
        .B2(\registers[22][22] ), .ZN(n2376) );
  AOI22_X1 U1698 ( .A1(net26933), .A2(\registers[23][23] ), .B1(net26939), 
        .B2(\registers[22][23] ), .ZN(n2359) );
  AOI22_X1 U1699 ( .A1(net26933), .A2(\registers[23][24] ), .B1(net26939), 
        .B2(\registers[22][24] ), .ZN(n2342) );
  AOI22_X1 U1700 ( .A1(net26933), .A2(\registers[23][25] ), .B1(net26939), 
        .B2(\registers[22][25] ), .ZN(n2325) );
  AOI22_X1 U1701 ( .A1(net26933), .A2(\registers[23][26] ), .B1(net26939), 
        .B2(\registers[22][26] ), .ZN(n2308) );
  AOI22_X1 U1702 ( .A1(net26933), .A2(\registers[23][27] ), .B1(net26939), 
        .B2(\registers[22][27] ), .ZN(n2291) );
  AOI22_X1 U1703 ( .A1(net26933), .A2(\registers[23][29] ), .B1(net26939), 
        .B2(\registers[22][29] ), .ZN(n2257) );
  AOI22_X1 U1704 ( .A1(net26933), .A2(\registers[23][30] ), .B1(net26939), 
        .B2(\registers[22][30] ), .ZN(n2240) );
  AOI22_X1 U1705 ( .A1(net26933), .A2(\registers[23][31] ), .B1(net26939), 
        .B2(\registers[22][31] ), .ZN(n2198) );
  AOI22_X1 U1706 ( .A1(net26743), .A2(\registers[23][0] ), .B1(net26749), .B2(
        \registers[22][0] ), .ZN(n2163) );
  AOI22_X1 U1707 ( .A1(net26743), .A2(\registers[23][1] ), .B1(net26749), .B2(
        \registers[22][1] ), .ZN(n2142) );
  AOI22_X1 U1708 ( .A1(net26743), .A2(\registers[23][2] ), .B1(net26749), .B2(
        \registers[22][2] ), .ZN(n2125) );
  AOI22_X1 U1709 ( .A1(net26743), .A2(\registers[23][3] ), .B1(net26749), .B2(
        \registers[22][3] ), .ZN(n2108) );
  AOI22_X1 U1710 ( .A1(net26743), .A2(\registers[23][4] ), .B1(net26749), .B2(
        \registers[22][4] ), .ZN(n2091) );
  AOI22_X1 U1711 ( .A1(net26743), .A2(\registers[23][5] ), .B1(net26749), .B2(
        \registers[22][5] ), .ZN(n2074) );
  AOI22_X1 U1712 ( .A1(net26743), .A2(\registers[23][6] ), .B1(net26749), .B2(
        \registers[22][6] ), .ZN(n2057) );
  AOI22_X1 U1713 ( .A1(net26743), .A2(\registers[23][7] ), .B1(net26749), .B2(
        \registers[22][7] ), .ZN(n2040) );
  AOI22_X1 U1714 ( .A1(net26743), .A2(\registers[23][8] ), .B1(net26749), .B2(
        \registers[22][8] ), .ZN(n2023) );
  AOI22_X1 U1715 ( .A1(net26743), .A2(\registers[23][9] ), .B1(net26749), .B2(
        \registers[22][9] ), .ZN(n2006) );
  AOI22_X1 U1716 ( .A1(net26743), .A2(\registers[23][10] ), .B1(net26749), 
        .B2(\registers[22][10] ), .ZN(n1989) );
  AOI22_X1 U1717 ( .A1(net26745), .A2(\registers[23][11] ), .B1(net26751), 
        .B2(\registers[22][11] ), .ZN(n1972) );
  AOI22_X1 U1718 ( .A1(net26745), .A2(\registers[23][12] ), .B1(net26751), 
        .B2(\registers[22][12] ), .ZN(n1955) );
  AOI22_X1 U1719 ( .A1(net26745), .A2(\registers[23][13] ), .B1(net26751), 
        .B2(\registers[22][13] ), .ZN(n1938) );
  AOI22_X1 U1720 ( .A1(net26745), .A2(\registers[23][14] ), .B1(net26751), 
        .B2(\registers[22][14] ), .ZN(n1921) );
  AOI22_X1 U1721 ( .A1(net26745), .A2(\registers[23][15] ), .B1(net26751), 
        .B2(\registers[22][15] ), .ZN(n1904) );
  AOI22_X1 U1722 ( .A1(net26745), .A2(\registers[23][16] ), .B1(net26751), 
        .B2(\registers[22][16] ), .ZN(n1887) );
  AOI22_X1 U1723 ( .A1(net26745), .A2(\registers[23][17] ), .B1(net26751), 
        .B2(\registers[22][17] ), .ZN(n1870) );
  AOI22_X1 U1724 ( .A1(net26745), .A2(\registers[23][18] ), .B1(net26751), 
        .B2(\registers[22][18] ), .ZN(n1853) );
  AOI22_X1 U1725 ( .A1(net26745), .A2(\registers[23][19] ), .B1(net26751), 
        .B2(\registers[22][19] ), .ZN(n1836) );
  AOI22_X1 U1726 ( .A1(net26745), .A2(\registers[23][20] ), .B1(net26751), 
        .B2(\registers[22][20] ), .ZN(n1819) );
  AOI22_X1 U1727 ( .A1(net26745), .A2(\registers[23][21] ), .B1(net26751), 
        .B2(\registers[22][21] ), .ZN(n1802) );
  AOI22_X1 U1728 ( .A1(net26929), .A2(\registers[23][0] ), .B1(net26935), .B2(
        \registers[22][0] ), .ZN(n2754) );
  AOI22_X1 U1729 ( .A1(net26929), .A2(\registers[23][1] ), .B1(net26935), .B2(
        \registers[22][1] ), .ZN(n2733) );
  AOI22_X1 U1730 ( .A1(net26929), .A2(\registers[23][2] ), .B1(net26935), .B2(
        \registers[22][2] ), .ZN(n2716) );
  AOI22_X1 U1731 ( .A1(net26929), .A2(\registers[23][3] ), .B1(net26935), .B2(
        \registers[22][3] ), .ZN(n2699) );
  AOI22_X1 U1732 ( .A1(net26929), .A2(\registers[23][4] ), .B1(net26935), .B2(
        \registers[22][4] ), .ZN(n2682) );
  AOI22_X1 U1733 ( .A1(net26929), .A2(\registers[23][5] ), .B1(net26935), .B2(
        \registers[22][5] ), .ZN(n2665) );
  AOI22_X1 U1734 ( .A1(net26929), .A2(\registers[23][6] ), .B1(net26935), .B2(
        \registers[22][6] ), .ZN(n2648) );
  AOI22_X1 U1735 ( .A1(net26929), .A2(\registers[23][7] ), .B1(net26935), .B2(
        \registers[22][7] ), .ZN(n2631) );
  AOI22_X1 U1736 ( .A1(net26929), .A2(\registers[23][8] ), .B1(net26935), .B2(
        \registers[22][8] ), .ZN(n2614) );
  AOI22_X1 U1737 ( .A1(net26929), .A2(\registers[23][9] ), .B1(net26935), .B2(
        \registers[22][9] ), .ZN(n2597) );
  AOI22_X1 U1738 ( .A1(net26929), .A2(\registers[23][10] ), .B1(net26935), 
        .B2(\registers[22][10] ), .ZN(n2580) );
  AOI22_X1 U1739 ( .A1(net26931), .A2(\registers[23][11] ), .B1(net26937), 
        .B2(\registers[22][11] ), .ZN(n2563) );
  AOI22_X1 U1740 ( .A1(net26931), .A2(\registers[23][12] ), .B1(net26937), 
        .B2(\registers[22][12] ), .ZN(n2546) );
  AOI22_X1 U1741 ( .A1(net26931), .A2(\registers[23][13] ), .B1(net26937), 
        .B2(\registers[22][13] ), .ZN(n2529) );
  AOI22_X1 U1742 ( .A1(net26931), .A2(\registers[23][14] ), .B1(net26937), 
        .B2(\registers[22][14] ), .ZN(n2512) );
  AOI22_X1 U1743 ( .A1(net26931), .A2(\registers[23][15] ), .B1(net26937), 
        .B2(\registers[22][15] ), .ZN(n2495) );
  AOI22_X1 U1744 ( .A1(net26931), .A2(\registers[23][16] ), .B1(net26937), 
        .B2(\registers[22][16] ), .ZN(n2478) );
  AOI22_X1 U1745 ( .A1(net26931), .A2(\registers[23][17] ), .B1(net26937), 
        .B2(\registers[22][17] ), .ZN(n2461) );
  AOI22_X1 U1746 ( .A1(net26931), .A2(\registers[23][18] ), .B1(net26937), 
        .B2(\registers[22][18] ), .ZN(n2444) );
  AOI22_X1 U1747 ( .A1(net26931), .A2(\registers[23][19] ), .B1(net26937), 
        .B2(\registers[22][19] ), .ZN(n2427) );
  AOI22_X1 U1748 ( .A1(net26931), .A2(\registers[23][20] ), .B1(net26937), 
        .B2(\registers[22][20] ), .ZN(n2410) );
  AOI22_X1 U1749 ( .A1(net26931), .A2(\registers[23][21] ), .B1(net26937), 
        .B2(\registers[22][21] ), .ZN(n2393) );
  AOI22_X1 U1750 ( .A1(n3467), .A2(\registers[25][22] ), .B1(n3464), .B2(
        \registers[24][22] ), .ZN(n1786) );
  AOI22_X1 U1751 ( .A1(n3467), .A2(\registers[25][23] ), .B1(n3464), .B2(
        \registers[24][23] ), .ZN(n1769) );
  AOI22_X1 U1752 ( .A1(n3467), .A2(\registers[25][24] ), .B1(n3464), .B2(
        \registers[24][24] ), .ZN(n1752) );
  AOI22_X1 U1753 ( .A1(n3467), .A2(\registers[25][25] ), .B1(n3464), .B2(
        \registers[24][25] ), .ZN(n1735) );
  AOI22_X1 U1754 ( .A1(n3467), .A2(\registers[25][26] ), .B1(n3464), .B2(
        \registers[24][26] ), .ZN(n1718) );
  AOI22_X1 U1755 ( .A1(n3467), .A2(\registers[25][27] ), .B1(n3464), .B2(
        \registers[24][27] ), .ZN(n1701) );
  AOI22_X1 U1756 ( .A1(n3467), .A2(\registers[25][28] ), .B1(n3464), .B2(
        \registers[24][28] ), .ZN(n1684) );
  AOI22_X1 U1757 ( .A1(n3467), .A2(\registers[25][29] ), .B1(n3464), .B2(
        \registers[24][29] ), .ZN(n1667) );
  AOI22_X1 U1758 ( .A1(n3467), .A2(\registers[25][30] ), .B1(n3464), .B2(
        \registers[24][30] ), .ZN(n1650) );
  AOI22_X1 U1759 ( .A1(n3467), .A2(\registers[25][31] ), .B1(n3464), .B2(
        \registers[24][31] ), .ZN(n1612) );
  AOI22_X1 U1760 ( .A1(n3380), .A2(\registers[25][22] ), .B1(n3377), .B2(
        \registers[24][22] ), .ZN(n2377) );
  AOI22_X1 U1761 ( .A1(n3380), .A2(\registers[25][23] ), .B1(n3377), .B2(
        \registers[24][23] ), .ZN(n2360) );
  AOI22_X1 U1762 ( .A1(n3380), .A2(\registers[25][24] ), .B1(n3377), .B2(
        \registers[24][24] ), .ZN(n2343) );
  AOI22_X1 U1763 ( .A1(n3380), .A2(\registers[25][25] ), .B1(n3377), .B2(
        \registers[24][25] ), .ZN(n2326) );
  AOI22_X1 U1764 ( .A1(n3380), .A2(\registers[25][26] ), .B1(n3377), .B2(
        \registers[24][26] ), .ZN(n2309) );
  AOI22_X1 U1765 ( .A1(n3380), .A2(\registers[25][27] ), .B1(n3377), .B2(
        \registers[24][27] ), .ZN(n2292) );
  AOI22_X1 U1766 ( .A1(n3380), .A2(\registers[25][28] ), .B1(n3377), .B2(
        \registers[24][28] ), .ZN(n2275) );
  AOI22_X1 U1767 ( .A1(n3380), .A2(\registers[25][29] ), .B1(n3377), .B2(
        \registers[24][29] ), .ZN(n2258) );
  AOI22_X1 U1768 ( .A1(n3380), .A2(\registers[25][30] ), .B1(n3377), .B2(
        \registers[24][30] ), .ZN(n2241) );
  AOI22_X1 U1769 ( .A1(n3380), .A2(\registers[25][31] ), .B1(n3377), .B2(
        \registers[24][31] ), .ZN(n2203) );
  AOI22_X1 U1770 ( .A1(n3465), .A2(\registers[25][0] ), .B1(n3462), .B2(
        \registers[24][0] ), .ZN(n2167) );
  AOI22_X1 U1771 ( .A1(n3465), .A2(\registers[25][1] ), .B1(n3462), .B2(
        \registers[24][1] ), .ZN(n2143) );
  AOI22_X1 U1772 ( .A1(n3465), .A2(\registers[25][2] ), .B1(n3462), .B2(
        \registers[24][2] ), .ZN(n2126) );
  AOI22_X1 U1773 ( .A1(n3465), .A2(\registers[25][3] ), .B1(n3462), .B2(
        \registers[24][3] ), .ZN(n2109) );
  AOI22_X1 U1774 ( .A1(n3465), .A2(\registers[25][4] ), .B1(n3462), .B2(
        \registers[24][4] ), .ZN(n2092) );
  AOI22_X1 U1775 ( .A1(n3465), .A2(\registers[25][5] ), .B1(n3462), .B2(
        \registers[24][5] ), .ZN(n2075) );
  AOI22_X1 U1776 ( .A1(n3465), .A2(\registers[25][6] ), .B1(n3462), .B2(
        \registers[24][6] ), .ZN(n2058) );
  AOI22_X1 U1777 ( .A1(n3465), .A2(\registers[25][7] ), .B1(n3462), .B2(
        \registers[24][7] ), .ZN(n2041) );
  AOI22_X1 U1778 ( .A1(n3465), .A2(\registers[25][8] ), .B1(n3462), .B2(
        \registers[24][8] ), .ZN(n2024) );
  AOI22_X1 U1779 ( .A1(n3465), .A2(\registers[25][9] ), .B1(n3462), .B2(
        \registers[24][9] ), .ZN(n2007) );
  AOI22_X1 U1780 ( .A1(n3465), .A2(\registers[25][10] ), .B1(n3462), .B2(
        \registers[24][10] ), .ZN(n1990) );
  AOI22_X1 U1781 ( .A1(n3466), .A2(\registers[25][11] ), .B1(n3463), .B2(
        \registers[24][11] ), .ZN(n1973) );
  AOI22_X1 U1782 ( .A1(n3466), .A2(\registers[25][12] ), .B1(n3463), .B2(
        \registers[24][12] ), .ZN(n1956) );
  AOI22_X1 U1783 ( .A1(n3466), .A2(\registers[25][13] ), .B1(n3463), .B2(
        \registers[24][13] ), .ZN(n1939) );
  AOI22_X1 U1784 ( .A1(n3466), .A2(\registers[25][14] ), .B1(n3463), .B2(
        \registers[24][14] ), .ZN(n1922) );
  AOI22_X1 U1785 ( .A1(n3466), .A2(\registers[25][15] ), .B1(n3463), .B2(
        \registers[24][15] ), .ZN(n1905) );
  AOI22_X1 U1786 ( .A1(n3466), .A2(\registers[25][16] ), .B1(n3463), .B2(
        \registers[24][16] ), .ZN(n1888) );
  AOI22_X1 U1787 ( .A1(n3466), .A2(\registers[25][17] ), .B1(n3463), .B2(
        \registers[24][17] ), .ZN(n1871) );
  AOI22_X1 U1788 ( .A1(n3466), .A2(\registers[25][18] ), .B1(n3463), .B2(
        \registers[24][18] ), .ZN(n1854) );
  AOI22_X1 U1789 ( .A1(n3466), .A2(\registers[25][19] ), .B1(n3463), .B2(
        \registers[24][19] ), .ZN(n1837) );
  AOI22_X1 U1790 ( .A1(n3466), .A2(\registers[25][20] ), .B1(n3463), .B2(
        \registers[24][20] ), .ZN(n1820) );
  AOI22_X1 U1791 ( .A1(n3466), .A2(\registers[25][21] ), .B1(n3463), .B2(
        \registers[24][21] ), .ZN(n1803) );
  AOI22_X1 U1792 ( .A1(n3378), .A2(\registers[25][0] ), .B1(n3375), .B2(
        \registers[24][0] ), .ZN(n2758) );
  AOI22_X1 U1793 ( .A1(n3378), .A2(\registers[25][1] ), .B1(n3375), .B2(
        \registers[24][1] ), .ZN(n2734) );
  AOI22_X1 U1794 ( .A1(n3378), .A2(\registers[25][2] ), .B1(n3375), .B2(
        \registers[24][2] ), .ZN(n2717) );
  AOI22_X1 U1795 ( .A1(n3378), .A2(\registers[25][3] ), .B1(n3375), .B2(
        \registers[24][3] ), .ZN(n2700) );
  AOI22_X1 U1796 ( .A1(n3378), .A2(\registers[25][4] ), .B1(n3375), .B2(
        \registers[24][4] ), .ZN(n2683) );
  AOI22_X1 U1797 ( .A1(n3378), .A2(\registers[25][5] ), .B1(n3375), .B2(
        \registers[24][5] ), .ZN(n2666) );
  AOI22_X1 U1798 ( .A1(n3378), .A2(\registers[25][6] ), .B1(n3375), .B2(
        \registers[24][6] ), .ZN(n2649) );
  AOI22_X1 U1799 ( .A1(n3378), .A2(\registers[25][7] ), .B1(n3375), .B2(
        \registers[24][7] ), .ZN(n2632) );
  AOI22_X1 U1800 ( .A1(n3378), .A2(\registers[25][8] ), .B1(n3375), .B2(
        \registers[24][8] ), .ZN(n2615) );
  AOI22_X1 U1801 ( .A1(n3378), .A2(\registers[25][9] ), .B1(n3375), .B2(
        \registers[24][9] ), .ZN(n2598) );
  AOI22_X1 U1802 ( .A1(n3378), .A2(\registers[25][10] ), .B1(n3375), .B2(
        \registers[24][10] ), .ZN(n2581) );
  AOI22_X1 U1803 ( .A1(n3379), .A2(\registers[25][11] ), .B1(n3376), .B2(
        \registers[24][11] ), .ZN(n2564) );
  AOI22_X1 U1804 ( .A1(n3379), .A2(\registers[25][12] ), .B1(n3376), .B2(
        \registers[24][12] ), .ZN(n2547) );
  AOI22_X1 U1805 ( .A1(n3379), .A2(\registers[25][13] ), .B1(n3376), .B2(
        \registers[24][13] ), .ZN(n2530) );
  AOI22_X1 U1806 ( .A1(n3379), .A2(\registers[25][14] ), .B1(n3376), .B2(
        \registers[24][14] ), .ZN(n2513) );
  AOI22_X1 U1807 ( .A1(n3379), .A2(\registers[25][15] ), .B1(n3376), .B2(
        \registers[24][15] ), .ZN(n2496) );
  AOI22_X1 U1808 ( .A1(n3379), .A2(\registers[25][16] ), .B1(n3376), .B2(
        \registers[24][16] ), .ZN(n2479) );
  AOI22_X1 U1809 ( .A1(n3379), .A2(\registers[25][17] ), .B1(n3376), .B2(
        \registers[24][17] ), .ZN(n2462) );
  AOI22_X1 U1810 ( .A1(n3379), .A2(\registers[25][18] ), .B1(n3376), .B2(
        \registers[24][18] ), .ZN(n2445) );
  AOI22_X1 U1811 ( .A1(n3379), .A2(\registers[25][19] ), .B1(n3376), .B2(
        \registers[24][19] ), .ZN(n2428) );
  AOI22_X1 U1812 ( .A1(n3379), .A2(\registers[25][20] ), .B1(n3376), .B2(
        \registers[24][20] ), .ZN(n2411) );
  AOI22_X1 U1813 ( .A1(n3379), .A2(\registers[25][21] ), .B1(n3376), .B2(
        \registers[24][21] ), .ZN(n2394) );
  AOI22_X1 U1814 ( .A1(n3455), .A2(\registers[29][22] ), .B1(n3452), .B2(
        \registers[28][22] ), .ZN(n1787) );
  AOI22_X1 U1815 ( .A1(n3455), .A2(\registers[29][23] ), .B1(n3452), .B2(
        \registers[28][23] ), .ZN(n1770) );
  AOI22_X1 U1816 ( .A1(n3455), .A2(\registers[29][24] ), .B1(n3452), .B2(
        \registers[28][24] ), .ZN(n1753) );
  AOI22_X1 U1817 ( .A1(n3455), .A2(\registers[29][25] ), .B1(n3452), .B2(
        \registers[28][25] ), .ZN(n1736) );
  AOI22_X1 U1818 ( .A1(n3455), .A2(\registers[29][26] ), .B1(n3452), .B2(
        \registers[28][26] ), .ZN(n1719) );
  AOI22_X1 U1819 ( .A1(n3455), .A2(\registers[29][27] ), .B1(n3452), .B2(
        \registers[28][27] ), .ZN(n1702) );
  AOI22_X1 U1820 ( .A1(n3455), .A2(\registers[29][28] ), .B1(n3452), .B2(
        \registers[28][28] ), .ZN(n1685) );
  AOI22_X1 U1821 ( .A1(n3455), .A2(\registers[29][29] ), .B1(n3452), .B2(
        \registers[28][29] ), .ZN(n1668) );
  AOI22_X1 U1822 ( .A1(n3455), .A2(\registers[29][30] ), .B1(n3452), .B2(
        \registers[28][30] ), .ZN(n1651) );
  AOI22_X1 U1823 ( .A1(n3455), .A2(\registers[29][31] ), .B1(n3452), .B2(
        \registers[28][31] ), .ZN(n1617) );
  AOI22_X1 U1824 ( .A1(n3368), .A2(\registers[29][22] ), .B1(n3365), .B2(
        \registers[28][22] ), .ZN(n2378) );
  AOI22_X1 U1825 ( .A1(n3368), .A2(\registers[29][23] ), .B1(n3365), .B2(
        \registers[28][23] ), .ZN(n2361) );
  AOI22_X1 U1826 ( .A1(n3368), .A2(\registers[29][24] ), .B1(n3365), .B2(
        \registers[28][24] ), .ZN(n2344) );
  AOI22_X1 U1827 ( .A1(n3368), .A2(\registers[29][25] ), .B1(n3365), .B2(
        \registers[28][25] ), .ZN(n2327) );
  AOI22_X1 U1828 ( .A1(n3368), .A2(\registers[29][26] ), .B1(n3365), .B2(
        \registers[28][26] ), .ZN(n2310) );
  AOI22_X1 U1829 ( .A1(n3368), .A2(\registers[29][27] ), .B1(n3365), .B2(
        \registers[28][27] ), .ZN(n2293) );
  AOI22_X1 U1830 ( .A1(n3368), .A2(\registers[29][28] ), .B1(n3365), .B2(
        \registers[28][28] ), .ZN(n2276) );
  AOI22_X1 U1831 ( .A1(n3368), .A2(\registers[29][29] ), .B1(n3365), .B2(
        \registers[28][29] ), .ZN(n2259) );
  AOI22_X1 U1832 ( .A1(n3368), .A2(\registers[29][30] ), .B1(n3365), .B2(
        \registers[28][30] ), .ZN(n2242) );
  AOI22_X1 U1833 ( .A1(n3368), .A2(\registers[29][31] ), .B1(n3365), .B2(
        \registers[28][31] ), .ZN(n2208) );
  AOI22_X1 U1834 ( .A1(n3453), .A2(\registers[29][0] ), .B1(n3450), .B2(
        \registers[28][0] ), .ZN(n2170) );
  AOI22_X1 U1835 ( .A1(n3453), .A2(\registers[29][1] ), .B1(n3450), .B2(
        \registers[28][1] ), .ZN(n2144) );
  AOI22_X1 U1836 ( .A1(n3453), .A2(\registers[29][2] ), .B1(n3450), .B2(
        \registers[28][2] ), .ZN(n2127) );
  AOI22_X1 U1837 ( .A1(n3453), .A2(\registers[29][3] ), .B1(n3450), .B2(
        \registers[28][3] ), .ZN(n2110) );
  AOI22_X1 U1838 ( .A1(n3453), .A2(\registers[29][4] ), .B1(n3450), .B2(
        \registers[28][4] ), .ZN(n2093) );
  AOI22_X1 U1839 ( .A1(n3453), .A2(\registers[29][5] ), .B1(n3450), .B2(
        \registers[28][5] ), .ZN(n2076) );
  AOI22_X1 U1840 ( .A1(n3453), .A2(\registers[29][6] ), .B1(n3450), .B2(
        \registers[28][6] ), .ZN(n2059) );
  AOI22_X1 U1841 ( .A1(n3453), .A2(\registers[29][7] ), .B1(n3450), .B2(
        \registers[28][7] ), .ZN(n2042) );
  AOI22_X1 U1842 ( .A1(n3453), .A2(\registers[29][8] ), .B1(n3450), .B2(
        \registers[28][8] ), .ZN(n2025) );
  AOI22_X1 U1843 ( .A1(n3453), .A2(\registers[29][9] ), .B1(n3450), .B2(
        \registers[28][9] ), .ZN(n2008) );
  AOI22_X1 U1844 ( .A1(n3453), .A2(\registers[29][10] ), .B1(n3450), .B2(
        \registers[28][10] ), .ZN(n1991) );
  AOI22_X1 U1845 ( .A1(n3454), .A2(\registers[29][11] ), .B1(n3451), .B2(
        \registers[28][11] ), .ZN(n1974) );
  AOI22_X1 U1846 ( .A1(n3454), .A2(\registers[29][12] ), .B1(n3451), .B2(
        \registers[28][12] ), .ZN(n1957) );
  AOI22_X1 U1847 ( .A1(n3454), .A2(\registers[29][13] ), .B1(n3451), .B2(
        \registers[28][13] ), .ZN(n1940) );
  AOI22_X1 U1848 ( .A1(n3454), .A2(\registers[29][14] ), .B1(n3451), .B2(
        \registers[28][14] ), .ZN(n1923) );
  AOI22_X1 U1849 ( .A1(n3454), .A2(\registers[29][15] ), .B1(n3451), .B2(
        \registers[28][15] ), .ZN(n1906) );
  AOI22_X1 U1850 ( .A1(n3454), .A2(\registers[29][16] ), .B1(n3451), .B2(
        \registers[28][16] ), .ZN(n1889) );
  AOI22_X1 U1851 ( .A1(n3454), .A2(\registers[29][17] ), .B1(n3451), .B2(
        \registers[28][17] ), .ZN(n1872) );
  AOI22_X1 U1852 ( .A1(n3454), .A2(\registers[29][18] ), .B1(n3451), .B2(
        \registers[28][18] ), .ZN(n1855) );
  AOI22_X1 U1853 ( .A1(n3454), .A2(\registers[29][19] ), .B1(n3451), .B2(
        \registers[28][19] ), .ZN(n1838) );
  AOI22_X1 U1854 ( .A1(n3454), .A2(\registers[29][20] ), .B1(n3451), .B2(
        \registers[28][20] ), .ZN(n1821) );
  AOI22_X1 U1855 ( .A1(n3454), .A2(\registers[29][21] ), .B1(n3451), .B2(
        \registers[28][21] ), .ZN(n1804) );
  AOI22_X1 U1856 ( .A1(n3366), .A2(\registers[29][0] ), .B1(n3363), .B2(
        \registers[28][0] ), .ZN(n2761) );
  AOI22_X1 U1857 ( .A1(n3366), .A2(\registers[29][1] ), .B1(n3363), .B2(
        \registers[28][1] ), .ZN(n2735) );
  AOI22_X1 U1858 ( .A1(n3366), .A2(\registers[29][2] ), .B1(n3363), .B2(
        \registers[28][2] ), .ZN(n2718) );
  AOI22_X1 U1859 ( .A1(n3366), .A2(\registers[29][3] ), .B1(n3363), .B2(
        \registers[28][3] ), .ZN(n2701) );
  AOI22_X1 U1860 ( .A1(n3366), .A2(\registers[29][4] ), .B1(n3363), .B2(
        \registers[28][4] ), .ZN(n2684) );
  AOI22_X1 U1861 ( .A1(n3366), .A2(\registers[29][5] ), .B1(n3363), .B2(
        \registers[28][5] ), .ZN(n2667) );
  AOI22_X1 U1862 ( .A1(n3366), .A2(\registers[29][6] ), .B1(n3363), .B2(
        \registers[28][6] ), .ZN(n2650) );
  AOI22_X1 U1863 ( .A1(n3366), .A2(\registers[29][7] ), .B1(n3363), .B2(
        \registers[28][7] ), .ZN(n2633) );
  AOI22_X1 U1864 ( .A1(n3366), .A2(\registers[29][8] ), .B1(n3363), .B2(
        \registers[28][8] ), .ZN(n2616) );
  AOI22_X1 U1865 ( .A1(n3366), .A2(\registers[29][9] ), .B1(n3363), .B2(
        \registers[28][9] ), .ZN(n2599) );
  AOI22_X1 U1866 ( .A1(n3366), .A2(\registers[29][10] ), .B1(n3363), .B2(
        \registers[28][10] ), .ZN(n2582) );
  AOI22_X1 U1867 ( .A1(n3367), .A2(\registers[29][11] ), .B1(n3364), .B2(
        \registers[28][11] ), .ZN(n2565) );
  AOI22_X1 U1868 ( .A1(n3367), .A2(\registers[29][12] ), .B1(n3364), .B2(
        \registers[28][12] ), .ZN(n2548) );
  AOI22_X1 U1869 ( .A1(n3367), .A2(\registers[29][13] ), .B1(n3364), .B2(
        \registers[28][13] ), .ZN(n2531) );
  AOI22_X1 U1870 ( .A1(n3367), .A2(\registers[29][14] ), .B1(n3364), .B2(
        \registers[28][14] ), .ZN(n2514) );
  AOI22_X1 U1871 ( .A1(n3367), .A2(\registers[29][15] ), .B1(n3364), .B2(
        \registers[28][15] ), .ZN(n2497) );
  AOI22_X1 U1872 ( .A1(n3367), .A2(\registers[29][16] ), .B1(n3364), .B2(
        \registers[28][16] ), .ZN(n2480) );
  AOI22_X1 U1873 ( .A1(n3367), .A2(\registers[29][17] ), .B1(n3364), .B2(
        \registers[28][17] ), .ZN(n2463) );
  AOI22_X1 U1874 ( .A1(n3367), .A2(\registers[29][18] ), .B1(n3364), .B2(
        \registers[28][18] ), .ZN(n2446) );
  AOI22_X1 U1875 ( .A1(n3367), .A2(\registers[29][19] ), .B1(n3364), .B2(
        \registers[28][19] ), .ZN(n2429) );
  AOI22_X1 U1876 ( .A1(n3367), .A2(\registers[29][20] ), .B1(n3364), .B2(
        \registers[28][20] ), .ZN(n2412) );
  AOI22_X1 U1877 ( .A1(n3367), .A2(\registers[29][21] ), .B1(n3364), .B2(
        \registers[28][21] ), .ZN(n2395) );
  OAI22_X1 U1878 ( .A1(n713), .A2(n4259), .B1(n718), .B2(n980), .ZN(n2786) );
  OAI22_X1 U1879 ( .A1(n598), .A2(n713), .B1(n718), .B2(n979), .ZN(n2787) );
  OAI22_X1 U1880 ( .A1(n716), .A2(n696), .B1(n719), .B2(n978), .ZN(n2788) );
  OAI22_X1 U1881 ( .A1(n714), .A2(n729), .B1(n720), .B2(n977), .ZN(n2789) );
  OAI22_X1 U1882 ( .A1(n715), .A2(n4256), .B1(n724), .B2(n976), .ZN(n2790) );
  OAI22_X1 U1883 ( .A1(n716), .A2(n4255), .B1(n721), .B2(n975), .ZN(n2791) );
  OAI22_X1 U1884 ( .A1(n4254), .A2(n714), .B1(n722), .B2(n974), .ZN(n2792) );
  OAI22_X1 U1885 ( .A1(n717), .A2(n745), .B1(n723), .B2(n973), .ZN(n2793) );
  OAI22_X1 U1886 ( .A1(n717), .A2(n208), .B1(n718), .B2(n972), .ZN(n2794) );
  OAI22_X1 U1887 ( .A1(n186), .A2(n717), .B1(n720), .B2(n971), .ZN(n2795) );
  OAI22_X1 U1888 ( .A1(n700), .A2(n714), .B1(n721), .B2(n970), .ZN(n2796) );
  OAI22_X1 U1889 ( .A1(n698), .A2(n715), .B1(n724), .B2(n969), .ZN(n2797) );
  OAI22_X1 U1890 ( .A1(n716), .A2(n4249), .B1(n723), .B2(n968), .ZN(n2798) );
  OAI22_X1 U1891 ( .A1(n716), .A2(n706), .B1(n725), .B2(n967), .ZN(n2799) );
  OAI22_X1 U1892 ( .A1(n713), .A2(n4247), .B1(n718), .B2(n966), .ZN(n2800) );
  OAI22_X1 U1893 ( .A1(n717), .A2(n4246), .B1(n720), .B2(n965), .ZN(n2801) );
  OAI22_X1 U1894 ( .A1(net39055), .A2(n713), .B1(n719), .B2(n964), .ZN(n2802)
         );
  OAI22_X1 U1895 ( .A1(n714), .A2(n742), .B1(n720), .B2(n963), .ZN(n2803) );
  OAI22_X1 U1896 ( .A1(n270), .A2(n715), .B1(n724), .B2(n962), .ZN(n2804) );
  OAI22_X1 U1897 ( .A1(n674), .A2(n713), .B1(n719), .B2(n982), .ZN(n2784) );
  OAI22_X1 U1898 ( .A1(n714), .A2(n4260), .B1(n719), .B2(n981), .ZN(n2785) );
  OAI22_X1 U1899 ( .A1(n716), .A2(n263), .B1(n721), .B2(n961), .ZN(n2805) );
  OAI22_X1 U1900 ( .A1(n3615), .A2(n4263), .B1(n3621), .B2(n856), .ZN(n2846)
         );
  OAI22_X1 U1901 ( .A1(n4262), .A2(n3615), .B1(n3621), .B2(n855), .ZN(n2847)
         );
  OAI22_X1 U1902 ( .A1(n201), .A2(n3606), .B1(n3609), .B2(n824), .ZN(n2878) );
  OAI22_X1 U1903 ( .A1(n179), .A2(n3606), .B1(n3609), .B2(n823), .ZN(n2879) );
  OAI22_X1 U1904 ( .A1(n730), .A2(n371), .B1(n381), .B2(n664), .ZN(n2910) );
  OAI22_X1 U1905 ( .A1(n179), .A2(n372), .B1(n377), .B2(n663), .ZN(n2911) );
  OAI22_X1 U1906 ( .A1(n730), .A2(n755), .B1(n754), .B2(n632), .ZN(n2942) );
  OAI22_X1 U1907 ( .A1(n4262), .A2(n756), .B1(n753), .B2(n631), .ZN(n2943) );
  OAI22_X1 U1908 ( .A1(n201), .A2(n995), .B1(n905), .B2(n504), .ZN(n3006) );
  OAI22_X1 U1909 ( .A1(n179), .A2(n996), .B1(n905), .B2(n503), .ZN(n3007) );
  OAI22_X1 U1910 ( .A1(n201), .A2(n1035), .B1(n192), .B2(n472), .ZN(n3038) );
  OAI22_X1 U1911 ( .A1(n601), .A2(n1036), .B1(n233), .B2(n471), .ZN(n3039) );
  OAI22_X1 U1912 ( .A1(n4263), .A2(net44474), .B1(net26421), .B2(n440), .ZN(
        n3070) );
  OAI22_X1 U1913 ( .A1(n600), .A2(net26413), .B1(net26421), .B2(n439), .ZN(
        n3071) );
  OAI22_X1 U1914 ( .A1(n4263), .A2(n3302), .B1(n3291), .B2(n344), .ZN(n3102)
         );
  OAI22_X1 U1915 ( .A1(n601), .A2(n3303), .B1(n3534), .B2(n343), .ZN(n3103) );
  OAI22_X1 U1916 ( .A1(n201), .A2(n1143), .B1(n1050), .B2(n312), .ZN(n3134) );
  OAI22_X1 U1917 ( .A1(n4262), .A2(n1201), .B1(n1057), .B2(n311), .ZN(n3135)
         );
  OAI22_X1 U1918 ( .A1(n730), .A2(n580), .B1(n583), .B2(n88), .ZN(n3230) );
  OAI22_X1 U1919 ( .A1(n601), .A2(n580), .B1(n589), .B2(n87), .ZN(n3231) );
  OAI22_X1 U1920 ( .A1(n4263), .A2(n565), .B1(n568), .B2(n56), .ZN(n3262) );
  OAI22_X1 U1921 ( .A1(n4262), .A2(n565), .B1(n573), .B2(n55), .ZN(n3263) );
  OAI22_X1 U1922 ( .A1(n4258), .A2(n1039), .B1(n192), .B2(n467), .ZN(n3043) );
  OAI22_X1 U1923 ( .A1(n18), .A2(n1041), .B1(n192), .B2(n465), .ZN(n3045) );
  OAI22_X1 U1924 ( .A1(n1035), .A2(n402), .B1(n1045), .B2(n463), .ZN(n3047) );
  OAI22_X1 U1925 ( .A1(n745), .A2(n1034), .B1(n232), .B2(n461), .ZN(n3049) );
  OAI22_X1 U1926 ( .A1(n178), .A2(n1038), .B1(n1045), .B2(n470), .ZN(n3040) );
  OAI22_X1 U1927 ( .A1(n195), .A2(n1037), .B1(n1045), .B2(n469), .ZN(n3041) );
  OAI22_X1 U1928 ( .A1(n546), .A2(n1032), .B1(n1046), .B2(n474), .ZN(n3036) );
  OAI22_X1 U1929 ( .A1(n732), .A2(n1029), .B1(n1044), .B2(n477), .ZN(n3033) );
  OAI22_X1 U1930 ( .A1(n275), .A2(n1030), .B1(n1046), .B2(n476), .ZN(n3034) );
  OAI22_X1 U1931 ( .A1(n1), .A2(n1031), .B1(n1046), .B2(n475), .ZN(n3035) );
  OAI22_X1 U1932 ( .A1(n715), .A2(n4263), .B1(n722), .B2(n984), .ZN(n2782) );
  OAI22_X1 U1933 ( .A1(n600), .A2(n715), .B1(n723), .B2(n983), .ZN(n2783) );
  OAI22_X1 U1934 ( .A1(n717), .A2(n606), .B1(n725), .B2(n992), .ZN(n2774) );
  OAI22_X1 U1935 ( .A1(n608), .A2(n714), .B1(n721), .B2(n991), .ZN(n2775) );
  OAI22_X1 U1936 ( .A1(n715), .A2(n268), .B1(n722), .B2(n990), .ZN(n2776) );
  OAI22_X1 U1937 ( .A1(n546), .A2(n713), .B1(n723), .B2(n986), .ZN(n2780) );
  OAI22_X1 U1938 ( .A1(n716), .A2(n4264), .B1(n725), .B2(n985), .ZN(n2781) );
  OAI22_X1 U1939 ( .A1(n713), .A2(n238), .B1(n724), .B2(n989), .ZN(n2777) );
  OAI22_X1 U1940 ( .A1(n714), .A2(n4267), .B1(n722), .B2(n988), .ZN(n2778) );
  OAI22_X1 U1941 ( .A1(n717), .A2(n4266), .B1(n725), .B2(n987), .ZN(n2779) );
  OAI22_X1 U1942 ( .A1(n606), .A2(n562), .B1(n3617), .B2(n864), .ZN(n2838) );
  OAI22_X1 U1943 ( .A1(n4270), .A2(n561), .B1(n3618), .B2(n863), .ZN(n2839) );
  OAI22_X1 U1944 ( .A1(n4269), .A2(n3616), .B1(n3621), .B2(n862), .ZN(n2840)
         );
  OAI22_X1 U1945 ( .A1(n606), .A2(n370), .B1(n382), .B2(n672), .ZN(n2902) );
  OAI22_X1 U1946 ( .A1(n608), .A2(n371), .B1(n375), .B2(n671), .ZN(n2903) );
  OAI22_X1 U1947 ( .A1(n194), .A2(n371), .B1(n383), .B2(n670), .ZN(n2904) );
  OAI22_X1 U1948 ( .A1(n4271), .A2(n288), .B1(n362), .B2(n160), .ZN(n3158) );
  OAI22_X1 U1949 ( .A1(n608), .A2(n353), .B1(n358), .B2(n159), .ZN(n3159) );
  OAI22_X1 U1950 ( .A1(n733), .A2(n353), .B1(n368), .B2(n158), .ZN(n3160) );
  OAI22_X1 U1951 ( .A1(n21), .A2(n3615), .B1(n3621), .B2(n852), .ZN(n2850) );
  OAI22_X1 U1952 ( .A1(n4258), .A2(n3615), .B1(n3620), .B2(n851), .ZN(n2851)
         );
  OAI22_X1 U1953 ( .A1(n696), .A2(n3615), .B1(n3618), .B2(n850), .ZN(n2852) );
  OAI22_X1 U1954 ( .A1(n188), .A2(n3615), .B1(n3620), .B2(n849), .ZN(n2853) );
  OAI22_X1 U1955 ( .A1(n4256), .A2(n3615), .B1(n3618), .B2(n848), .ZN(n2854)
         );
  OAI22_X1 U1956 ( .A1(n3614), .A2(n4255), .B1(n3617), .B2(n847), .ZN(n2855)
         );
  OAI22_X1 U1957 ( .A1(n4254), .A2(n562), .B1(n3619), .B2(n846), .ZN(n2856) );
  OAI22_X1 U1958 ( .A1(n745), .A2(n561), .B1(n3618), .B2(n845), .ZN(n2857) );
  OAI22_X1 U1959 ( .A1(n396), .A2(n562), .B1(n3618), .B2(n844), .ZN(n2858) );
  OAI22_X1 U1960 ( .A1(n186), .A2(n561), .B1(n3617), .B2(n843), .ZN(n2859) );
  OAI22_X1 U1961 ( .A1(n700), .A2(n3616), .B1(n3619), .B2(n842), .ZN(n2860) );
  OAI22_X1 U1962 ( .A1(n697), .A2(n3614), .B1(n3620), .B2(n841), .ZN(n2861) );
  OAI22_X1 U1963 ( .A1(n4249), .A2(n562), .B1(n3621), .B2(n840), .ZN(n2862) );
  OAI22_X1 U1964 ( .A1(n561), .A2(n184), .B1(n3617), .B2(n839), .ZN(n2863) );
  OAI22_X1 U1965 ( .A1(n3616), .A2(n4247), .B1(n3619), .B2(n838), .ZN(n2864)
         );
  OAI22_X1 U1966 ( .A1(n3614), .A2(n4246), .B1(n3621), .B2(n837), .ZN(n2865)
         );
  OAI22_X1 U1967 ( .A1(net39055), .A2(n562), .B1(n3621), .B2(n836), .ZN(n2866)
         );
  OAI22_X1 U1968 ( .A1(n4245), .A2(n561), .B1(n3620), .B2(n835), .ZN(n2867) );
  OAI22_X1 U1969 ( .A1(n399), .A2(n3616), .B1(n3618), .B2(n834), .ZN(n2868) );
  OAI22_X1 U1970 ( .A1(n181), .A2(n372), .B1(n380), .B2(n660), .ZN(n2914) );
  OAI22_X1 U1971 ( .A1(n177), .A2(n370), .B1(n377), .B2(n659), .ZN(n2915) );
  OAI22_X1 U1972 ( .A1(n4257), .A2(n371), .B1(n384), .B2(n658), .ZN(n2916) );
  OAI22_X1 U1973 ( .A1(n180), .A2(n372), .B1(n381), .B2(n657), .ZN(n2917) );
  OAI22_X1 U1974 ( .A1(n552), .A2(n371), .B1(n376), .B2(n656), .ZN(n2918) );
  OAI22_X1 U1975 ( .A1(n402), .A2(n371), .B1(n377), .B2(n655), .ZN(n2919) );
  OAI22_X1 U1976 ( .A1(n415), .A2(n371), .B1(n376), .B2(n654), .ZN(n2920) );
  OAI22_X1 U1977 ( .A1(n260), .A2(n370), .B1(n376), .B2(n653), .ZN(n2921) );
  OAI22_X1 U1978 ( .A1(n186), .A2(n371), .B1(n382), .B2(n651), .ZN(n2923) );
  OAI22_X1 U1979 ( .A1(n699), .A2(n370), .B1(n384), .B2(n650), .ZN(n2924) );
  OAI22_X1 U1980 ( .A1(n224), .A2(n370), .B1(n378), .B2(n649), .ZN(n2925) );
  OAI22_X1 U1981 ( .A1(n744), .A2(n370), .B1(n374), .B2(n648), .ZN(n2926) );
  OAI22_X1 U1982 ( .A1(n28), .A2(n370), .B1(n377), .B2(n647), .ZN(n2927) );
  OAI22_X1 U1983 ( .A1(n592), .A2(n372), .B1(n383), .B2(n646), .ZN(n2928) );
  OAI22_X1 U1984 ( .A1(n594), .A2(n370), .B1(n378), .B2(n645), .ZN(n2929) );
  OAI22_X1 U1985 ( .A1(n197), .A2(n372), .B1(n374), .B2(n644), .ZN(n2930) );
  OAI22_X1 U1986 ( .A1(n5), .A2(n371), .B1(n381), .B2(n643), .ZN(n2931) );
  OAI22_X1 U1987 ( .A1(n4244), .A2(n372), .B1(n378), .B2(n642), .ZN(n2932) );
  OAI22_X1 U1988 ( .A1(n4252), .A2(n1027), .B1(n1005), .B2(n524), .ZN(n2986)
         );
  OAI22_X1 U1989 ( .A1(n709), .A2(n1021), .B1(n1006), .B2(n523), .ZN(n2987) );
  OAI22_X1 U1990 ( .A1(n183), .A2(n1022), .B1(n1007), .B2(n522), .ZN(n2988) );
  OAI22_X1 U1991 ( .A1(n224), .A2(n1025), .B1(n1016), .B2(n521), .ZN(n2989) );
  OAI22_X1 U1992 ( .A1(n280), .A2(n1024), .B1(n1007), .B2(n520), .ZN(n2990) );
  OAI22_X1 U1993 ( .A1(n707), .A2(n1026), .B1(n1016), .B2(n519), .ZN(n2991) );
  OAI22_X1 U1994 ( .A1(n1021), .A2(n735), .B1(n1016), .B2(n518), .ZN(n2992) );
  OAI22_X1 U1995 ( .A1(n1022), .A2(n734), .B1(n1016), .B2(n517), .ZN(n2993) );
  OAI22_X1 U1996 ( .A1(net44818), .A2(n1023), .B1(n1016), .B2(n516), .ZN(n2994) );
  OAI22_X1 U1997 ( .A1(n5), .A2(n1028), .B1(n1017), .B2(n515), .ZN(n2995) );
  OAI22_X1 U1998 ( .A1(n4244), .A2(n1023), .B1(n1005), .B2(n514), .ZN(n2996)
         );
  OAI22_X1 U1999 ( .A1(n740), .A2(n353), .B1(n366), .B2(n148), .ZN(n3170) );
  OAI22_X1 U2000 ( .A1(n599), .A2(n354), .B1(n360), .B2(n147), .ZN(n3171) );
  OAI22_X1 U2001 ( .A1(n4257), .A2(n354), .B1(n365), .B2(n146), .ZN(n3172) );
  OAI22_X1 U2002 ( .A1(n728), .A2(n288), .B1(n360), .B2(n145), .ZN(n3173) );
  OAI22_X1 U2003 ( .A1(n552), .A2(n353), .B1(n369), .B2(n144), .ZN(n3174) );
  OAI22_X1 U2004 ( .A1(n739), .A2(n354), .B1(n366), .B2(n143), .ZN(n3175) );
  OAI22_X1 U2005 ( .A1(n415), .A2(n353), .B1(n359), .B2(n142), .ZN(n3176) );
  OAI22_X1 U2006 ( .A1(n260), .A2(n353), .B1(n360), .B2(n141), .ZN(n3177) );
  OAI22_X1 U2007 ( .A1(n701), .A2(n353), .B1(n361), .B2(n140), .ZN(n3178) );
  OAI22_X1 U2008 ( .A1(n708), .A2(n288), .B1(n357), .B2(n139), .ZN(n3179) );
  OAI22_X1 U2009 ( .A1(n4251), .A2(n288), .B1(n362), .B2(n138), .ZN(n3180) );
  OAI22_X1 U2010 ( .A1(n697), .A2(n288), .B1(n367), .B2(n137), .ZN(n3181) );
  OAI22_X1 U2011 ( .A1(n744), .A2(n288), .B1(n369), .B2(n136), .ZN(n3182) );
  OAI22_X1 U2012 ( .A1(n706), .A2(n354), .B1(n365), .B2(n135), .ZN(n3183) );
  OAI22_X1 U2013 ( .A1(n735), .A2(n288), .B1(n358), .B2(n134), .ZN(n3184) );
  OAI22_X1 U2014 ( .A1(n593), .A2(n354), .B1(n358), .B2(n133), .ZN(n3185) );
  OAI22_X1 U2015 ( .A1(net39055), .A2(n353), .B1(n362), .B2(n132), .ZN(n3186)
         );
  OAI22_X1 U2016 ( .A1(n4245), .A2(n288), .B1(n368), .B2(n131), .ZN(n3187) );
  OAI22_X1 U2017 ( .A1(n4244), .A2(n354), .B1(n361), .B2(n130), .ZN(n3188) );
  OAI22_X1 U2018 ( .A1(n178), .A2(n3616), .B1(n3619), .B2(n854), .ZN(n2848) );
  OAI22_X1 U2019 ( .A1(n575), .A2(n3614), .B1(n3617), .B2(n853), .ZN(n2849) );
  OAI22_X1 U2020 ( .A1(n674), .A2(n371), .B1(n381), .B2(n662), .ZN(n2912) );
  OAI22_X1 U2021 ( .A1(n4260), .A2(n370), .B1(n384), .B2(n661), .ZN(n2913) );
  OAI22_X1 U2022 ( .A1(n547), .A2(n3614), .B1(n3620), .B2(n858), .ZN(n2844) );
  OAI22_X1 U2023 ( .A1(n9), .A2(n562), .B1(n3619), .B2(n857), .ZN(n2845) );
  OAI22_X1 U2024 ( .A1(n547), .A2(n371), .B1(n380), .B2(n666), .ZN(n2908) );
  OAI22_X1 U2025 ( .A1(n212), .A2(n372), .B1(n375), .B2(n665), .ZN(n2909) );
  OAI22_X1 U2026 ( .A1(n546), .A2(n353), .B1(n361), .B2(n154), .ZN(n3164) );
  OAI22_X1 U2027 ( .A1(n235), .A2(n354), .B1(n357), .B2(n153), .ZN(n3165) );
  OAI22_X1 U2028 ( .A1(n400), .A2(n561), .B1(n3620), .B2(n861), .ZN(n2841) );
  OAI22_X1 U2029 ( .A1(n275), .A2(n3616), .B1(n3619), .B2(n860), .ZN(n2842) );
  OAI22_X1 U2030 ( .A1(n3614), .A2(n4266), .B1(n3618), .B2(n859), .ZN(n2843)
         );
  OAI22_X1 U2031 ( .A1(n239), .A2(n372), .B1(n380), .B2(n669), .ZN(n2905) );
  OAI22_X1 U2032 ( .A1(n7), .A2(n370), .B1(n382), .B2(n668), .ZN(n2906) );
  OAI22_X1 U2033 ( .A1(n1), .A2(n372), .B1(n375), .B2(n667), .ZN(n2907) );
  OAI22_X1 U2034 ( .A1(n4268), .A2(n354), .B1(n365), .B2(n157), .ZN(n3161) );
  OAI22_X1 U2035 ( .A1(n731), .A2(n288), .B1(n367), .B2(n156), .ZN(n3162) );
  OAI22_X1 U2036 ( .A1(n738), .A2(n354), .B1(n357), .B2(n155), .ZN(n3163) );
  OAI22_X1 U2037 ( .A1(n605), .A2(n3614), .B1(n3617), .B2(n833), .ZN(n2869) );
  OAI22_X1 U2038 ( .A1(n172), .A2(n372), .B1(n383), .B2(n641), .ZN(n2933) );
  OAI22_X1 U2039 ( .A1(n172), .A2(n1024), .B1(n1017), .B2(n513), .ZN(n2997) );
  OAI22_X1 U2040 ( .A1(n263), .A2(n354), .B1(n368), .B2(n129), .ZN(n3189) );
  OAI22_X1 U2041 ( .A1(n198), .A2(n3302), .B1(n1421), .B2(n352), .ZN(n3094) );
  OAI22_X1 U2042 ( .A1(n191), .A2(n3303), .B1(n1437), .B2(n351), .ZN(n3095) );
  OAI22_X1 U2043 ( .A1(n170), .A2(n3304), .B1(n1474), .B2(n350), .ZN(n3096) );
  OAI22_X1 U2044 ( .A1(n181), .A2(n3306), .B1(n3286), .B2(n340), .ZN(n3106) );
  OAI22_X1 U2045 ( .A1(n4258), .A2(n3308), .B1(n1538), .B2(n339), .ZN(n3107)
         );
  OAI22_X1 U2046 ( .A1(n269), .A2(n3309), .B1(n3289), .B2(n338), .ZN(n3108) );
  OAI22_X1 U2047 ( .A1(n401), .A2(n3310), .B1(n3288), .B2(n337), .ZN(n3109) );
  OAI22_X1 U2048 ( .A1(n3311), .A2(n553), .B1(n3287), .B2(n336), .ZN(n3110) );
  OAI22_X1 U2049 ( .A1(n739), .A2(n3312), .B1(n3286), .B2(n335), .ZN(n3111) );
  OAI22_X1 U2050 ( .A1(n602), .A2(n3302), .B1(n1538), .B2(n334), .ZN(n3112) );
  OAI22_X1 U2051 ( .A1(n26), .A2(n3309), .B1(n1474), .B2(n333), .ZN(n3113) );
  OAI22_X1 U2052 ( .A1(n702), .A2(n3313), .B1(n1437), .B2(n332), .ZN(n3114) );
  OAI22_X1 U2053 ( .A1(n708), .A2(n3314), .B1(n1421), .B2(n331), .ZN(n3115) );
  OAI22_X1 U2054 ( .A1(n10), .A2(n3307), .B1(n3535), .B2(n330), .ZN(n3116) );
  OAI22_X1 U2055 ( .A1(n698), .A2(n3316), .B1(n3299), .B2(n329), .ZN(n3117) );
  OAI22_X1 U2056 ( .A1(n280), .A2(n3302), .B1(n3298), .B2(n328), .ZN(n3118) );
  OAI22_X1 U2057 ( .A1(n4248), .A2(n3309), .B1(n3297), .B2(n327), .ZN(n3119)
         );
  OAI22_X1 U2058 ( .A1(n592), .A2(n3309), .B1(n3296), .B2(n326), .ZN(n3120) );
  OAI22_X1 U2059 ( .A1(n594), .A2(n3310), .B1(n3296), .B2(n325), .ZN(n3121) );
  OAI22_X1 U2060 ( .A1(net17879), .A2(n3311), .B1(n3295), .B2(n324), .ZN(n3122) );
  OAI22_X1 U2061 ( .A1(n742), .A2(n3312), .B1(n173), .B2(n323), .ZN(n3123) );
  OAI22_X1 U2062 ( .A1(n4244), .A2(n3315), .B1(n3534), .B2(n322), .ZN(n3124)
         );
  OAI22_X1 U2063 ( .A1(n607), .A2(n581), .B1(n583), .B2(n96), .ZN(n3222) );
  OAI22_X1 U2064 ( .A1(n673), .A2(n581), .B1(n583), .B2(n95), .ZN(n3223) );
  OAI22_X1 U2065 ( .A1(n225), .A2(n580), .B1(n585), .B2(n94), .ZN(n3224) );
  OAI22_X1 U2066 ( .A1(n274), .A2(n580), .B1(n588), .B2(n84), .ZN(n3234) );
  OAI22_X1 U2067 ( .A1(n599), .A2(n580), .B1(n585), .B2(n83), .ZN(n3235) );
  OAI22_X1 U2068 ( .A1(n4257), .A2(n580), .B1(n585), .B2(n82), .ZN(n3236) );
  OAI22_X1 U2069 ( .A1(n180), .A2(n580), .B1(n588), .B2(n81), .ZN(n3237) );
  OAI22_X1 U2070 ( .A1(n727), .A2(n580), .B1(n583), .B2(n80), .ZN(n3238) );
  OAI22_X1 U2071 ( .A1(n403), .A2(n580), .B1(n589), .B2(n79), .ZN(n3239) );
  OAI22_X1 U2072 ( .A1(n602), .A2(n580), .B1(n587), .B2(n78), .ZN(n3240) );
  OAI22_X1 U2073 ( .A1(n560), .A2(n581), .B1(n587), .B2(n77), .ZN(n3241) );
  OAI22_X1 U2074 ( .A1(n702), .A2(n580), .B1(n584), .B2(n76), .ZN(n3242) );
  OAI22_X1 U2075 ( .A1(n185), .A2(n581), .B1(n584), .B2(n75), .ZN(n3243) );
  OAI22_X1 U2076 ( .A1(n699), .A2(n580), .B1(n588), .B2(n74), .ZN(n3244) );
  OAI22_X1 U2077 ( .A1(n697), .A2(n581), .B1(n584), .B2(n73), .ZN(n3245) );
  OAI22_X1 U2078 ( .A1(n280), .A2(n580), .B1(n583), .B2(n72), .ZN(n3246) );
  OAI22_X1 U2079 ( .A1(n4248), .A2(n581), .B1(n589), .B2(n71), .ZN(n3247) );
  OAI22_X1 U2080 ( .A1(n591), .A2(n581), .B1(n588), .B2(n70), .ZN(n3248) );
  OAI22_X1 U2081 ( .A1(n593), .A2(n581), .B1(n587), .B2(n69), .ZN(n3249) );
  OAI22_X1 U2082 ( .A1(net44818), .A2(n581), .B1(n585), .B2(n68), .ZN(n3250)
         );
  OAI22_X1 U2083 ( .A1(n271), .A2(n581), .B1(n587), .B2(n67), .ZN(n3251) );
  OAI22_X1 U2084 ( .A1(n270), .A2(n580), .B1(n585), .B2(n66), .ZN(n3252) );
  OAI22_X1 U2085 ( .A1(n178), .A2(n3304), .B1(n3295), .B2(n342), .ZN(n3104) );
  OAI22_X1 U2086 ( .A1(n4260), .A2(n3306), .B1(n3287), .B2(n341), .ZN(n3105)
         );
  OAI22_X1 U2087 ( .A1(n674), .A2(n581), .B1(n588), .B2(n86), .ZN(n3232) );
  OAI22_X1 U2088 ( .A1(n575), .A2(n580), .B1(n584), .B2(n85), .ZN(n3233) );
  OAI22_X1 U2089 ( .A1(n547), .A2(n3315), .B1(n3292), .B2(n346), .ZN(n3100) );
  OAI22_X1 U2090 ( .A1(n705), .A2(n3308), .B1(n3293), .B2(n345), .ZN(n3101) );
  OAI22_X1 U2091 ( .A1(n547), .A2(n581), .B1(n584), .B2(n90), .ZN(n3228) );
  OAI22_X1 U2092 ( .A1(n235), .A2(n581), .B1(n583), .B2(n89), .ZN(n3229) );
  OAI22_X1 U2093 ( .A1(n238), .A2(n3305), .B1(n3288), .B2(n349), .ZN(n3097) );
  OAI22_X1 U2094 ( .A1(n731), .A2(n3302), .B1(n3289), .B2(n348), .ZN(n3098) );
  OAI22_X1 U2095 ( .A1(n738), .A2(n3306), .B1(n3290), .B2(n347), .ZN(n3099) );
  OAI22_X1 U2096 ( .A1(n605), .A2(n3306), .B1(n3294), .B2(n321), .ZN(n3125) );
  OAI22_X1 U2097 ( .A1(n732), .A2(n581), .B1(n589), .B2(n93), .ZN(n3225) );
  OAI22_X1 U2098 ( .A1(n7), .A2(n581), .B1(n587), .B2(n92), .ZN(n3226) );
  OAI22_X1 U2099 ( .A1(n554), .A2(n580), .B1(n589), .B2(n91), .ZN(n3227) );
  OAI22_X1 U2100 ( .A1(n4243), .A2(n581), .B1(n584), .B2(n65), .ZN(n3253) );
  OAI22_X1 U2101 ( .A1(n741), .A2(net26415), .B1(net26423), .B2(n436), .ZN(
        n3074) );
  OAI22_X1 U2102 ( .A1(n598), .A2(net26417), .B1(net26423), .B2(n435), .ZN(
        n3075) );
  OAI22_X1 U2103 ( .A1(n696), .A2(net26413), .B1(net26423), .B2(n434), .ZN(
        n3076) );
  OAI22_X1 U2104 ( .A1(n728), .A2(net44474), .B1(net26425), .B2(n433), .ZN(
        n3077) );
  OAI22_X1 U2105 ( .A1(net44473), .A2(n4256), .B1(net26425), .B2(n432), .ZN(
        n3078) );
  OAI22_X1 U2106 ( .A1(n4255), .A2(net26417), .B1(net26425), .B2(n431), .ZN(
        n3079) );
  OAI22_X1 U2107 ( .A1(n4254), .A2(net26415), .B1(net26425), .B2(n430), .ZN(
        n3080) );
  OAI22_X1 U2108 ( .A1(n260), .A2(net26417), .B1(net26425), .B2(n429), .ZN(
        n3081) );
  OAI22_X1 U2109 ( .A1(n208), .A2(net26413), .B1(net26427), .B2(n428), .ZN(
        n3082) );
  OAI22_X1 U2110 ( .A1(n185), .A2(net26417), .B1(net26427), .B2(n427), .ZN(
        n3083) );
  OAI22_X1 U2111 ( .A1(n182), .A2(net26417), .B1(net26427), .B2(n426), .ZN(
        n3084) );
  OAI22_X1 U2112 ( .A1(n224), .A2(net44473), .B1(net26427), .B2(n425), .ZN(
        n3085) );
  OAI22_X1 U2113 ( .A1(n4249), .A2(net44474), .B1(net26427), .B2(n424), .ZN(
        n3086) );
  OAI22_X1 U2114 ( .A1(net26415), .A2(n4248), .B1(net26429), .B2(n423), .ZN(
        n3087) );
  OAI22_X1 U2115 ( .A1(n4247), .A2(net26415), .B1(net26429), .B2(n422), .ZN(
        n3088) );
  OAI22_X1 U2116 ( .A1(net44473), .A2(n4246), .B1(net26429), .B2(n421), .ZN(
        n3089) );
  OAI22_X1 U2117 ( .A1(n197), .A2(net44474), .B1(net26429), .B2(n420), .ZN(
        n3090) );
  OAI22_X1 U2118 ( .A1(n743), .A2(net44473), .B1(net26429), .B2(n419), .ZN(
        n3091) );
  OAI22_X1 U2119 ( .A1(n270), .A2(net26415), .B1(net33812), .B2(n418), .ZN(
        n3092) );
  OAI22_X1 U2120 ( .A1(n607), .A2(n1143), .B1(n1049), .B2(n320), .ZN(n3126) );
  OAI22_X1 U2121 ( .A1(n4270), .A2(n1201), .B1(n1050), .B2(n319), .ZN(n3127)
         );
  OAI22_X1 U2122 ( .A1(n268), .A2(n1204), .B1(n1051), .B2(n318), .ZN(n3128) );
  OAI22_X1 U2123 ( .A1(n741), .A2(n1281), .B1(n1053), .B2(n308), .ZN(n3138) );
  OAI22_X1 U2124 ( .A1(n599), .A2(n1349), .B1(n1052), .B2(n307), .ZN(n3139) );
  OAI22_X1 U2125 ( .A1(n4257), .A2(n1269), .B1(n1055), .B2(n306), .ZN(n3140)
         );
  OAI22_X1 U2126 ( .A1(n281), .A2(n1271), .B1(n1054), .B2(n305), .ZN(n3141) );
  OAI22_X1 U2127 ( .A1(n553), .A2(n1281), .B1(n1062), .B2(n304), .ZN(n3142) );
  OAI22_X1 U2128 ( .A1(n739), .A2(n1349), .B1(n1053), .B2(n303), .ZN(n3143) );
  OAI22_X1 U2129 ( .A1(n415), .A2(n1204), .B1(n1052), .B2(n302), .ZN(n3144) );
  OAI22_X1 U2130 ( .A1(n4253), .A2(n1353), .B1(n1051), .B2(n301), .ZN(n3145)
         );
  OAI22_X1 U2131 ( .A1(n702), .A2(n1143), .B1(n1050), .B2(n300), .ZN(n3146) );
  OAI22_X1 U2132 ( .A1(n185), .A2(n1271), .B1(n1049), .B2(n299), .ZN(n3147) );
  OAI22_X1 U2133 ( .A1(n182), .A2(n1370), .B1(n1141), .B2(n298), .ZN(n3148) );
  OAI22_X1 U2134 ( .A1(n698), .A2(n1143), .B1(n1115), .B2(n297), .ZN(n3149) );
  OAI22_X1 U2135 ( .A1(n280), .A2(n1201), .B1(n1098), .B2(n296), .ZN(n3150) );
  OAI22_X1 U2136 ( .A1(n1400), .A2(n707), .B1(n1067), .B2(n295), .ZN(n3151) );
  OAI22_X1 U2137 ( .A1(n23), .A2(n1269), .B1(n1066), .B2(n294), .ZN(n3152) );
  OAI22_X1 U2138 ( .A1(n1271), .A2(n594), .B1(n1065), .B2(n293), .ZN(n3153) );
  OAI22_X1 U2139 ( .A1(net44818), .A2(n1281), .B1(n1063), .B2(n292), .ZN(n3154) );
  OAI22_X1 U2140 ( .A1(n743), .A2(n1349), .B1(n1062), .B2(n291), .ZN(n3155) );
  OAI22_X1 U2141 ( .A1(n4244), .A2(n1261), .B1(n1050), .B2(n290), .ZN(n3156)
         );
  OAI22_X1 U2142 ( .A1(n198), .A2(n566), .B1(n568), .B2(n64), .ZN(n3254) );
  OAI22_X1 U2143 ( .A1(n191), .A2(n566), .B1(n568), .B2(n63), .ZN(n3255) );
  OAI22_X1 U2144 ( .A1(n733), .A2(n565), .B1(n570), .B2(n62), .ZN(n3256) );
  OAI22_X1 U2145 ( .A1(n181), .A2(n566), .B1(n572), .B2(n52), .ZN(n3266) );
  OAI22_X1 U2146 ( .A1(n4258), .A2(n566), .B1(n570), .B2(n51), .ZN(n3267) );
  OAI22_X1 U2147 ( .A1(n269), .A2(n566), .B1(n570), .B2(n50), .ZN(n3268) );
  OAI22_X1 U2148 ( .A1(n188), .A2(n566), .B1(n572), .B2(n49), .ZN(n3269) );
  OAI22_X1 U2149 ( .A1(n727), .A2(n566), .B1(n568), .B2(n48), .ZN(n3270) );
  OAI22_X1 U2150 ( .A1(n739), .A2(n566), .B1(n573), .B2(n47), .ZN(n3271) );
  OAI22_X1 U2151 ( .A1(n415), .A2(n565), .B1(n571), .B2(n46), .ZN(n3272) );
  OAI22_X1 U2152 ( .A1(n4253), .A2(n566), .B1(n571), .B2(n45), .ZN(n3273) );
  OAI22_X1 U2153 ( .A1(n396), .A2(n565), .B1(n569), .B2(n44), .ZN(n3274) );
  OAI22_X1 U2154 ( .A1(n709), .A2(n566), .B1(n569), .B2(n43), .ZN(n3275) );
  OAI22_X1 U2155 ( .A1(n699), .A2(n565), .B1(n572), .B2(n42), .ZN(n3276) );
  OAI22_X1 U2156 ( .A1(n224), .A2(n566), .B1(n569), .B2(n41), .ZN(n3277) );
  OAI22_X1 U2157 ( .A1(n744), .A2(n565), .B1(n568), .B2(n40), .ZN(n3278) );
  OAI22_X1 U2158 ( .A1(n566), .A2(n706), .B1(n573), .B2(n39), .ZN(n3279) );
  OAI22_X1 U2159 ( .A1(n24), .A2(n565), .B1(n572), .B2(n38), .ZN(n3280) );
  OAI22_X1 U2160 ( .A1(n593), .A2(n565), .B1(n571), .B2(n37), .ZN(n3281) );
  OAI22_X1 U2161 ( .A1(net17879), .A2(n565), .B1(n570), .B2(n36), .ZN(n3282)
         );
  OAI22_X1 U2162 ( .A1(n743), .A2(n565), .B1(n571), .B2(n35), .ZN(n3283) );
  OAI22_X1 U2163 ( .A1(n221), .A2(n566), .B1(n570), .B2(n34), .ZN(n3284) );
  OAI22_X1 U2164 ( .A1(n4261), .A2(net26413), .B1(net26423), .B2(n438), .ZN(
        n3072) );
  OAI22_X1 U2165 ( .A1(n195), .A2(net26417), .B1(net26423), .B2(n437), .ZN(
        n3073) );
  OAI22_X1 U2166 ( .A1(n675), .A2(n1204), .B1(n1057), .B2(n310), .ZN(n3136) );
  OAI22_X1 U2167 ( .A1(n195), .A2(n1218), .B1(n1063), .B2(n309), .ZN(n3137) );
  OAI22_X1 U2168 ( .A1(n4261), .A2(n566), .B1(n572), .B2(n54), .ZN(n3264) );
  OAI22_X1 U2169 ( .A1(n574), .A2(n566), .B1(n569), .B2(n53), .ZN(n3265) );
  OAI22_X1 U2170 ( .A1(n4265), .A2(net26417), .B1(net26421), .B2(n442), .ZN(
        n3068) );
  OAI22_X1 U2171 ( .A1(n4264), .A2(net26413), .B1(net26421), .B2(n441), .ZN(
        n3069) );
  OAI22_X1 U2172 ( .A1(n546), .A2(n1281), .B1(n1059), .B2(n314), .ZN(n3132) );
  OAI22_X1 U2173 ( .A1(n212), .A2(n1349), .B1(n1060), .B2(n313), .ZN(n3133) );
  OAI22_X1 U2174 ( .A1(n547), .A2(n565), .B1(n569), .B2(n58), .ZN(n3260) );
  OAI22_X1 U2175 ( .A1(n235), .A2(n565), .B1(n568), .B2(n57), .ZN(n3261) );
  OAI22_X1 U2176 ( .A1(n172), .A2(net44474), .B1(net33812), .B2(n417), .ZN(
        n3093) );
  OAI22_X1 U2177 ( .A1(n4), .A2(n1218), .B1(n1054), .B2(n317), .ZN(n3129) );
  OAI22_X1 U2178 ( .A1(n193), .A2(n1261), .B1(n1055), .B2(n316), .ZN(n3130) );
  OAI22_X1 U2179 ( .A1(n1), .A2(n1261), .B1(n1050), .B2(n315), .ZN(n3131) );
  OAI22_X1 U2180 ( .A1(n263), .A2(n1269), .B1(n1061), .B2(n289), .ZN(n3157) );
  OAI22_X1 U2181 ( .A1(n4268), .A2(n565), .B1(n573), .B2(n61), .ZN(n3257) );
  OAI22_X1 U2182 ( .A1(n4267), .A2(n565), .B1(n571), .B2(n60), .ZN(n3258) );
  OAI22_X1 U2183 ( .A1(n738), .A2(n566), .B1(n573), .B2(n59), .ZN(n3259) );
  OAI22_X1 U2184 ( .A1(n4243), .A2(n565), .B1(n569), .B2(n33), .ZN(n3285) );
  OAI22_X1 U2185 ( .A1(n198), .A2(n3607), .B1(n3608), .B2(n832), .ZN(n2870) );
  OAI22_X1 U2186 ( .A1(n191), .A2(n3607), .B1(n3608), .B2(n831), .ZN(n2871) );
  OAI22_X1 U2187 ( .A1(n733), .A2(n3607), .B1(n3608), .B2(n830), .ZN(n2872) );
  OAI22_X1 U2188 ( .A1(n4271), .A2(n755), .B1(n754), .B2(n640), .ZN(n2934) );
  OAI22_X1 U2189 ( .A1(n673), .A2(n756), .B1(n205), .B2(n639), .ZN(n2935) );
  OAI22_X1 U2190 ( .A1(n268), .A2(n755), .B1(n3576), .B2(n638), .ZN(n2936) );
  OAI22_X1 U2191 ( .A1(n4271), .A2(n749), .B1(n3504), .B2(n128), .ZN(n3190) );
  OAI22_X1 U2192 ( .A1(n4270), .A2(n750), .B1(n8), .B2(n127), .ZN(n3191) );
  OAI22_X1 U2193 ( .A1(n194), .A2(n749), .B1(n748), .B2(n126), .ZN(n3192) );
  OAI22_X1 U2194 ( .A1(n4252), .A2(net38965), .B1(net38970), .B2(n940), .ZN(
        n2826) );
  OAI22_X1 U2195 ( .A1(n708), .A2(net38965), .B1(net38973), .B2(n939), .ZN(
        n2827) );
  OAI22_X1 U2196 ( .A1(n4251), .A2(net38966), .B1(net38968), .B2(n938), .ZN(
        n2828) );
  OAI22_X1 U2197 ( .A1(n4250), .A2(net38966), .B1(net38973), .B2(n937), .ZN(
        n2829) );
  OAI22_X1 U2198 ( .A1(n4249), .A2(net38966), .B1(net38974), .B2(n936), .ZN(
        n2830) );
  OAI22_X1 U2199 ( .A1(n28), .A2(net38964), .B1(net38973), .B2(n935), .ZN(
        n2831) );
  OAI22_X1 U2200 ( .A1(n21), .A2(n3606), .B1(n3610), .B2(n820), .ZN(n2882) );
  OAI22_X1 U2201 ( .A1(n177), .A2(n3606), .B1(n3610), .B2(n819), .ZN(n2883) );
  OAI22_X1 U2202 ( .A1(n696), .A2(n3606), .B1(n3610), .B2(n818), .ZN(n2884) );
  OAI22_X1 U2203 ( .A1(n729), .A2(n3606), .B1(n3611), .B2(n817), .ZN(n2885) );
  OAI22_X1 U2204 ( .A1(n4256), .A2(n3606), .B1(n3611), .B2(n816), .ZN(n2886)
         );
  OAI22_X1 U2205 ( .A1(n4255), .A2(n3606), .B1(n3611), .B2(n815), .ZN(n2887)
         );
  OAI22_X1 U2206 ( .A1(n4254), .A2(n3606), .B1(n3611), .B2(n814), .ZN(n2888)
         );
  OAI22_X1 U2207 ( .A1(n745), .A2(n3606), .B1(n3611), .B2(n813), .ZN(n2889) );
  OAI22_X1 U2208 ( .A1(n15), .A2(n756), .B1(n753), .B2(n628), .ZN(n2946) );
  OAI22_X1 U2209 ( .A1(n177), .A2(n757), .B1(n205), .B2(n627), .ZN(n2947) );
  OAI22_X1 U2210 ( .A1(n269), .A2(n755), .B1(n3578), .B2(n626), .ZN(n2948) );
  OAI22_X1 U2211 ( .A1(n401), .A2(n757), .B1(n3577), .B2(n625), .ZN(n2949) );
  OAI22_X1 U2212 ( .A1(n727), .A2(n756), .B1(n753), .B2(n624), .ZN(n2950) );
  OAI22_X1 U2213 ( .A1(n403), .A2(n757), .B1(n3578), .B2(n623), .ZN(n2951) );
  OAI22_X1 U2214 ( .A1(n602), .A2(n755), .B1(n205), .B2(n622), .ZN(n2952) );
  OAI22_X1 U2215 ( .A1(n26), .A2(n755), .B1(n3578), .B2(n621), .ZN(n2953) );
  OAI22_X1 U2216 ( .A1(n208), .A2(n757), .B1(n3576), .B2(n620), .ZN(n2954) );
  OAI22_X1 U2217 ( .A1(n183), .A2(n755), .B1(n3576), .B2(n618), .ZN(n2956) );
  OAI22_X1 U2218 ( .A1(n697), .A2(n757), .B1(n753), .B2(n617), .ZN(n2957) );
  OAI22_X1 U2219 ( .A1(n744), .A2(n756), .B1(n753), .B2(n616), .ZN(n2958) );
  OAI22_X1 U2220 ( .A1(n707), .A2(n757), .B1(n3578), .B2(n615), .ZN(n2959) );
  OAI22_X1 U2221 ( .A1(n591), .A2(n755), .B1(n3576), .B2(n614), .ZN(n2960) );
  OAI22_X1 U2222 ( .A1(n29), .A2(n755), .B1(n754), .B2(n613), .ZN(n2961) );
  OAI22_X1 U2223 ( .A1(n197), .A2(n756), .B1(n205), .B2(n612), .ZN(n2962) );
  OAI22_X1 U2224 ( .A1(n271), .A2(n756), .B1(n205), .B2(n611), .ZN(n2963) );
  OAI22_X1 U2225 ( .A1(n270), .A2(n755), .B1(n3576), .B2(n610), .ZN(n2964) );
  OAI22_X1 U2226 ( .A1(n4271), .A2(n926), .B1(n911), .B2(n512), .ZN(n2998) );
  OAI22_X1 U2227 ( .A1(n4270), .A2(n927), .B1(n911), .B2(n511), .ZN(n2999) );
  OAI22_X1 U2228 ( .A1(n4269), .A2(n928), .B1(n917), .B2(n510), .ZN(n3000) );
  OAI22_X1 U2229 ( .A1(n740), .A2(n928), .B1(n909), .B2(n500), .ZN(n3010) );
  OAI22_X1 U2230 ( .A1(n599), .A2(n993), .B1(n910), .B2(n499), .ZN(n3011) );
  OAI22_X1 U2231 ( .A1(n4257), .A2(n997), .B1(n912), .B2(n498), .ZN(n3012) );
  OAI22_X1 U2232 ( .A1(n281), .A2(n994), .B1(n913), .B2(n497), .ZN(n3013) );
  OAI22_X1 U2233 ( .A1(n995), .A2(n727), .B1(n916), .B2(n496), .ZN(n3014) );
  OAI22_X1 U2234 ( .A1(n403), .A2(n996), .B1(n914), .B2(n495), .ZN(n3015) );
  OAI22_X1 U2235 ( .A1(n602), .A2(n994), .B1(n915), .B2(n494), .ZN(n3016) );
  OAI22_X1 U2236 ( .A1(n560), .A2(n998), .B1(n918), .B2(n493), .ZN(n3017) );
  OAI22_X1 U2237 ( .A1(n6), .A2(n994), .B1(n909), .B2(n492), .ZN(n3018) );
  OAI22_X1 U2238 ( .A1(n709), .A2(n999), .B1(n908), .B2(n491), .ZN(n3019) );
  OAI22_X1 U2239 ( .A1(n10), .A2(n1000), .B1(n907), .B2(n490), .ZN(n3020) );
  OAI22_X1 U2240 ( .A1(n698), .A2(n1001), .B1(n906), .B2(n489), .ZN(n3021) );
  OAI22_X1 U2241 ( .A1(n744), .A2(n997), .B1(n920), .B2(n488), .ZN(n3022) );
  OAI22_X1 U2242 ( .A1(n184), .A2(n1002), .B1(n915), .B2(n487), .ZN(n3023) );
  OAI22_X1 U2243 ( .A1(n735), .A2(n994), .B1(n905), .B2(n486), .ZN(n3024) );
  OAI22_X1 U2244 ( .A1(n734), .A2(n997), .B1(n905), .B2(n485), .ZN(n3025) );
  OAI22_X1 U2245 ( .A1(net17879), .A2(n924), .B1(n920), .B2(n484), .ZN(n3026)
         );
  OAI22_X1 U2246 ( .A1(n743), .A2(n925), .B1(n919), .B2(n483), .ZN(n3027) );
  OAI22_X1 U2247 ( .A1(n4244), .A2(n926), .B1(n917), .B2(n482), .ZN(n3028) );
  OAI22_X1 U2248 ( .A1(n701), .A2(n751), .B1(n746), .B2(n108), .ZN(n3210) );
  OAI22_X1 U2249 ( .A1(n185), .A2(n749), .B1(n748), .B2(n107), .ZN(n3211) );
  OAI22_X1 U2250 ( .A1(n24), .A2(n751), .B1(n3503), .B2(n102), .ZN(n3216) );
  OAI22_X1 U2251 ( .A1(n734), .A2(n750), .B1(n8), .B2(n101), .ZN(n3217) );
  OAI22_X1 U2252 ( .A1(net39055), .A2(n751), .B1(n3503), .B2(n100), .ZN(n3218)
         );
  OAI22_X1 U2253 ( .A1(n5), .A2(n749), .B1(n3503), .B2(n99), .ZN(n3219) );
  OAI22_X1 U2254 ( .A1(n270), .A2(n749), .B1(n3503), .B2(n98), .ZN(n3220) );
  OAI22_X1 U2255 ( .A1(n674), .A2(n3606), .B1(n3610), .B2(n822), .ZN(n2880) );
  OAI22_X1 U2256 ( .A1(n574), .A2(n3606), .B1(n3610), .B2(n821), .ZN(n2881) );
  OAI22_X1 U2257 ( .A1(n675), .A2(n756), .B1(n3576), .B2(n630), .ZN(n2944) );
  OAI22_X1 U2258 ( .A1(n604), .A2(n756), .B1(n3576), .B2(n629), .ZN(n2945) );
  OAI22_X1 U2259 ( .A1(n675), .A2(n994), .B1(n912), .B2(n502), .ZN(n3008) );
  OAI22_X1 U2260 ( .A1(n575), .A2(n998), .B1(n908), .B2(n501), .ZN(n3009) );
  OAI22_X1 U2261 ( .A1(n4265), .A2(n3607), .B1(n3609), .B2(n826), .ZN(n2876)
         );
  OAI22_X1 U2262 ( .A1(n212), .A2(n3607), .B1(n3609), .B2(n825), .ZN(n2877) );
  OAI22_X1 U2263 ( .A1(n4265), .A2(n757), .B1(n3576), .B2(n634), .ZN(n2940) );
  OAI22_X1 U2264 ( .A1(n704), .A2(n755), .B1(n753), .B2(n633), .ZN(n2941) );
  OAI22_X1 U2265 ( .A1(n4265), .A2(n751), .B1(n3504), .B2(n122), .ZN(n3196) );
  OAI22_X1 U2266 ( .A1(n704), .A2(n749), .B1(n8), .B2(n121), .ZN(n3197) );
  OAI22_X1 U2267 ( .A1(n4265), .A2(n924), .B1(n910), .B2(n506), .ZN(n3004) );
  OAI22_X1 U2268 ( .A1(n9), .A2(n925), .B1(n918), .B2(n505), .ZN(n3005) );
  OAI22_X1 U2269 ( .A1(n22), .A2(n3607), .B1(n3608), .B2(n829), .ZN(n2873) );
  OAI22_X1 U2270 ( .A1(n731), .A2(n3607), .B1(n3608), .B2(n828), .ZN(n2874) );
  OAI22_X1 U2271 ( .A1(n4266), .A2(n3607), .B1(n3609), .B2(n827), .ZN(n2875)
         );
  OAI22_X1 U2272 ( .A1(n238), .A2(n756), .B1(n3577), .B2(n637), .ZN(n2937) );
  OAI22_X1 U2273 ( .A1(n193), .A2(n756), .B1(n3576), .B2(n636), .ZN(n2938) );
  OAI22_X1 U2274 ( .A1(n27), .A2(n757), .B1(n3578), .B2(n635), .ZN(n2939) );
  OAI22_X1 U2275 ( .A1(n239), .A2(n750), .B1(n3502), .B2(n125), .ZN(n3193) );
  OAI22_X1 U2276 ( .A1(n240), .A2(n750), .B1(n748), .B2(n124), .ZN(n3194) );
  OAI22_X1 U2277 ( .A1(n555), .A2(n751), .B1(n3502), .B2(n123), .ZN(n3195) );
  OAI22_X1 U2278 ( .A1(n605), .A2(n757), .B1(n3576), .B2(n609), .ZN(n2965) );
  OAI22_X1 U2279 ( .A1(n22), .A2(n993), .B1(n907), .B2(n509), .ZN(n3001) );
  OAI22_X1 U2280 ( .A1(n240), .A2(n1003), .B1(n906), .B2(n508), .ZN(n3002) );
  OAI22_X1 U2281 ( .A1(n554), .A2(n994), .B1(n920), .B2(n507), .ZN(n3003) );
  OAI22_X1 U2282 ( .A1(n4243), .A2(n927), .B1(n916), .B2(n481), .ZN(n3029) );
  OAI22_X1 U2283 ( .A1(n4243), .A2(n751), .B1(n746), .B2(n97), .ZN(n3221) );
  AND2_X1 U2284 ( .A1(ADD_RD2[0]), .A2(n2171), .ZN(n2169) );
  AND2_X1 U2285 ( .A1(ADD_RD1[0]), .A2(n2762), .ZN(n2760) );
  NAND4_X1 U2286 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(N343)
         );
  AOI221_X1 U2287 ( .B1(n3416), .B2(\registers[9][22] ), .C1(n3413), .C2(
        \registers[8][22] ), .A(n1792), .ZN(n1776) );
  AOI221_X1 U2288 ( .B1(n3428), .B2(\registers[13][22] ), .C1(n3425), .C2(
        \registers[12][22] ), .A(n1791), .ZN(n1777) );
  AOI211_X1 U2289 ( .C1(n3449), .C2(\registers[1][22] ), .A(n1788), .B(n1789), 
        .ZN(n1778) );
  NAND4_X1 U2290 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(N344)
         );
  AOI221_X1 U2291 ( .B1(n3416), .B2(\registers[9][23] ), .C1(n3413), .C2(
        \registers[8][23] ), .A(n1775), .ZN(n1759) );
  AOI221_X1 U2292 ( .B1(n3428), .B2(\registers[13][23] ), .C1(n3425), .C2(
        \registers[12][23] ), .A(n1774), .ZN(n1760) );
  AOI211_X1 U2293 ( .C1(n3449), .C2(\registers[1][23] ), .A(n1771), .B(n1772), 
        .ZN(n1761) );
  NAND4_X1 U2294 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(N345)
         );
  AOI221_X1 U2295 ( .B1(n3416), .B2(\registers[9][24] ), .C1(n3413), .C2(
        \registers[8][24] ), .A(n1758), .ZN(n1742) );
  AOI221_X1 U2296 ( .B1(n3428), .B2(\registers[13][24] ), .C1(n3425), .C2(
        \registers[12][24] ), .A(n1757), .ZN(n1743) );
  AOI211_X1 U2297 ( .C1(n3449), .C2(\registers[1][24] ), .A(n1754), .B(n1755), 
        .ZN(n1744) );
  NAND4_X1 U2298 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(N346)
         );
  AOI221_X1 U2299 ( .B1(n3416), .B2(\registers[9][25] ), .C1(n3413), .C2(
        \registers[8][25] ), .A(n1741), .ZN(n1725) );
  AOI221_X1 U2300 ( .B1(n3428), .B2(\registers[13][25] ), .C1(n3425), .C2(
        \registers[12][25] ), .A(n1740), .ZN(n1726) );
  AOI211_X1 U2301 ( .C1(n3449), .C2(\registers[1][25] ), .A(n1737), .B(n1738), 
        .ZN(n1727) );
  NAND4_X1 U2302 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(N347)
         );
  AOI221_X1 U2303 ( .B1(n3416), .B2(\registers[9][26] ), .C1(n3413), .C2(
        \registers[8][26] ), .A(n1724), .ZN(n1708) );
  AOI221_X1 U2304 ( .B1(n3428), .B2(\registers[13][26] ), .C1(n3425), .C2(
        \registers[12][26] ), .A(n1723), .ZN(n1709) );
  AOI211_X1 U2305 ( .C1(n3449), .C2(\registers[1][26] ), .A(n1720), .B(n1721), 
        .ZN(n1710) );
  NAND4_X1 U2306 ( .A1(n1691), .A2(n1692), .A3(n1693), .A4(n1694), .ZN(N348)
         );
  AOI221_X1 U2307 ( .B1(n3416), .B2(\registers[9][27] ), .C1(n3413), .C2(
        \registers[8][27] ), .A(n1707), .ZN(n1691) );
  AOI221_X1 U2308 ( .B1(n3428), .B2(\registers[13][27] ), .C1(n3425), .C2(
        \registers[12][27] ), .A(n1706), .ZN(n1692) );
  AOI211_X1 U2309 ( .C1(n3449), .C2(\registers[1][27] ), .A(n1703), .B(n1704), 
        .ZN(n1693) );
  NAND4_X1 U2310 ( .A1(n1674), .A2(n1675), .A3(n1676), .A4(n1677), .ZN(N349)
         );
  AOI221_X1 U2311 ( .B1(n3416), .B2(\registers[9][28] ), .C1(n3413), .C2(
        \registers[8][28] ), .A(n1690), .ZN(n1674) );
  AOI221_X1 U2312 ( .B1(n3428), .B2(\registers[13][28] ), .C1(n3425), .C2(
        \registers[12][28] ), .A(n1689), .ZN(n1675) );
  AOI211_X1 U2313 ( .C1(n3449), .C2(\registers[1][28] ), .A(n1686), .B(n1687), 
        .ZN(n1676) );
  NAND4_X1 U2314 ( .A1(n1657), .A2(n1658), .A3(n1659), .A4(n1660), .ZN(N350)
         );
  AOI221_X1 U2315 ( .B1(n3416), .B2(\registers[9][29] ), .C1(n3413), .C2(
        \registers[8][29] ), .A(n1673), .ZN(n1657) );
  AOI221_X1 U2316 ( .B1(n3428), .B2(\registers[13][29] ), .C1(n3425), .C2(
        \registers[12][29] ), .A(n1672), .ZN(n1658) );
  AOI211_X1 U2317 ( .C1(n3449), .C2(\registers[1][29] ), .A(n1669), .B(n1670), 
        .ZN(n1659) );
  NAND4_X1 U2318 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .ZN(N351)
         );
  AOI221_X1 U2319 ( .B1(n3416), .B2(\registers[9][30] ), .C1(n3413), .C2(
        \registers[8][30] ), .A(n1656), .ZN(n1640) );
  AOI221_X1 U2320 ( .B1(n3428), .B2(\registers[13][30] ), .C1(n3425), .C2(
        \registers[12][30] ), .A(n1655), .ZN(n1641) );
  AOI211_X1 U2321 ( .C1(n3449), .C2(\registers[1][30] ), .A(n1652), .B(n1653), 
        .ZN(n1642) );
  NAND4_X1 U2322 ( .A1(n1592), .A2(n1593), .A3(n1594), .A4(n1595), .ZN(N352)
         );
  AOI221_X1 U2323 ( .B1(n3416), .B2(\registers[9][31] ), .C1(n3413), .C2(
        \registers[8][31] ), .A(n1637), .ZN(n1592) );
  AOI221_X1 U2324 ( .B1(n3428), .B2(\registers[13][31] ), .C1(n3425), .C2(
        \registers[12][31] ), .A(n1632), .ZN(n1593) );
  AOI211_X1 U2325 ( .C1(n3449), .C2(\registers[1][31] ), .A(n1621), .B(n1622), 
        .ZN(n1594) );
  NAND4_X1 U2326 ( .A1(n2367), .A2(n2368), .A3(n2369), .A4(n2370), .ZN(N208)
         );
  AOI221_X1 U2327 ( .B1(n3329), .B2(\registers[9][22] ), .C1(n3326), .C2(
        \registers[8][22] ), .A(n2383), .ZN(n2367) );
  AOI221_X1 U2328 ( .B1(n3341), .B2(\registers[13][22] ), .C1(n3338), .C2(
        \registers[12][22] ), .A(n2382), .ZN(n2368) );
  AOI211_X1 U2329 ( .C1(n3362), .C2(\registers[1][22] ), .A(n2379), .B(n2380), 
        .ZN(n2369) );
  NAND4_X1 U2330 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(N209)
         );
  AOI221_X1 U2331 ( .B1(n3329), .B2(\registers[9][23] ), .C1(n3326), .C2(
        \registers[8][23] ), .A(n2366), .ZN(n2350) );
  AOI221_X1 U2332 ( .B1(n3341), .B2(\registers[13][23] ), .C1(n3338), .C2(
        \registers[12][23] ), .A(n2365), .ZN(n2351) );
  AOI211_X1 U2333 ( .C1(n3362), .C2(\registers[1][23] ), .A(n2362), .B(n2363), 
        .ZN(n2352) );
  NAND4_X1 U2334 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(N210)
         );
  AOI221_X1 U2335 ( .B1(n3329), .B2(\registers[9][24] ), .C1(n3326), .C2(
        \registers[8][24] ), .A(n2349), .ZN(n2333) );
  AOI221_X1 U2336 ( .B1(n3341), .B2(\registers[13][24] ), .C1(n3338), .C2(
        \registers[12][24] ), .A(n2348), .ZN(n2334) );
  AOI211_X1 U2337 ( .C1(n3362), .C2(\registers[1][24] ), .A(n2345), .B(n2346), 
        .ZN(n2335) );
  NAND4_X1 U2338 ( .A1(n2316), .A2(n2317), .A3(n2318), .A4(n2319), .ZN(N211)
         );
  AOI221_X1 U2339 ( .B1(n3329), .B2(\registers[9][25] ), .C1(n3326), .C2(
        \registers[8][25] ), .A(n2332), .ZN(n2316) );
  AOI221_X1 U2340 ( .B1(n3341), .B2(\registers[13][25] ), .C1(n3338), .C2(
        \registers[12][25] ), .A(n2331), .ZN(n2317) );
  AOI211_X1 U2341 ( .C1(n3362), .C2(\registers[1][25] ), .A(n2328), .B(n2329), 
        .ZN(n2318) );
  NAND4_X1 U2342 ( .A1(n2299), .A2(n2300), .A3(n2301), .A4(n2302), .ZN(N212)
         );
  AOI221_X1 U2343 ( .B1(n3329), .B2(\registers[9][26] ), .C1(n3326), .C2(
        \registers[8][26] ), .A(n2315), .ZN(n2299) );
  AOI221_X1 U2344 ( .B1(n3341), .B2(\registers[13][26] ), .C1(n3338), .C2(
        \registers[12][26] ), .A(n2314), .ZN(n2300) );
  AOI211_X1 U2345 ( .C1(n3362), .C2(\registers[1][26] ), .A(n2311), .B(n2312), 
        .ZN(n2301) );
  NAND4_X1 U2346 ( .A1(n2282), .A2(n2283), .A3(n2284), .A4(n2285), .ZN(N213)
         );
  AOI221_X1 U2347 ( .B1(n3329), .B2(\registers[9][27] ), .C1(n3326), .C2(
        \registers[8][27] ), .A(n2298), .ZN(n2282) );
  AOI221_X1 U2348 ( .B1(n3341), .B2(\registers[13][27] ), .C1(n3338), .C2(
        \registers[12][27] ), .A(n2297), .ZN(n2283) );
  AOI211_X1 U2349 ( .C1(n3362), .C2(\registers[1][27] ), .A(n2294), .B(n2295), 
        .ZN(n2284) );
  NAND4_X1 U2350 ( .A1(n2265), .A2(n2266), .A3(n2267), .A4(n2268), .ZN(N214)
         );
  AOI221_X1 U2351 ( .B1(n3329), .B2(\registers[9][28] ), .C1(n3326), .C2(
        \registers[8][28] ), .A(n2281), .ZN(n2265) );
  AOI221_X1 U2352 ( .B1(n3341), .B2(\registers[13][28] ), .C1(n3338), .C2(
        \registers[12][28] ), .A(n2280), .ZN(n2266) );
  AOI211_X1 U2353 ( .C1(n3362), .C2(\registers[1][28] ), .A(n2277), .B(n2278), 
        .ZN(n2267) );
  NAND4_X1 U2354 ( .A1(n2248), .A2(n2249), .A3(n2250), .A4(n2251), .ZN(N215)
         );
  AOI221_X1 U2355 ( .B1(n3329), .B2(\registers[9][29] ), .C1(n3326), .C2(
        \registers[8][29] ), .A(n2264), .ZN(n2248) );
  AOI221_X1 U2356 ( .B1(n3341), .B2(\registers[13][29] ), .C1(n3338), .C2(
        \registers[12][29] ), .A(n2263), .ZN(n2249) );
  AOI211_X1 U2357 ( .C1(n3362), .C2(\registers[1][29] ), .A(n2260), .B(n2261), 
        .ZN(n2250) );
  NAND4_X1 U2358 ( .A1(n2231), .A2(n2232), .A3(n2233), .A4(n2234), .ZN(N216)
         );
  AOI221_X1 U2359 ( .B1(n3329), .B2(\registers[9][30] ), .C1(n3326), .C2(
        \registers[8][30] ), .A(n2247), .ZN(n2231) );
  AOI221_X1 U2360 ( .B1(n3341), .B2(\registers[13][30] ), .C1(n3338), .C2(
        \registers[12][30] ), .A(n2246), .ZN(n2232) );
  AOI211_X1 U2361 ( .C1(n3362), .C2(\registers[1][30] ), .A(n2243), .B(n2244), 
        .ZN(n2233) );
  NAND4_X1 U2362 ( .A1(n2183), .A2(n2184), .A3(n2185), .A4(n2186), .ZN(N217)
         );
  AOI221_X1 U2363 ( .B1(n3329), .B2(\registers[9][31] ), .C1(n3326), .C2(
        \registers[8][31] ), .A(n2228), .ZN(n2183) );
  AOI221_X1 U2364 ( .B1(n3341), .B2(\registers[13][31] ), .C1(n3338), .C2(
        \registers[12][31] ), .A(n2223), .ZN(n2184) );
  AOI211_X1 U2365 ( .C1(n3362), .C2(\registers[1][31] ), .A(n2212), .B(n2213), 
        .ZN(n2185) );
  NAND4_X1 U2366 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .ZN(N321)
         );
  AOI221_X1 U2367 ( .B1(n3414), .B2(\registers[9][0] ), .C1(n3411), .C2(
        \registers[8][0] ), .A(n2181), .ZN(n2150) );
  AOI221_X1 U2368 ( .B1(n3426), .B2(\registers[13][0] ), .C1(n3423), .C2(
        \registers[12][0] ), .A(n2178), .ZN(n2151) );
  AOI211_X1 U2369 ( .C1(n3447), .C2(\registers[1][0] ), .A(n2172), .B(n2173), 
        .ZN(n2152) );
  NAND4_X1 U2370 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(N322)
         );
  AOI221_X1 U2371 ( .B1(n3414), .B2(\registers[9][1] ), .C1(n3411), .C2(
        \registers[8][1] ), .A(n2149), .ZN(n2133) );
  AOI221_X1 U2372 ( .B1(n3426), .B2(\registers[13][1] ), .C1(n3423), .C2(
        \registers[12][1] ), .A(n2148), .ZN(n2134) );
  AOI211_X1 U2373 ( .C1(n3447), .C2(\registers[1][1] ), .A(n2145), .B(n2146), 
        .ZN(n2135) );
  NAND4_X1 U2374 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(N323)
         );
  AOI221_X1 U2375 ( .B1(n3414), .B2(\registers[9][2] ), .C1(n3411), .C2(
        \registers[8][2] ), .A(n2132), .ZN(n2116) );
  AOI221_X1 U2376 ( .B1(n3426), .B2(\registers[13][2] ), .C1(n3423), .C2(
        \registers[12][2] ), .A(n2131), .ZN(n2117) );
  AOI211_X1 U2377 ( .C1(n3447), .C2(\registers[1][2] ), .A(n2128), .B(n2129), 
        .ZN(n2118) );
  NAND4_X1 U2378 ( .A1(n2099), .A2(n2100), .A3(n2101), .A4(n2102), .ZN(N324)
         );
  AOI221_X1 U2379 ( .B1(n3414), .B2(\registers[9][3] ), .C1(n3411), .C2(
        \registers[8][3] ), .A(n2115), .ZN(n2099) );
  AOI221_X1 U2380 ( .B1(n3426), .B2(\registers[13][3] ), .C1(n3423), .C2(
        \registers[12][3] ), .A(n2114), .ZN(n2100) );
  AOI211_X1 U2381 ( .C1(n3447), .C2(\registers[1][3] ), .A(n2111), .B(n2112), 
        .ZN(n2101) );
  NAND4_X1 U2382 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(N325)
         );
  AOI221_X1 U2383 ( .B1(n3414), .B2(\registers[9][4] ), .C1(n3411), .C2(
        \registers[8][4] ), .A(n2098), .ZN(n2082) );
  AOI221_X1 U2384 ( .B1(n3426), .B2(\registers[13][4] ), .C1(n3423), .C2(
        \registers[12][4] ), .A(n2097), .ZN(n2083) );
  AOI211_X1 U2385 ( .C1(n3447), .C2(\registers[1][4] ), .A(n2094), .B(n2095), 
        .ZN(n2084) );
  NAND4_X1 U2386 ( .A1(n2065), .A2(n2066), .A3(n2067), .A4(n2068), .ZN(N326)
         );
  AOI221_X1 U2387 ( .B1(n3414), .B2(\registers[9][5] ), .C1(n3411), .C2(
        \registers[8][5] ), .A(n2081), .ZN(n2065) );
  AOI221_X1 U2388 ( .B1(n3426), .B2(\registers[13][5] ), .C1(n3423), .C2(
        \registers[12][5] ), .A(n2080), .ZN(n2066) );
  AOI211_X1 U2389 ( .C1(n3447), .C2(\registers[1][5] ), .A(n2077), .B(n2078), 
        .ZN(n2067) );
  NAND4_X1 U2390 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(N327)
         );
  AOI221_X1 U2391 ( .B1(n3414), .B2(\registers[9][6] ), .C1(n3411), .C2(
        \registers[8][6] ), .A(n2064), .ZN(n2048) );
  AOI221_X1 U2392 ( .B1(n3426), .B2(\registers[13][6] ), .C1(n3423), .C2(
        \registers[12][6] ), .A(n2063), .ZN(n2049) );
  AOI211_X1 U2393 ( .C1(n3447), .C2(\registers[1][6] ), .A(n2060), .B(n2061), 
        .ZN(n2050) );
  NAND4_X1 U2394 ( .A1(n2031), .A2(n2032), .A3(n2033), .A4(n2034), .ZN(N328)
         );
  AOI221_X1 U2395 ( .B1(n3414), .B2(\registers[9][7] ), .C1(n3411), .C2(
        \registers[8][7] ), .A(n2047), .ZN(n2031) );
  AOI221_X1 U2396 ( .B1(n3426), .B2(\registers[13][7] ), .C1(n3423), .C2(
        \registers[12][7] ), .A(n2046), .ZN(n2032) );
  AOI211_X1 U2397 ( .C1(n3447), .C2(\registers[1][7] ), .A(n2043), .B(n2044), 
        .ZN(n2033) );
  NAND4_X1 U2398 ( .A1(n2014), .A2(n2015), .A3(n2016), .A4(n2017), .ZN(N329)
         );
  AOI221_X1 U2399 ( .B1(n3414), .B2(\registers[9][8] ), .C1(n3411), .C2(
        \registers[8][8] ), .A(n2030), .ZN(n2014) );
  AOI221_X1 U2400 ( .B1(n3426), .B2(\registers[13][8] ), .C1(n3423), .C2(
        \registers[12][8] ), .A(n2029), .ZN(n2015) );
  AOI211_X1 U2401 ( .C1(n3447), .C2(\registers[1][8] ), .A(n2026), .B(n2027), 
        .ZN(n2016) );
  NAND4_X1 U2402 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(N330)
         );
  AOI221_X1 U2403 ( .B1(n3414), .B2(\registers[9][9] ), .C1(n3411), .C2(
        \registers[8][9] ), .A(n2013), .ZN(n1997) );
  AOI221_X1 U2404 ( .B1(n3426), .B2(\registers[13][9] ), .C1(n3423), .C2(
        \registers[12][9] ), .A(n2012), .ZN(n1998) );
  AOI211_X1 U2405 ( .C1(n3447), .C2(\registers[1][9] ), .A(n2009), .B(n2010), 
        .ZN(n1999) );
  NAND4_X1 U2406 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .ZN(N331)
         );
  AOI221_X1 U2407 ( .B1(n3414), .B2(\registers[9][10] ), .C1(n3411), .C2(
        \registers[8][10] ), .A(n1996), .ZN(n1980) );
  AOI221_X1 U2408 ( .B1(n3426), .B2(\registers[13][10] ), .C1(n3423), .C2(
        \registers[12][10] ), .A(n1995), .ZN(n1981) );
  AOI211_X1 U2409 ( .C1(n3447), .C2(\registers[1][10] ), .A(n1992), .B(n1993), 
        .ZN(n1982) );
  NAND4_X1 U2410 ( .A1(n1963), .A2(n1964), .A3(n1965), .A4(n1966), .ZN(N332)
         );
  AOI221_X1 U2411 ( .B1(n3415), .B2(\registers[9][11] ), .C1(n3412), .C2(
        \registers[8][11] ), .A(n1979), .ZN(n1963) );
  AOI221_X1 U2412 ( .B1(n3427), .B2(\registers[13][11] ), .C1(n3424), .C2(
        \registers[12][11] ), .A(n1978), .ZN(n1964) );
  AOI211_X1 U2413 ( .C1(n3448), .C2(\registers[1][11] ), .A(n1975), .B(n1976), 
        .ZN(n1965) );
  NAND4_X1 U2414 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(N333)
         );
  AOI221_X1 U2415 ( .B1(n3415), .B2(\registers[9][12] ), .C1(n3412), .C2(
        \registers[8][12] ), .A(n1962), .ZN(n1946) );
  AOI221_X1 U2416 ( .B1(n3427), .B2(\registers[13][12] ), .C1(n3424), .C2(
        \registers[12][12] ), .A(n1961), .ZN(n1947) );
  AOI211_X1 U2417 ( .C1(n3448), .C2(\registers[1][12] ), .A(n1958), .B(n1959), 
        .ZN(n1948) );
  NAND4_X1 U2418 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(N334)
         );
  AOI221_X1 U2419 ( .B1(n3415), .B2(\registers[9][13] ), .C1(n3412), .C2(
        \registers[8][13] ), .A(n1945), .ZN(n1929) );
  AOI221_X1 U2420 ( .B1(n3427), .B2(\registers[13][13] ), .C1(n3424), .C2(
        \registers[12][13] ), .A(n1944), .ZN(n1930) );
  AOI211_X1 U2421 ( .C1(n3448), .C2(\registers[1][13] ), .A(n1941), .B(n1942), 
        .ZN(n1931) );
  NAND4_X1 U2422 ( .A1(n1912), .A2(n1913), .A3(n1914), .A4(n1915), .ZN(N335)
         );
  AOI221_X1 U2423 ( .B1(n3415), .B2(\registers[9][14] ), .C1(n3412), .C2(
        \registers[8][14] ), .A(n1928), .ZN(n1912) );
  AOI221_X1 U2424 ( .B1(n3427), .B2(\registers[13][14] ), .C1(n3424), .C2(
        \registers[12][14] ), .A(n1927), .ZN(n1913) );
  AOI211_X1 U2425 ( .C1(n3448), .C2(\registers[1][14] ), .A(n1924), .B(n1925), 
        .ZN(n1914) );
  NAND4_X1 U2426 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(N336)
         );
  AOI221_X1 U2427 ( .B1(n3415), .B2(\registers[9][15] ), .C1(n3412), .C2(
        \registers[8][15] ), .A(n1911), .ZN(n1895) );
  AOI221_X1 U2428 ( .B1(n3427), .B2(\registers[13][15] ), .C1(n3424), .C2(
        \registers[12][15] ), .A(n1910), .ZN(n1896) );
  AOI211_X1 U2429 ( .C1(n3448), .C2(\registers[1][15] ), .A(n1907), .B(n1908), 
        .ZN(n1897) );
  NAND4_X1 U2430 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .ZN(N337)
         );
  AOI221_X1 U2431 ( .B1(n3415), .B2(\registers[9][16] ), .C1(n3412), .C2(
        \registers[8][16] ), .A(n1894), .ZN(n1878) );
  AOI221_X1 U2432 ( .B1(n3427), .B2(\registers[13][16] ), .C1(n3424), .C2(
        \registers[12][16] ), .A(n1893), .ZN(n1879) );
  AOI211_X1 U2433 ( .C1(n3448), .C2(\registers[1][16] ), .A(n1890), .B(n1891), 
        .ZN(n1880) );
  NAND4_X1 U2434 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .ZN(N338)
         );
  AOI221_X1 U2435 ( .B1(n3415), .B2(\registers[9][17] ), .C1(n3412), .C2(
        \registers[8][17] ), .A(n1877), .ZN(n1861) );
  AOI221_X1 U2436 ( .B1(n3427), .B2(\registers[13][17] ), .C1(n3424), .C2(
        \registers[12][17] ), .A(n1876), .ZN(n1862) );
  AOI211_X1 U2437 ( .C1(n3448), .C2(\registers[1][17] ), .A(n1873), .B(n1874), 
        .ZN(n1863) );
  NAND4_X1 U2438 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .ZN(N339)
         );
  AOI221_X1 U2439 ( .B1(n3415), .B2(\registers[9][18] ), .C1(n3412), .C2(
        \registers[8][18] ), .A(n1860), .ZN(n1844) );
  AOI221_X1 U2440 ( .B1(n3427), .B2(\registers[13][18] ), .C1(n3424), .C2(
        \registers[12][18] ), .A(n1859), .ZN(n1845) );
  AOI211_X1 U2441 ( .C1(n3448), .C2(\registers[1][18] ), .A(n1856), .B(n1857), 
        .ZN(n1846) );
  NAND4_X1 U2442 ( .A1(n1827), .A2(n1828), .A3(n1829), .A4(n1830), .ZN(N340)
         );
  AOI221_X1 U2443 ( .B1(n3415), .B2(\registers[9][19] ), .C1(n3412), .C2(
        \registers[8][19] ), .A(n1843), .ZN(n1827) );
  AOI221_X1 U2444 ( .B1(n3427), .B2(\registers[13][19] ), .C1(n3424), .C2(
        \registers[12][19] ), .A(n1842), .ZN(n1828) );
  AOI211_X1 U2445 ( .C1(n3448), .C2(\registers[1][19] ), .A(n1839), .B(n1840), 
        .ZN(n1829) );
  NAND4_X1 U2446 ( .A1(n1810), .A2(n1811), .A3(n1812), .A4(n1813), .ZN(N341)
         );
  AOI221_X1 U2447 ( .B1(n3415), .B2(\registers[9][20] ), .C1(n3412), .C2(
        \registers[8][20] ), .A(n1826), .ZN(n1810) );
  AOI221_X1 U2448 ( .B1(n3427), .B2(\registers[13][20] ), .C1(n3424), .C2(
        \registers[12][20] ), .A(n1825), .ZN(n1811) );
  AOI211_X1 U2449 ( .C1(n3448), .C2(\registers[1][20] ), .A(n1822), .B(n1823), 
        .ZN(n1812) );
  NAND4_X1 U2450 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .ZN(N342)
         );
  AOI221_X1 U2451 ( .B1(n3415), .B2(\registers[9][21] ), .C1(n3412), .C2(
        \registers[8][21] ), .A(n1809), .ZN(n1793) );
  AOI221_X1 U2452 ( .B1(n3427), .B2(\registers[13][21] ), .C1(n3424), .C2(
        \registers[12][21] ), .A(n1808), .ZN(n1794) );
  AOI211_X1 U2453 ( .C1(n3448), .C2(\registers[1][21] ), .A(n1805), .B(n1806), 
        .ZN(n1795) );
  NAND4_X1 U2454 ( .A1(n2741), .A2(n2742), .A3(n2743), .A4(n2744), .ZN(N186)
         );
  AOI221_X1 U2455 ( .B1(n3327), .B2(\registers[9][0] ), .C1(n3324), .C2(
        \registers[8][0] ), .A(n2772), .ZN(n2741) );
  AOI221_X1 U2456 ( .B1(n3339), .B2(\registers[13][0] ), .C1(n3336), .C2(
        \registers[12][0] ), .A(n2769), .ZN(n2742) );
  AOI211_X1 U2457 ( .C1(n3360), .C2(\registers[1][0] ), .A(n2763), .B(n2764), 
        .ZN(n2743) );
  NAND4_X1 U2458 ( .A1(n2724), .A2(n2725), .A3(n2726), .A4(n2727), .ZN(N187)
         );
  AOI221_X1 U2459 ( .B1(n3327), .B2(\registers[9][1] ), .C1(n3324), .C2(
        \registers[8][1] ), .A(n2740), .ZN(n2724) );
  AOI221_X1 U2460 ( .B1(n3339), .B2(\registers[13][1] ), .C1(n3336), .C2(
        \registers[12][1] ), .A(n2739), .ZN(n2725) );
  AOI211_X1 U2461 ( .C1(n3360), .C2(\registers[1][1] ), .A(n2736), .B(n2737), 
        .ZN(n2726) );
  NAND4_X1 U2462 ( .A1(n2707), .A2(n2708), .A3(n2709), .A4(n2710), .ZN(N188)
         );
  AOI221_X1 U2463 ( .B1(n3327), .B2(\registers[9][2] ), .C1(n3324), .C2(
        \registers[8][2] ), .A(n2723), .ZN(n2707) );
  AOI221_X1 U2464 ( .B1(n3339), .B2(\registers[13][2] ), .C1(n3336), .C2(
        \registers[12][2] ), .A(n2722), .ZN(n2708) );
  AOI211_X1 U2465 ( .C1(n3360), .C2(\registers[1][2] ), .A(n2719), .B(n2720), 
        .ZN(n2709) );
  NAND4_X1 U2466 ( .A1(n2690), .A2(n2691), .A3(n2692), .A4(n2693), .ZN(N189)
         );
  AOI221_X1 U2467 ( .B1(n3327), .B2(\registers[9][3] ), .C1(n3324), .C2(
        \registers[8][3] ), .A(n2706), .ZN(n2690) );
  AOI221_X1 U2468 ( .B1(n3339), .B2(\registers[13][3] ), .C1(n3336), .C2(
        \registers[12][3] ), .A(n2705), .ZN(n2691) );
  AOI211_X1 U2469 ( .C1(n3360), .C2(\registers[1][3] ), .A(n2702), .B(n2703), 
        .ZN(n2692) );
  NAND4_X1 U2470 ( .A1(n2673), .A2(n2674), .A3(n2675), .A4(n2676), .ZN(N190)
         );
  AOI221_X1 U2471 ( .B1(n3327), .B2(\registers[9][4] ), .C1(n3324), .C2(
        \registers[8][4] ), .A(n2689), .ZN(n2673) );
  AOI221_X1 U2472 ( .B1(n3339), .B2(\registers[13][4] ), .C1(n3336), .C2(
        \registers[12][4] ), .A(n2688), .ZN(n2674) );
  AOI211_X1 U2473 ( .C1(n3360), .C2(\registers[1][4] ), .A(n2685), .B(n2686), 
        .ZN(n2675) );
  NAND4_X1 U2474 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(N191)
         );
  AOI221_X1 U2475 ( .B1(n3327), .B2(\registers[9][5] ), .C1(n3324), .C2(
        \registers[8][5] ), .A(n2672), .ZN(n2656) );
  AOI221_X1 U2476 ( .B1(n3339), .B2(\registers[13][5] ), .C1(n3336), .C2(
        \registers[12][5] ), .A(n2671), .ZN(n2657) );
  AOI211_X1 U2477 ( .C1(n3360), .C2(\registers[1][5] ), .A(n2668), .B(n2669), 
        .ZN(n2658) );
  NAND4_X1 U2478 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2642), .ZN(N192)
         );
  AOI221_X1 U2479 ( .B1(n3327), .B2(\registers[9][6] ), .C1(n3324), .C2(
        \registers[8][6] ), .A(n2655), .ZN(n2639) );
  AOI221_X1 U2480 ( .B1(n3339), .B2(\registers[13][6] ), .C1(n3336), .C2(
        \registers[12][6] ), .A(n2654), .ZN(n2640) );
  AOI211_X1 U2481 ( .C1(n3360), .C2(\registers[1][6] ), .A(n2651), .B(n2652), 
        .ZN(n2641) );
  NAND4_X1 U2482 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(N193)
         );
  AOI221_X1 U2483 ( .B1(n3327), .B2(\registers[9][7] ), .C1(n3324), .C2(
        \registers[8][7] ), .A(n2638), .ZN(n2622) );
  AOI221_X1 U2484 ( .B1(n3339), .B2(\registers[13][7] ), .C1(n3336), .C2(
        \registers[12][7] ), .A(n2637), .ZN(n2623) );
  AOI211_X1 U2485 ( .C1(n3360), .C2(\registers[1][7] ), .A(n2634), .B(n2635), 
        .ZN(n2624) );
  NAND4_X1 U2486 ( .A1(n2605), .A2(n2606), .A3(n2607), .A4(n2608), .ZN(N194)
         );
  AOI221_X1 U2487 ( .B1(n3327), .B2(\registers[9][8] ), .C1(n3324), .C2(
        \registers[8][8] ), .A(n2621), .ZN(n2605) );
  AOI221_X1 U2488 ( .B1(n3339), .B2(\registers[13][8] ), .C1(n3336), .C2(
        \registers[12][8] ), .A(n2620), .ZN(n2606) );
  AOI211_X1 U2489 ( .C1(n3360), .C2(\registers[1][8] ), .A(n2617), .B(n2618), 
        .ZN(n2607) );
  NAND4_X1 U2490 ( .A1(n2588), .A2(n2589), .A3(n2590), .A4(n2591), .ZN(N195)
         );
  AOI221_X1 U2491 ( .B1(n3327), .B2(\registers[9][9] ), .C1(n3324), .C2(
        \registers[8][9] ), .A(n2604), .ZN(n2588) );
  AOI221_X1 U2492 ( .B1(n3339), .B2(\registers[13][9] ), .C1(n3336), .C2(
        \registers[12][9] ), .A(n2603), .ZN(n2589) );
  AOI211_X1 U2493 ( .C1(n3360), .C2(\registers[1][9] ), .A(n2600), .B(n2601), 
        .ZN(n2590) );
  NAND4_X1 U2494 ( .A1(n2571), .A2(n2572), .A3(n2573), .A4(n2574), .ZN(N196)
         );
  AOI221_X1 U2495 ( .B1(n3327), .B2(\registers[9][10] ), .C1(n3324), .C2(
        \registers[8][10] ), .A(n2587), .ZN(n2571) );
  AOI221_X1 U2496 ( .B1(n3339), .B2(\registers[13][10] ), .C1(n3336), .C2(
        \registers[12][10] ), .A(n2586), .ZN(n2572) );
  AOI211_X1 U2497 ( .C1(n3360), .C2(\registers[1][10] ), .A(n2583), .B(n2584), 
        .ZN(n2573) );
  NAND4_X1 U2498 ( .A1(n2554), .A2(n2555), .A3(n2556), .A4(n2557), .ZN(N197)
         );
  AOI221_X1 U2499 ( .B1(n3328), .B2(\registers[9][11] ), .C1(n3325), .C2(
        \registers[8][11] ), .A(n2570), .ZN(n2554) );
  AOI221_X1 U2500 ( .B1(n3340), .B2(\registers[13][11] ), .C1(n3337), .C2(
        \registers[12][11] ), .A(n2569), .ZN(n2555) );
  AOI211_X1 U2501 ( .C1(n3361), .C2(\registers[1][11] ), .A(n2566), .B(n2567), 
        .ZN(n2556) );
  NAND4_X1 U2502 ( .A1(n2537), .A2(n2538), .A3(n2539), .A4(n2540), .ZN(N198)
         );
  AOI221_X1 U2503 ( .B1(n3328), .B2(\registers[9][12] ), .C1(n3325), .C2(
        \registers[8][12] ), .A(n2553), .ZN(n2537) );
  AOI221_X1 U2504 ( .B1(n3340), .B2(\registers[13][12] ), .C1(n3337), .C2(
        \registers[12][12] ), .A(n2552), .ZN(n2538) );
  AOI211_X1 U2505 ( .C1(n3361), .C2(\registers[1][12] ), .A(n2549), .B(n2550), 
        .ZN(n2539) );
  NAND4_X1 U2506 ( .A1(n2520), .A2(n2521), .A3(n2522), .A4(n2523), .ZN(N199)
         );
  AOI221_X1 U2507 ( .B1(n3328), .B2(\registers[9][13] ), .C1(n3325), .C2(
        \registers[8][13] ), .A(n2536), .ZN(n2520) );
  AOI221_X1 U2508 ( .B1(n3340), .B2(\registers[13][13] ), .C1(n3337), .C2(
        \registers[12][13] ), .A(n2535), .ZN(n2521) );
  AOI211_X1 U2509 ( .C1(n3361), .C2(\registers[1][13] ), .A(n2532), .B(n2533), 
        .ZN(n2522) );
  NAND4_X1 U2510 ( .A1(n2503), .A2(n2504), .A3(n2505), .A4(n2506), .ZN(N200)
         );
  AOI221_X1 U2511 ( .B1(n3328), .B2(\registers[9][14] ), .C1(n3325), .C2(
        \registers[8][14] ), .A(n2519), .ZN(n2503) );
  AOI221_X1 U2512 ( .B1(n3340), .B2(\registers[13][14] ), .C1(n3337), .C2(
        \registers[12][14] ), .A(n2518), .ZN(n2504) );
  AOI211_X1 U2513 ( .C1(n3361), .C2(\registers[1][14] ), .A(n2515), .B(n2516), 
        .ZN(n2505) );
  NAND4_X1 U2514 ( .A1(n2486), .A2(n2487), .A3(n2488), .A4(n2489), .ZN(N201)
         );
  AOI221_X1 U2515 ( .B1(n3328), .B2(\registers[9][15] ), .C1(n3325), .C2(
        \registers[8][15] ), .A(n2502), .ZN(n2486) );
  AOI221_X1 U2516 ( .B1(n3340), .B2(\registers[13][15] ), .C1(n3337), .C2(
        \registers[12][15] ), .A(n2501), .ZN(n2487) );
  AOI211_X1 U2517 ( .C1(n3361), .C2(\registers[1][15] ), .A(n2498), .B(n2499), 
        .ZN(n2488) );
  NAND4_X1 U2518 ( .A1(n2469), .A2(n2470), .A3(n2471), .A4(n2472), .ZN(N202)
         );
  AOI221_X1 U2519 ( .B1(n3328), .B2(\registers[9][16] ), .C1(n3325), .C2(
        \registers[8][16] ), .A(n2485), .ZN(n2469) );
  AOI221_X1 U2520 ( .B1(n3340), .B2(\registers[13][16] ), .C1(n3337), .C2(
        \registers[12][16] ), .A(n2484), .ZN(n2470) );
  AOI211_X1 U2521 ( .C1(n3361), .C2(\registers[1][16] ), .A(n2481), .B(n2482), 
        .ZN(n2471) );
  NAND4_X1 U2522 ( .A1(n2452), .A2(n2453), .A3(n2454), .A4(n2455), .ZN(N203)
         );
  AOI221_X1 U2523 ( .B1(n3328), .B2(\registers[9][17] ), .C1(n3325), .C2(
        \registers[8][17] ), .A(n2468), .ZN(n2452) );
  AOI221_X1 U2524 ( .B1(n3340), .B2(\registers[13][17] ), .C1(n3337), .C2(
        \registers[12][17] ), .A(n2467), .ZN(n2453) );
  AOI211_X1 U2525 ( .C1(n3361), .C2(\registers[1][17] ), .A(n2464), .B(n2465), 
        .ZN(n2454) );
  NAND4_X1 U2526 ( .A1(n2435), .A2(n2436), .A3(n2437), .A4(n2438), .ZN(N204)
         );
  AOI221_X1 U2527 ( .B1(n3328), .B2(\registers[9][18] ), .C1(n3325), .C2(
        \registers[8][18] ), .A(n2451), .ZN(n2435) );
  AOI221_X1 U2528 ( .B1(n3340), .B2(\registers[13][18] ), .C1(n3337), .C2(
        \registers[12][18] ), .A(n2450), .ZN(n2436) );
  AOI211_X1 U2529 ( .C1(n3361), .C2(\registers[1][18] ), .A(n2447), .B(n2448), 
        .ZN(n2437) );
  NAND4_X1 U2530 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(N205)
         );
  AOI221_X1 U2531 ( .B1(n3328), .B2(\registers[9][19] ), .C1(n3325), .C2(
        \registers[8][19] ), .A(n2434), .ZN(n2418) );
  AOI221_X1 U2532 ( .B1(n3340), .B2(\registers[13][19] ), .C1(n3337), .C2(
        \registers[12][19] ), .A(n2433), .ZN(n2419) );
  AOI211_X1 U2533 ( .C1(n3361), .C2(\registers[1][19] ), .A(n2430), .B(n2431), 
        .ZN(n2420) );
  NAND4_X1 U2534 ( .A1(n2401), .A2(n2402), .A3(n2403), .A4(n2404), .ZN(N206)
         );
  AOI221_X1 U2535 ( .B1(n3328), .B2(\registers[9][20] ), .C1(n3325), .C2(
        \registers[8][20] ), .A(n2417), .ZN(n2401) );
  AOI221_X1 U2536 ( .B1(n3340), .B2(\registers[13][20] ), .C1(n3337), .C2(
        \registers[12][20] ), .A(n2416), .ZN(n2402) );
  AOI211_X1 U2537 ( .C1(n3361), .C2(\registers[1][20] ), .A(n2413), .B(n2414), 
        .ZN(n2403) );
  NAND4_X1 U2538 ( .A1(n2384), .A2(n2385), .A3(n2386), .A4(n2387), .ZN(N207)
         );
  AOI221_X1 U2539 ( .B1(n3328), .B2(\registers[9][21] ), .C1(n3325), .C2(
        \registers[8][21] ), .A(n2400), .ZN(n2384) );
  AOI221_X1 U2540 ( .B1(n3340), .B2(\registers[13][21] ), .C1(n3337), .C2(
        \registers[12][21] ), .A(n2399), .ZN(n2385) );
  AOI211_X1 U2541 ( .C1(n3361), .C2(\registers[1][21] ), .A(n2396), .B(n2397), 
        .ZN(n2386) );
  NOR2_X1 U2542 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n2177) );
  NOR2_X1 U2543 ( .A1(n4240), .A2(ADD_RD2[4]), .ZN(n2182) );
  NOR2_X1 U2544 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n2768) );
  NOR2_X1 U2545 ( .A1(n4237), .A2(ADD_RD1[4]), .ZN(n2773) );
  AND2_X1 U2546 ( .A1(n2166), .A2(ADD_RD2[0]), .ZN(n2161) );
  AND2_X1 U2547 ( .A1(n2177), .A2(ADD_RD2[0]), .ZN(n2174) );
  AND2_X1 U2548 ( .A1(n2182), .A2(ADD_RD2[0]), .ZN(n2179) );
  AND2_X1 U2549 ( .A1(n2757), .A2(ADD_RD1[0]), .ZN(n2752) );
  AND2_X1 U2550 ( .A1(n2768), .A2(ADD_RD1[0]), .ZN(n2765) );
  AND2_X1 U2551 ( .A1(n2773), .A2(ADD_RD1[0]), .ZN(n2770) );
  INV_X1 U2552 ( .A(ADD_RD2[0]), .ZN(n4242) );
  INV_X1 U2553 ( .A(ADD_RD1[0]), .ZN(n4239) );
  INV_X1 U2554 ( .A(ADD_RD2[1]), .ZN(n4241) );
  INV_X1 U2555 ( .A(ADD_RD2[3]), .ZN(n4240) );
  INV_X1 U2556 ( .A(ADD_RD1[1]), .ZN(n4238) );
  INV_X1 U2557 ( .A(ADD_RD1[3]), .ZN(n4237) );
  AND2_X1 U2558 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n2171) );
  AND2_X1 U2559 ( .A1(ADD_RD2[4]), .A2(n4240), .ZN(n2166) );
  AND2_X1 U2560 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2762) );
  AND2_X1 U2561 ( .A1(ADD_RD1[4]), .A2(n4237), .ZN(n2757) );
  INV_X1 U2562 ( .A(n1325), .ZN(n3994) );
  AOI22_X1 U2563 ( .A1(n30), .A2(n3562), .B1(n3565), .B2(\registers[18][8] ), 
        .ZN(n1325) );
  INV_X1 U2564 ( .A(n1326), .ZN(n3995) );
  AOI22_X1 U2565 ( .A1(n780), .A2(n3563), .B1(n3565), .B2(\registers[18][9] ), 
        .ZN(n1326) );
  INV_X1 U2566 ( .A(n1292), .ZN(n4026) );
  AOI22_X1 U2567 ( .A1(n30), .A2(n760), .B1(n3572), .B2(\registers[19][8] ), 
        .ZN(n1292) );
  INV_X1 U2568 ( .A(n1293), .ZN(n4027) );
  AOI22_X1 U2569 ( .A1(n282), .A2(n761), .B1(n3572), .B2(\registers[19][9] ), 
        .ZN(n1293) );
  INV_X1 U2570 ( .A(n1154), .ZN(n4147) );
  AOI22_X1 U2571 ( .A1(n782), .A2(n3595), .B1(n3603), .B2(\registers[25][8] ), 
        .ZN(n1154) );
  INV_X1 U2572 ( .A(n1155), .ZN(n4148) );
  AOI22_X1 U2573 ( .A1(n780), .A2(n737), .B1(n3600), .B2(\registers[25][9] ), 
        .ZN(n1155) );
  INV_X1 U2574 ( .A(n1363), .ZN(n3867) );
  AOI22_X1 U2575 ( .A1(n782), .A2(n3545), .B1(n220), .B2(\registers[13][8] ), 
        .ZN(n1363) );
  INV_X1 U2576 ( .A(n1364), .ZN(n3868) );
  AOI22_X1 U2577 ( .A1(n282), .A2(n776), .B1(n17), .B2(\registers[13][9] ), 
        .ZN(n1364) );
  INV_X1 U2578 ( .A(n1396), .ZN(n3836) );
  AOI22_X1 U2579 ( .A1(n782), .A2(n203), .B1(n3542), .B2(\registers[12][8] ), 
        .ZN(n1396) );
  INV_X1 U2580 ( .A(n1397), .ZN(n3837) );
  AOI22_X1 U2581 ( .A1(n282), .A2(n770), .B1(n3540), .B2(\registers[12][9] ), 
        .ZN(n1397) );
  INV_X1 U2582 ( .A(n1082), .ZN(n4210) );
  AOI22_X1 U2583 ( .A1(n30), .A2(n3633), .B1(n3636), .B2(\registers[29][8] ), 
        .ZN(n1082) );
  INV_X1 U2584 ( .A(n1083), .ZN(n4211) );
  AOI22_X1 U2585 ( .A1(n780), .A2(n3634), .B1(n3637), .B2(\registers[29][9] ), 
        .ZN(n1083) );
  INV_X1 U2586 ( .A(n1116), .ZN(n4178) );
  AOI22_X1 U2587 ( .A1(n782), .A2(n767), .B1(n3626), .B2(\registers[28][8] ), 
        .ZN(n1116) );
  INV_X1 U2588 ( .A(n1117), .ZN(n4179) );
  AOI22_X1 U2589 ( .A1(n780), .A2(n688), .B1(n3626), .B2(\registers[28][9] ), 
        .ZN(n1117) );
  INV_X1 U2590 ( .A(n1223), .ZN(n4085) );
  AOI22_X1 U2591 ( .A1(n782), .A2(n3582), .B1(n3586), .B2(\registers[23][8] ), 
        .ZN(n1223) );
  INV_X1 U2592 ( .A(n1224), .ZN(n4086) );
  AOI22_X1 U2593 ( .A1(n282), .A2(n3582), .B1(n3585), .B2(\registers[23][9] ), 
        .ZN(n1224) );
  INV_X1 U2594 ( .A(n1497), .ZN(n3961) );
  AOI22_X1 U2595 ( .A1(n30), .A2(n682), .B1(n3507), .B2(\registers[7][8] ), 
        .ZN(n1497) );
  INV_X1 U2596 ( .A(n1498), .ZN(n3962) );
  AOI22_X1 U2597 ( .A1(n780), .A2(n764), .B1(n3508), .B2(\registers[7][9] ), 
        .ZN(n1498) );
  INV_X1 U2598 ( .A(n1431), .ZN(n3805) );
  AOI22_X1 U2599 ( .A1(n782), .A2(n3520), .B1(n3526), .B2(\registers[9][8] ), 
        .ZN(n1431) );
  INV_X1 U2600 ( .A(n1432), .ZN(n3806) );
  AOI22_X1 U2601 ( .A1(n282), .A2(n3519), .B1(n3526), .B2(\registers[9][9] ), 
        .ZN(n1432) );
  INV_X1 U2602 ( .A(n1568), .ZN(n3898) );
  AOI22_X1 U2603 ( .A1(n30), .A2(n3493), .B1(n3500), .B2(\registers[1][8] ), 
        .ZN(n1568) );
  INV_X1 U2604 ( .A(n1569), .ZN(n3899) );
  AOI22_X1 U2605 ( .A1(n780), .A2(n3493), .B1(n3500), .B2(\registers[1][9] ), 
        .ZN(n1569) );
  INV_X1 U2606 ( .A(n1257), .ZN(n4058) );
  AOI22_X1 U2607 ( .A1(n782), .A2(net26243), .B1(net26249), .B2(
        \registers[22][8] ), .ZN(n1257) );
  INV_X1 U2608 ( .A(n1258), .ZN(n4059) );
  AOI22_X1 U2609 ( .A1(n282), .A2(net26247), .B1(n20), .B2(\registers[22][9] ), 
        .ZN(n1258) );
  INV_X1 U2610 ( .A(n1531), .ZN(n3930) );
  AOI22_X1 U2611 ( .A1(n782), .A2(n229), .B1(net26585), .B2(\registers[6][8] ), 
        .ZN(n1531) );
  INV_X1 U2612 ( .A(n1532), .ZN(n3931) );
  AOI22_X1 U2613 ( .A1(n780), .A2(n228), .B1(net26589), .B2(\registers[6][9] ), 
        .ZN(n1532) );
  INV_X1 U2614 ( .A(n1464), .ZN(n3774) );
  AOI22_X1 U2615 ( .A1(n30), .A2(n3512), .B1(n3516), .B2(\registers[8][8] ), 
        .ZN(n1464) );
  INV_X1 U2616 ( .A(n1465), .ZN(n3775) );
  AOI22_X1 U2617 ( .A1(n282), .A2(n277), .B1(n3516), .B2(\registers[8][9] ), 
        .ZN(n1465) );
  INV_X1 U2618 ( .A(n1188), .ZN(n4117) );
  AOI22_X1 U2619 ( .A1(n782), .A2(n14), .B1(n3593), .B2(\registers[24][8] ), 
        .ZN(n1188) );
  INV_X1 U2620 ( .A(n1189), .ZN(n4118) );
  AOI22_X1 U2621 ( .A1(n282), .A2(n3588), .B1(n3592), .B2(\registers[24][9] ), 
        .ZN(n1189) );
  INV_X1 U2622 ( .A(n1073), .ZN(n4202) );
  AOI22_X1 U2623 ( .A1(n388), .A2(n16), .B1(n3635), .B2(\registers[29][0] ), 
        .ZN(n1073) );
  INV_X1 U2624 ( .A(n1075), .ZN(n4203) );
  AOI22_X1 U2625 ( .A1(n902), .A2(n690), .B1(n3638), .B2(\registers[29][1] ), 
        .ZN(n1075) );
  INV_X1 U2626 ( .A(n1076), .ZN(n4204) );
  AOI22_X1 U2627 ( .A1(n189), .A2(n763), .B1(n3637), .B2(\registers[29][2] ), 
        .ZN(n1076) );
  INV_X1 U2628 ( .A(n1107), .ZN(n4171) );
  AOI22_X1 U2629 ( .A1(n387), .A2(n689), .B1(n3627), .B2(\registers[28][0] ), 
        .ZN(n1107) );
  INV_X1 U2630 ( .A(n1109), .ZN(n4172) );
  AOI22_X1 U2631 ( .A1(n279), .A2(n767), .B1(n3628), .B2(\registers[28][1] ), 
        .ZN(n1109) );
  INV_X1 U2632 ( .A(n1110), .ZN(n4173) );
  AOI22_X1 U2633 ( .A1(n900), .A2(n767), .B1(n3626), .B2(\registers[28][2] ), 
        .ZN(n1110) );
  INV_X1 U2634 ( .A(n1145), .ZN(n4139) );
  AOI22_X1 U2635 ( .A1(n388), .A2(n777), .B1(n13), .B2(\registers[25][0] ), 
        .ZN(n1145) );
  INV_X1 U2636 ( .A(n1147), .ZN(n4140) );
  AOI22_X1 U2637 ( .A1(n902), .A2(n777), .B1(n3598), .B2(\registers[25][1] ), 
        .ZN(n1147) );
  INV_X1 U2638 ( .A(n1148), .ZN(n4141) );
  AOI22_X1 U2639 ( .A1(n190), .A2(n778), .B1(n234), .B2(\registers[25][2] ), 
        .ZN(n1148) );
  INV_X1 U2640 ( .A(n1179), .ZN(n4109) );
  AOI22_X1 U2641 ( .A1(n904), .A2(n3590), .B1(n3593), .B2(\registers[24][0] ), 
        .ZN(n1179) );
  INV_X1 U2642 ( .A(n1181), .ZN(n4110) );
  AOI22_X1 U2643 ( .A1(n279), .A2(n171), .B1(n3592), .B2(\registers[24][1] ), 
        .ZN(n1181) );
  INV_X1 U2644 ( .A(n1182), .ZN(n4111) );
  AOI22_X1 U2645 ( .A1(n900), .A2(n3588), .B1(n3591), .B2(\registers[24][2] ), 
        .ZN(n1182) );
  INV_X1 U2646 ( .A(n1214), .ZN(n4078) );
  AOI22_X1 U2647 ( .A1(n387), .A2(n765), .B1(n3584), .B2(\registers[23][0] ), 
        .ZN(n1214) );
  INV_X1 U2648 ( .A(n1216), .ZN(n4079) );
  AOI22_X1 U2649 ( .A1(n902), .A2(n765), .B1(n3585), .B2(\registers[23][1] ), 
        .ZN(n1216) );
  INV_X1 U2650 ( .A(n1217), .ZN(n4080) );
  AOI22_X1 U2651 ( .A1(n189), .A2(n765), .B1(n3583), .B2(\registers[23][2] ), 
        .ZN(n1217) );
  INV_X1 U2652 ( .A(n1248), .ZN(n4050) );
  AOI22_X1 U2653 ( .A1(n387), .A2(n25), .B1(net44860), .B2(\registers[22][0] ), 
        .ZN(n1248) );
  INV_X1 U2654 ( .A(n1250), .ZN(n4051) );
  AOI22_X1 U2655 ( .A1(n279), .A2(net44303), .B1(net44604), .B2(
        \registers[22][1] ), .ZN(n1250) );
  INV_X1 U2656 ( .A(n1251), .ZN(n4052) );
  AOI22_X1 U2657 ( .A1(n189), .A2(net26247), .B1(n20), .B2(\registers[22][2] ), 
        .ZN(n1251) );
  INV_X1 U2658 ( .A(n1283), .ZN(n4018) );
  AOI22_X1 U2659 ( .A1(n388), .A2(n761), .B1(n3), .B2(\registers[19][0] ), 
        .ZN(n1283) );
  INV_X1 U2660 ( .A(n1285), .ZN(n4019) );
  AOI22_X1 U2661 ( .A1(n279), .A2(n3570), .B1(n3571), .B2(\registers[19][1] ), 
        .ZN(n1285) );
  INV_X1 U2662 ( .A(n1286), .ZN(n4020) );
  AOI22_X1 U2663 ( .A1(n189), .A2(n3569), .B1(n3572), .B2(\registers[19][2] ), 
        .ZN(n1286) );
  INV_X1 U2664 ( .A(n1316), .ZN(n3986) );
  AOI22_X1 U2665 ( .A1(n904), .A2(n3564), .B1(n3565), .B2(\registers[18][0] ), 
        .ZN(n1316) );
  INV_X1 U2666 ( .A(n1318), .ZN(n3987) );
  AOI22_X1 U2667 ( .A1(n902), .A2(n3564), .B1(n3565), .B2(\registers[18][1] ), 
        .ZN(n1318) );
  INV_X1 U2668 ( .A(n1319), .ZN(n3988) );
  AOI22_X1 U2669 ( .A1(n190), .A2(n3562), .B1(n3565), .B2(\registers[18][2] ), 
        .ZN(n1319) );
  INV_X1 U2670 ( .A(n1354), .ZN(n3859) );
  AOI22_X1 U2671 ( .A1(n387), .A2(n3546), .B1(n216), .B2(\registers[13][0] ), 
        .ZN(n1354) );
  INV_X1 U2672 ( .A(n1356), .ZN(n3860) );
  AOI22_X1 U2673 ( .A1(n279), .A2(n776), .B1(n216), .B2(\registers[13][1] ), 
        .ZN(n1356) );
  INV_X1 U2674 ( .A(n1357), .ZN(n3861) );
  AOI22_X1 U2675 ( .A1(n190), .A2(n776), .B1(n216), .B2(\registers[13][2] ), 
        .ZN(n1357) );
  INV_X1 U2676 ( .A(n1387), .ZN(n3828) );
  AOI22_X1 U2677 ( .A1(n388), .A2(n204), .B1(n3540), .B2(\registers[12][0] ), 
        .ZN(n1387) );
  INV_X1 U2678 ( .A(n1389), .ZN(n3829) );
  AOI22_X1 U2679 ( .A1(n902), .A2(n692), .B1(n3542), .B2(\registers[12][1] ), 
        .ZN(n1389) );
  INV_X1 U2680 ( .A(n1390), .ZN(n3830) );
  AOI22_X1 U2681 ( .A1(n190), .A2(n204), .B1(n3539), .B2(\registers[12][2] ), 
        .ZN(n1390) );
  INV_X1 U2682 ( .A(n1422), .ZN(n3797) );
  AOI22_X1 U2683 ( .A1(n904), .A2(n774), .B1(n3521), .B2(\registers[9][0] ), 
        .ZN(n1422) );
  INV_X1 U2684 ( .A(n1424), .ZN(n3798) );
  AOI22_X1 U2685 ( .A1(n279), .A2(n774), .B1(n3523), .B2(\registers[9][1] ), 
        .ZN(n1424) );
  INV_X1 U2686 ( .A(n1425), .ZN(n3799) );
  AOI22_X1 U2687 ( .A1(n190), .A2(n679), .B1(n3525), .B2(\registers[9][2] ), 
        .ZN(n1425) );
  INV_X1 U2688 ( .A(n1455), .ZN(n3766) );
  AOI22_X1 U2689 ( .A1(n904), .A2(n3513), .B1(n3516), .B2(\registers[8][0] ), 
        .ZN(n1455) );
  INV_X1 U2690 ( .A(n1457), .ZN(n3767) );
  AOI22_X1 U2691 ( .A1(n902), .A2(n389), .B1(n3514), .B2(\registers[8][1] ), 
        .ZN(n1457) );
  INV_X1 U2692 ( .A(n1458), .ZN(n3768) );
  AOI22_X1 U2693 ( .A1(n189), .A2(n390), .B1(n3516), .B2(\registers[8][2] ), 
        .ZN(n1458) );
  INV_X1 U2694 ( .A(n1488), .ZN(n3953) );
  AOI22_X1 U2695 ( .A1(n388), .A2(n214), .B1(n3510), .B2(\registers[7][0] ), 
        .ZN(n1488) );
  INV_X1 U2696 ( .A(n1490), .ZN(n3954) );
  AOI22_X1 U2697 ( .A1(n902), .A2(n214), .B1(n3509), .B2(\registers[7][1] ), 
        .ZN(n1490) );
  INV_X1 U2698 ( .A(n1491), .ZN(n3955) );
  AOI22_X1 U2699 ( .A1(n900), .A2(n3505), .B1(n3508), .B2(\registers[7][2] ), 
        .ZN(n1491) );
  INV_X1 U2700 ( .A(n1522), .ZN(n3922) );
  AOI22_X1 U2701 ( .A1(n387), .A2(net26583), .B1(net26585), .B2(
        \registers[6][0] ), .ZN(n1522) );
  INV_X1 U2702 ( .A(n1524), .ZN(n3923) );
  AOI22_X1 U2703 ( .A1(net39089), .A2(n279), .B1(net26595), .B2(
        \registers[6][1] ), .ZN(n1524) );
  INV_X1 U2704 ( .A(n1525), .ZN(n3924) );
  AOI22_X1 U2705 ( .A1(n190), .A2(net26581), .B1(net26589), .B2(
        \registers[6][2] ), .ZN(n1525) );
  INV_X1 U2706 ( .A(n1559), .ZN(n3890) );
  AOI22_X1 U2707 ( .A1(n904), .A2(n3494), .B1(n3497), .B2(\registers[1][0] ), 
        .ZN(n1559) );
  INV_X1 U2708 ( .A(n1561), .ZN(n3891) );
  AOI22_X1 U2709 ( .A1(n902), .A2(n3494), .B1(n3500), .B2(\registers[1][1] ), 
        .ZN(n1561) );
  INV_X1 U2710 ( .A(n1562), .ZN(n3892) );
  AOI22_X1 U2711 ( .A1(n189), .A2(n3493), .B1(n3497), .B2(\registers[1][2] ), 
        .ZN(n1562) );
  INV_X1 U2712 ( .A(n1320), .ZN(n3989) );
  AOI22_X1 U2713 ( .A1(n249), .A2(n3563), .B1(n3565), .B2(\registers[18][3] ), 
        .ZN(n1320) );
  INV_X1 U2714 ( .A(n1321), .ZN(n3990) );
  AOI22_X1 U2715 ( .A1(n267), .A2(n595), .B1(n3566), .B2(\registers[18][4] ), 
        .ZN(n1321) );
  INV_X1 U2716 ( .A(n1322), .ZN(n3991) );
  AOI22_X1 U2717 ( .A1(n412), .A2(n595), .B1(n3565), .B2(\registers[18][5] ), 
        .ZN(n1322) );
  INV_X1 U2718 ( .A(n1323), .ZN(n3992) );
  AOI22_X1 U2719 ( .A1(n795), .A2(n3564), .B1(n3566), .B2(\registers[18][6] ), 
        .ZN(n1323) );
  INV_X1 U2720 ( .A(n1324), .ZN(n3993) );
  AOI22_X1 U2721 ( .A1(n211), .A2(n3563), .B1(n3565), .B2(\registers[18][7] ), 
        .ZN(n1324) );
  INV_X1 U2722 ( .A(n1287), .ZN(n4021) );
  AOI22_X1 U2723 ( .A1(n249), .A2(n3569), .B1(n3573), .B2(\registers[19][3] ), 
        .ZN(n1287) );
  INV_X1 U2724 ( .A(n1288), .ZN(n4022) );
  AOI22_X1 U2725 ( .A1(n163), .A2(n3570), .B1(n3572), .B2(\registers[19][4] ), 
        .ZN(n1288) );
  INV_X1 U2726 ( .A(n1289), .ZN(n4023) );
  AOI22_X1 U2727 ( .A1(n787), .A2(n577), .B1(n3573), .B2(\registers[19][5] ), 
        .ZN(n1289) );
  INV_X1 U2728 ( .A(n1290), .ZN(n4024) );
  AOI22_X1 U2729 ( .A1(n278), .A2(n3568), .B1(n31), .B2(\registers[19][6] ), 
        .ZN(n1290) );
  INV_X1 U2730 ( .A(n1291), .ZN(n4025) );
  AOI22_X1 U2731 ( .A1(n162), .A2(n577), .B1(n3572), .B2(\registers[19][7] ), 
        .ZN(n1291) );
  INV_X1 U2732 ( .A(n1149), .ZN(n4142) );
  AOI22_X1 U2733 ( .A1(n167), .A2(n3596), .B1(n234), .B2(\registers[25][3] ), 
        .ZN(n1149) );
  INV_X1 U2734 ( .A(n1150), .ZN(n4143) );
  AOI22_X1 U2735 ( .A1(n789), .A2(n736), .B1(n3602), .B2(\registers[25][4] ), 
        .ZN(n1150) );
  INV_X1 U2736 ( .A(n1151), .ZN(n4144) );
  AOI22_X1 U2737 ( .A1(n413), .A2(n736), .B1(n3601), .B2(\registers[25][5] ), 
        .ZN(n1151) );
  INV_X1 U2738 ( .A(n1152), .ZN(n4145) );
  AOI22_X1 U2739 ( .A1(n278), .A2(n3595), .B1(n234), .B2(\registers[25][6] ), 
        .ZN(n1152) );
  INV_X1 U2740 ( .A(n1153), .ZN(n4146) );
  AOI22_X1 U2741 ( .A1(n211), .A2(n3596), .B1(n3598), .B2(\registers[25][7] ), 
        .ZN(n1153) );
  INV_X1 U2742 ( .A(n1358), .ZN(n3862) );
  AOI22_X1 U2743 ( .A1(n167), .A2(n196), .B1(n215), .B2(\registers[13][3] ), 
        .ZN(n1358) );
  INV_X1 U2744 ( .A(n1359), .ZN(n3863) );
  AOI22_X1 U2745 ( .A1(n789), .A2(n776), .B1(n216), .B2(\registers[13][4] ), 
        .ZN(n1359) );
  INV_X1 U2746 ( .A(n1360), .ZN(n3864) );
  AOI22_X1 U2747 ( .A1(n413), .A2(n776), .B1(n219), .B2(\registers[13][5] ), 
        .ZN(n1360) );
  INV_X1 U2748 ( .A(n1361), .ZN(n3865) );
  AOI22_X1 U2749 ( .A1(n795), .A2(n775), .B1(n17), .B2(\registers[13][6] ), 
        .ZN(n1361) );
  INV_X1 U2750 ( .A(n1362), .ZN(n3866) );
  AOI22_X1 U2751 ( .A1(n793), .A2(n3546), .B1(n17), .B2(\registers[13][7] ), 
        .ZN(n1362) );
  INV_X1 U2752 ( .A(n1391), .ZN(n3831) );
  AOI22_X1 U2753 ( .A1(n791), .A2(n692), .B1(n3541), .B2(\registers[12][3] ), 
        .ZN(n1391) );
  INV_X1 U2754 ( .A(n1392), .ZN(n3832) );
  AOI22_X1 U2755 ( .A1(n789), .A2(n204), .B1(n3540), .B2(\registers[12][4] ), 
        .ZN(n1392) );
  INV_X1 U2756 ( .A(n1393), .ZN(n3833) );
  AOI22_X1 U2757 ( .A1(n787), .A2(n770), .B1(n3542), .B2(\registers[12][5] ), 
        .ZN(n1393) );
  INV_X1 U2758 ( .A(n1394), .ZN(n3834) );
  AOI22_X1 U2759 ( .A1(n795), .A2(n3537), .B1(n3539), .B2(\registers[12][6] ), 
        .ZN(n1394) );
  INV_X1 U2760 ( .A(n1395), .ZN(n3835) );
  AOI22_X1 U2761 ( .A1(n162), .A2(n693), .B1(n3542), .B2(\registers[12][7] ), 
        .ZN(n1395) );
  INV_X1 U2762 ( .A(n1077), .ZN(n4205) );
  AOI22_X1 U2763 ( .A1(n791), .A2(n691), .B1(n3636), .B2(\registers[29][3] ), 
        .ZN(n1077) );
  INV_X1 U2764 ( .A(n1078), .ZN(n4206) );
  AOI22_X1 U2765 ( .A1(n267), .A2(n691), .B1(n3636), .B2(\registers[29][4] ), 
        .ZN(n1078) );
  INV_X1 U2766 ( .A(n1079), .ZN(n4207) );
  AOI22_X1 U2767 ( .A1(n413), .A2(n3632), .B1(n3637), .B2(\registers[29][5] ), 
        .ZN(n1079) );
  INV_X1 U2768 ( .A(n1080), .ZN(n4208) );
  AOI22_X1 U2769 ( .A1(n795), .A2(n3633), .B1(n3637), .B2(\registers[29][6] ), 
        .ZN(n1080) );
  INV_X1 U2770 ( .A(n1081), .ZN(n4209) );
  AOI22_X1 U2771 ( .A1(n211), .A2(n3634), .B1(n3636), .B2(\registers[29][7] ), 
        .ZN(n1081) );
  INV_X1 U2772 ( .A(n1111), .ZN(n4174) );
  AOI22_X1 U2773 ( .A1(n167), .A2(n3625), .B1(n3629), .B2(\registers[28][3] ), 
        .ZN(n1111) );
  INV_X1 U2774 ( .A(n1112), .ZN(n4175) );
  AOI22_X1 U2775 ( .A1(n267), .A2(n3625), .B1(n3630), .B2(\registers[28][4] ), 
        .ZN(n1112) );
  INV_X1 U2776 ( .A(n1113), .ZN(n4176) );
  AOI22_X1 U2777 ( .A1(n412), .A2(n3623), .B1(n3626), .B2(\registers[28][5] ), 
        .ZN(n1113) );
  INV_X1 U2778 ( .A(n1114), .ZN(n4177) );
  AOI22_X1 U2779 ( .A1(n278), .A2(n768), .B1(n3626), .B2(\registers[28][6] ), 
        .ZN(n1114) );
  INV_X1 U2780 ( .A(n1219), .ZN(n4081) );
  AOI22_X1 U2781 ( .A1(n789), .A2(n3580), .B1(n3585), .B2(\registers[23][4] ), 
        .ZN(n1219) );
  INV_X1 U2782 ( .A(n1220), .ZN(n4082) );
  AOI22_X1 U2783 ( .A1(n787), .A2(n3581), .B1(n3586), .B2(\registers[23][5] ), 
        .ZN(n1220) );
  INV_X1 U2784 ( .A(n1221), .ZN(n4083) );
  AOI22_X1 U2785 ( .A1(n278), .A2(n206), .B1(n3584), .B2(\registers[23][6] ), 
        .ZN(n1221) );
  INV_X1 U2786 ( .A(n1222), .ZN(n4084) );
  AOI22_X1 U2787 ( .A1(n793), .A2(n206), .B1(n3585), .B2(\registers[23][7] ), 
        .ZN(n1222) );
  INV_X1 U2788 ( .A(n1492), .ZN(n3956) );
  AOI22_X1 U2789 ( .A1(n167), .A2(n214), .B1(n3509), .B2(\registers[7][3] ), 
        .ZN(n1492) );
  INV_X1 U2790 ( .A(n1493), .ZN(n3957) );
  AOI22_X1 U2791 ( .A1(n163), .A2(n683), .B1(n3510), .B2(\registers[7][4] ), 
        .ZN(n1493) );
  INV_X1 U2792 ( .A(n1494), .ZN(n3958) );
  AOI22_X1 U2793 ( .A1(n413), .A2(n213), .B1(n3508), .B2(\registers[7][5] ), 
        .ZN(n1494) );
  INV_X1 U2794 ( .A(n1495), .ZN(n3959) );
  AOI22_X1 U2795 ( .A1(n795), .A2(n3506), .B1(n3509), .B2(\registers[7][6] ), 
        .ZN(n1495) );
  INV_X1 U2796 ( .A(n1496), .ZN(n3960) );
  AOI22_X1 U2797 ( .A1(n162), .A2(n683), .B1(n3510), .B2(\registers[7][7] ), 
        .ZN(n1496) );
  INV_X1 U2798 ( .A(n1426), .ZN(n3800) );
  AOI22_X1 U2799 ( .A1(n167), .A2(n679), .B1(n3524), .B2(\registers[9][3] ), 
        .ZN(n1426) );
  INV_X1 U2800 ( .A(n1427), .ZN(n3801) );
  AOI22_X1 U2801 ( .A1(n163), .A2(n773), .B1(n3524), .B2(\registers[9][4] ), 
        .ZN(n1427) );
  INV_X1 U2802 ( .A(n1428), .ZN(n3802) );
  AOI22_X1 U2803 ( .A1(n412), .A2(n679), .B1(n3521), .B2(\registers[9][5] ), 
        .ZN(n1428) );
  INV_X1 U2804 ( .A(n1429), .ZN(n3803) );
  AOI22_X1 U2805 ( .A1(n278), .A2(n3519), .B1(n3522), .B2(\registers[9][6] ), 
        .ZN(n1429) );
  INV_X1 U2806 ( .A(n1430), .ZN(n3804) );
  AOI22_X1 U2807 ( .A1(n211), .A2(n3518), .B1(n3523), .B2(\registers[9][7] ), 
        .ZN(n1430) );
  INV_X1 U2808 ( .A(n1563), .ZN(n3893) );
  AOI22_X1 U2809 ( .A1(n249), .A2(n771), .B1(n3496), .B2(\registers[1][3] ), 
        .ZN(n1563) );
  INV_X1 U2810 ( .A(n1564), .ZN(n3894) );
  AOI22_X1 U2811 ( .A1(n163), .A2(n677), .B1(n3496), .B2(\registers[1][4] ), 
        .ZN(n1564) );
  INV_X1 U2812 ( .A(n1565), .ZN(n3895) );
  AOI22_X1 U2813 ( .A1(n787), .A2(n677), .B1(n3495), .B2(\registers[1][5] ), 
        .ZN(n1565) );
  INV_X1 U2814 ( .A(n1566), .ZN(n3896) );
  AOI22_X1 U2815 ( .A1(n278), .A2(n3494), .B1(n3500), .B2(\registers[1][6] ), 
        .ZN(n1566) );
  INV_X1 U2816 ( .A(n1567), .ZN(n3897) );
  AOI22_X1 U2817 ( .A1(n211), .A2(n3492), .B1(n3495), .B2(\registers[1][7] ), 
        .ZN(n1567) );
  INV_X1 U2818 ( .A(n1252), .ZN(n4053) );
  AOI22_X1 U2819 ( .A1(n249), .A2(net26247), .B1(net44322), .B2(
        \registers[22][3] ), .ZN(n1252) );
  INV_X1 U2820 ( .A(n1253), .ZN(n4054) );
  AOI22_X1 U2821 ( .A1(n789), .A2(n25), .B1(n241), .B2(\registers[22][4] ), 
        .ZN(n1253) );
  INV_X1 U2822 ( .A(n1254), .ZN(n4055) );
  AOI22_X1 U2823 ( .A1(n413), .A2(net26243), .B1(net44605), .B2(
        \registers[22][5] ), .ZN(n1254) );
  INV_X1 U2824 ( .A(n1255), .ZN(n4056) );
  AOI22_X1 U2825 ( .A1(n795), .A2(net44304), .B1(net44605), .B2(
        \registers[22][6] ), .ZN(n1255) );
  INV_X1 U2826 ( .A(n1256), .ZN(n4057) );
  AOI22_X1 U2827 ( .A1(n162), .A2(net44304), .B1(net44605), .B2(
        \registers[22][7] ), .ZN(n1256) );
  INV_X1 U2828 ( .A(n1526), .ZN(n3925) );
  AOI22_X1 U2829 ( .A1(n249), .A2(net38993), .B1(net26593), .B2(
        \registers[6][3] ), .ZN(n1526) );
  INV_X1 U2830 ( .A(n1527), .ZN(n3926) );
  AOI22_X1 U2831 ( .A1(n267), .A2(net39090), .B1(net26589), .B2(
        \registers[6][4] ), .ZN(n1527) );
  INV_X1 U2832 ( .A(n1528), .ZN(n3927) );
  AOI22_X1 U2833 ( .A1(n413), .A2(net26583), .B1(net26595), .B2(
        \registers[6][5] ), .ZN(n1528) );
  INV_X1 U2834 ( .A(n1529), .ZN(n3928) );
  AOI22_X1 U2835 ( .A1(n229), .A2(n795), .B1(net26585), .B2(\registers[6][6] ), 
        .ZN(n1529) );
  INV_X1 U2836 ( .A(n1530), .ZN(n3929) );
  AOI22_X1 U2837 ( .A1(n793), .A2(net26579), .B1(net26589), .B2(
        \registers[6][7] ), .ZN(n1530) );
  INV_X1 U2838 ( .A(n1459), .ZN(n3769) );
  AOI22_X1 U2839 ( .A1(n167), .A2(n3512), .B1(n3516), .B2(\registers[8][3] ), 
        .ZN(n1459) );
  INV_X1 U2840 ( .A(n1460), .ZN(n3770) );
  AOI22_X1 U2841 ( .A1(n789), .A2(n3513), .B1(n3516), .B2(\registers[8][4] ), 
        .ZN(n1460) );
  INV_X1 U2842 ( .A(n1461), .ZN(n3771) );
  AOI22_X1 U2843 ( .A1(n412), .A2(n390), .B1(n3515), .B2(\registers[8][5] ), 
        .ZN(n1461) );
  INV_X1 U2844 ( .A(n1462), .ZN(n3772) );
  AOI22_X1 U2845 ( .A1(n795), .A2(n277), .B1(n3514), .B2(\registers[8][6] ), 
        .ZN(n1462) );
  INV_X1 U2846 ( .A(n1463), .ZN(n3773) );
  AOI22_X1 U2847 ( .A1(n211), .A2(n390), .B1(n3516), .B2(\registers[8][7] ), 
        .ZN(n1463) );
  INV_X1 U2848 ( .A(n1183), .ZN(n4112) );
  AOI22_X1 U2849 ( .A1(n791), .A2(n3589), .B1(n3592), .B2(\registers[24][3] ), 
        .ZN(n1183) );
  INV_X1 U2850 ( .A(n1184), .ZN(n4113) );
  AOI22_X1 U2851 ( .A1(n267), .A2(n3588), .B1(n3591), .B2(\registers[24][4] ), 
        .ZN(n1184) );
  INV_X1 U2852 ( .A(n1185), .ZN(n4114) );
  AOI22_X1 U2853 ( .A1(n787), .A2(n3588), .B1(n3592), .B2(\registers[24][5] ), 
        .ZN(n1185) );
  INV_X1 U2854 ( .A(n1186), .ZN(n4115) );
  AOI22_X1 U2855 ( .A1(n278), .A2(n3588), .B1(n3591), .B2(\registers[24][6] ), 
        .ZN(n1186) );
  INV_X1 U2856 ( .A(n1187), .ZN(n4116) );
  AOI22_X1 U2857 ( .A1(n793), .A2(n14), .B1(n3592), .B2(\registers[24][7] ), 
        .ZN(n1187) );
  INV_X1 U2858 ( .A(n1084), .ZN(n4212) );
  AOI22_X1 U2859 ( .A1(n283), .A2(n762), .B1(n3636), .B2(\registers[29][10] ), 
        .ZN(n1084) );
  INV_X1 U2860 ( .A(n1085), .ZN(n4213) );
  AOI22_X1 U2861 ( .A1(n548), .A2(n763), .B1(n3638), .B2(\registers[29][11] ), 
        .ZN(n1085) );
  INV_X1 U2862 ( .A(n1086), .ZN(n4214) );
  AOI22_X1 U2863 ( .A1(n166), .A2(n16), .B1(n3638), .B2(\registers[29][12] ), 
        .ZN(n1086) );
  INV_X1 U2864 ( .A(n1087), .ZN(n4215) );
  AOI22_X1 U2865 ( .A1(n284), .A2(n763), .B1(n3637), .B2(\registers[29][13] ), 
        .ZN(n1087) );
  INV_X1 U2866 ( .A(n1088), .ZN(n4216) );
  AOI22_X1 U2867 ( .A1(n894), .A2(n3632), .B1(n3638), .B2(\registers[29][14] ), 
        .ZN(n1088) );
  INV_X1 U2868 ( .A(n1089), .ZN(n4217) );
  AOI22_X1 U2869 ( .A1(n892), .A2(n691), .B1(n3637), .B2(\registers[29][15] ), 
        .ZN(n1089) );
  INV_X1 U2870 ( .A(n1090), .ZN(n4218) );
  AOI22_X1 U2871 ( .A1(n890), .A2(n3632), .B1(n3636), .B2(\registers[29][16] ), 
        .ZN(n1090) );
  INV_X1 U2872 ( .A(n1091), .ZN(n4219) );
  AOI22_X1 U2873 ( .A1(n250), .A2(n3632), .B1(n3637), .B2(\registers[29][17] ), 
        .ZN(n1091) );
  INV_X1 U2874 ( .A(n1092), .ZN(n4220) );
  AOI22_X1 U2875 ( .A1(n886), .A2(n762), .B1(n3635), .B2(\registers[29][18] ), 
        .ZN(n1092) );
  INV_X1 U2876 ( .A(n1093), .ZN(n4221) );
  AOI22_X1 U2877 ( .A1(n545), .A2(n763), .B1(n3638), .B2(\registers[29][19] ), 
        .ZN(n1093) );
  INV_X1 U2878 ( .A(n1094), .ZN(n4222) );
  AOI22_X1 U2879 ( .A1(n161), .A2(n3634), .B1(n3636), .B2(\registers[29][20] ), 
        .ZN(n1094) );
  INV_X1 U2880 ( .A(n1095), .ZN(n4223) );
  AOI22_X1 U2881 ( .A1(n880), .A2(n691), .B1(n3638), .B2(\registers[29][21] ), 
        .ZN(n1095) );
  INV_X1 U2882 ( .A(n1096), .ZN(n4224) );
  AOI22_X1 U2883 ( .A1(n877), .A2(n16), .B1(n3637), .B2(\registers[29][22] ), 
        .ZN(n1096) );
  INV_X1 U2884 ( .A(n1097), .ZN(n4225) );
  AOI22_X1 U2885 ( .A1(n264), .A2(n3633), .B1(n3638), .B2(\registers[29][23] ), 
        .ZN(n1097) );
  INV_X1 U2886 ( .A(n1099), .ZN(n4226) );
  AOI22_X1 U2887 ( .A1(n200), .A2(n762), .B1(n3636), .B2(\registers[29][25] ), 
        .ZN(n1099) );
  INV_X1 U2888 ( .A(n1100), .ZN(n4227) );
  AOI22_X1 U2889 ( .A1(n870), .A2(n16), .B1(n3635), .B2(\registers[29][26] ), 
        .ZN(n1100) );
  INV_X1 U2890 ( .A(n1101), .ZN(n4228) );
  AOI22_X1 U2891 ( .A1(n557), .A2(n762), .B1(n3638), .B2(\registers[29][27] ), 
        .ZN(n1101) );
  INV_X1 U2892 ( .A(n1102), .ZN(n4229) );
  AOI22_X1 U2893 ( .A1(net28529), .A2(n690), .B1(n3636), .B2(
        \registers[29][28] ), .ZN(n1102) );
  INV_X1 U2894 ( .A(n1103), .ZN(n4230) );
  AOI22_X1 U2895 ( .A1(n230), .A2(n690), .B1(n3636), .B2(\registers[29][29] ), 
        .ZN(n1103) );
  INV_X1 U2896 ( .A(n1104), .ZN(n4231) );
  AOI22_X1 U2897 ( .A1(n395), .A2(n690), .B1(n3636), .B2(\registers[29][30] ), 
        .ZN(n1104) );
  INV_X1 U2898 ( .A(n1118), .ZN(n4180) );
  AOI22_X1 U2899 ( .A1(n799), .A2(n689), .B1(n3627), .B2(\registers[28][10] ), 
        .ZN(n1118) );
  INV_X1 U2900 ( .A(n1119), .ZN(n4181) );
  AOI22_X1 U2901 ( .A1(n796), .A2(n768), .B1(n3627), .B2(\registers[28][11] ), 
        .ZN(n1119) );
  INV_X1 U2902 ( .A(n1120), .ZN(n4182) );
  AOI22_X1 U2903 ( .A1(n165), .A2(n3624), .B1(n3627), .B2(\registers[28][12] ), 
        .ZN(n1120) );
  INV_X1 U2904 ( .A(n1121), .ZN(n4183) );
  AOI22_X1 U2905 ( .A1(n896), .A2(n3624), .B1(n3627), .B2(\registers[28][13] ), 
        .ZN(n1121) );
  INV_X1 U2906 ( .A(n1122), .ZN(n4184) );
  AOI22_X1 U2907 ( .A1(n223), .A2(n3625), .B1(n3627), .B2(\registers[28][14] ), 
        .ZN(n1122) );
  INV_X1 U2908 ( .A(n1123), .ZN(n4185) );
  AOI22_X1 U2909 ( .A1(n892), .A2(n3623), .B1(n3628), .B2(\registers[28][15] ), 
        .ZN(n1123) );
  INV_X1 U2910 ( .A(n1124), .ZN(n4186) );
  AOI22_X1 U2911 ( .A1(n262), .A2(n3623), .B1(n3628), .B2(\registers[28][16] ), 
        .ZN(n1124) );
  INV_X1 U2912 ( .A(n1125), .ZN(n4187) );
  AOI22_X1 U2913 ( .A1(n250), .A2(n3623), .B1(n3628), .B2(\registers[28][17] ), 
        .ZN(n1125) );
  INV_X1 U2914 ( .A(n1126), .ZN(n4188) );
  AOI22_X1 U2915 ( .A1(n259), .A2(n3624), .B1(n3628), .B2(\registers[28][18] ), 
        .ZN(n1126) );
  INV_X1 U2916 ( .A(n1127), .ZN(n4189) );
  AOI22_X1 U2917 ( .A1(n883), .A2(n689), .B1(n3628), .B2(\registers[28][19] ), 
        .ZN(n1127) );
  INV_X1 U2918 ( .A(n1128), .ZN(n4190) );
  AOI22_X1 U2919 ( .A1(n207), .A2(n3624), .B1(n3629), .B2(\registers[28][20] ), 
        .ZN(n1128) );
  INV_X1 U2920 ( .A(n1129), .ZN(n4191) );
  AOI22_X1 U2921 ( .A1(n880), .A2(n768), .B1(n3629), .B2(\registers[28][21] ), 
        .ZN(n1129) );
  INV_X1 U2922 ( .A(n1130), .ZN(n4192) );
  AOI22_X1 U2923 ( .A1(n19), .A2(n688), .B1(n3629), .B2(\registers[28][22] ), 
        .ZN(n1130) );
  INV_X1 U2924 ( .A(n1131), .ZN(n4193) );
  AOI22_X1 U2925 ( .A1(n876), .A2(n3624), .B1(n3629), .B2(\registers[28][23] ), 
        .ZN(n1131) );
  INV_X1 U2926 ( .A(n1132), .ZN(n4194) );
  AOI22_X1 U2927 ( .A1(n398), .A2(n767), .B1(n3629), .B2(\registers[28][24] ), 
        .ZN(n1132) );
  INV_X1 U2928 ( .A(n1133), .ZN(n4195) );
  AOI22_X1 U2929 ( .A1(n872), .A2(n688), .B1(n3630), .B2(\registers[28][25] ), 
        .ZN(n1133) );
  INV_X1 U2930 ( .A(n1134), .ZN(n4196) );
  AOI22_X1 U2931 ( .A1(n559), .A2(n3623), .B1(n3630), .B2(\registers[28][26] ), 
        .ZN(n1134) );
  INV_X1 U2932 ( .A(n1135), .ZN(n4197) );
  AOI22_X1 U2933 ( .A1(n868), .A2(n689), .B1(n3630), .B2(\registers[28][27] ), 
        .ZN(n1135) );
  INV_X1 U2934 ( .A(n1136), .ZN(n4198) );
  AOI22_X1 U2935 ( .A1(n246), .A2(n3625), .B1(n3630), .B2(\registers[28][28] ), 
        .ZN(n1136) );
  INV_X1 U2936 ( .A(n1137), .ZN(n4199) );
  AOI22_X1 U2937 ( .A1(n866), .A2(n768), .B1(n3630), .B2(\registers[28][29] ), 
        .ZN(n1137) );
  INV_X1 U2938 ( .A(n1138), .ZN(n4200) );
  AOI22_X1 U2939 ( .A1(n394), .A2(n688), .B1(n3631), .B2(\registers[28][30] ), 
        .ZN(n1138) );
  INV_X1 U2940 ( .A(n1156), .ZN(n4149) );
  AOI22_X1 U2941 ( .A1(n283), .A2(n736), .B1(n234), .B2(\registers[25][10] ), 
        .ZN(n1156) );
  INV_X1 U2942 ( .A(n1157), .ZN(n4150) );
  AOI22_X1 U2943 ( .A1(n548), .A2(n777), .B1(n3598), .B2(\registers[25][11] ), 
        .ZN(n1157) );
  INV_X1 U2944 ( .A(n1158), .ZN(n4151) );
  AOI22_X1 U2945 ( .A1(n898), .A2(n3597), .B1(n3603), .B2(\registers[25][12] ), 
        .ZN(n1158) );
  INV_X1 U2946 ( .A(n1159), .ZN(n4152) );
  AOI22_X1 U2947 ( .A1(n284), .A2(n778), .B1(n3598), .B2(\registers[25][13] ), 
        .ZN(n1159) );
  INV_X1 U2948 ( .A(n1160), .ZN(n4153) );
  AOI22_X1 U2949 ( .A1(n223), .A2(n3595), .B1(n3598), .B2(\registers[25][14] ), 
        .ZN(n1160) );
  INV_X1 U2950 ( .A(n1161), .ZN(n4154) );
  AOI22_X1 U2951 ( .A1(n210), .A2(n3596), .B1(n3602), .B2(\registers[25][15] ), 
        .ZN(n1161) );
  INV_X1 U2952 ( .A(n1162), .ZN(n4155) );
  AOI22_X1 U2953 ( .A1(n261), .A2(n3595), .B1(n3600), .B2(\registers[25][16] ), 
        .ZN(n1162) );
  INV_X1 U2954 ( .A(n1163), .ZN(n4156) );
  AOI22_X1 U2955 ( .A1(n888), .A2(n3595), .B1(n3602), .B2(\registers[25][17] ), 
        .ZN(n1163) );
  INV_X1 U2956 ( .A(n1164), .ZN(n4157) );
  AOI22_X1 U2957 ( .A1(n259), .A2(n737), .B1(n3599), .B2(\registers[25][18] ), 
        .ZN(n1164) );
  INV_X1 U2958 ( .A(n1165), .ZN(n4158) );
  AOI22_X1 U2959 ( .A1(n416), .A2(n3596), .B1(n234), .B2(\registers[25][19] ), 
        .ZN(n1165) );
  INV_X1 U2960 ( .A(n1166), .ZN(n4159) );
  AOI22_X1 U2961 ( .A1(n161), .A2(n778), .B1(n3601), .B2(\registers[25][20] ), 
        .ZN(n1166) );
  INV_X1 U2962 ( .A(n1167), .ZN(n4160) );
  AOI22_X1 U2963 ( .A1(n242), .A2(n778), .B1(n3603), .B2(\registers[25][21] ), 
        .ZN(n1167) );
  INV_X1 U2964 ( .A(n1168), .ZN(n4161) );
  AOI22_X1 U2965 ( .A1(n877), .A2(n3597), .B1(n3599), .B2(\registers[25][22] ), 
        .ZN(n1168) );
  INV_X1 U2966 ( .A(n1169), .ZN(n4162) );
  AOI22_X1 U2967 ( .A1(n264), .A2(n737), .B1(n3602), .B2(\registers[25][23] ), 
        .ZN(n1169) );
  INV_X1 U2968 ( .A(n1170), .ZN(n4163) );
  AOI22_X1 U2969 ( .A1(n410), .A2(n737), .B1(n3601), .B2(\registers[25][24] ), 
        .ZN(n1170) );
  INV_X1 U2970 ( .A(n1171), .ZN(n4164) );
  AOI22_X1 U2971 ( .A1(n200), .A2(n3597), .B1(n3602), .B2(\registers[25][25] ), 
        .ZN(n1171) );
  INV_X1 U2972 ( .A(n1172), .ZN(n4165) );
  AOI22_X1 U2973 ( .A1(n558), .A2(n777), .B1(n3599), .B2(\registers[25][26] ), 
        .ZN(n1172) );
  INV_X1 U2974 ( .A(n1173), .ZN(n4166) );
  AOI22_X1 U2975 ( .A1(n557), .A2(n3597), .B1(n3603), .B2(\registers[25][27] ), 
        .ZN(n1173) );
  INV_X1 U2976 ( .A(n1174), .ZN(n4167) );
  AOI22_X1 U2977 ( .A1(n246), .A2(n3597), .B1(n3600), .B2(\registers[25][28] ), 
        .ZN(n1174) );
  INV_X1 U2978 ( .A(n1175), .ZN(n4168) );
  AOI22_X1 U2979 ( .A1(n231), .A2(n737), .B1(n3600), .B2(\registers[25][29] ), 
        .ZN(n1175) );
  INV_X1 U2980 ( .A(n1176), .ZN(n4169) );
  AOI22_X1 U2981 ( .A1(n800), .A2(n736), .B1(n597), .B2(\registers[25][30] ), 
        .ZN(n1176) );
  INV_X1 U2982 ( .A(n1190), .ZN(n4119) );
  AOI22_X1 U2983 ( .A1(n799), .A2(n168), .B1(n3592), .B2(\registers[24][10] ), 
        .ZN(n1190) );
  INV_X1 U2984 ( .A(n1191), .ZN(n4120) );
  AOI22_X1 U2985 ( .A1(n549), .A2(n603), .B1(n3593), .B2(\registers[24][11] ), 
        .ZN(n1191) );
  INV_X1 U2986 ( .A(n1192), .ZN(n4121) );
  AOI22_X1 U2987 ( .A1(n166), .A2(n168), .B1(n3592), .B2(\registers[24][12] ), 
        .ZN(n1192) );
  INV_X1 U2988 ( .A(n1193), .ZN(n4122) );
  AOI22_X1 U2989 ( .A1(n896), .A2(n14), .B1(n3592), .B2(\registers[24][13] ), 
        .ZN(n1193) );
  INV_X1 U2990 ( .A(n1194), .ZN(n4123) );
  AOI22_X1 U2991 ( .A1(n894), .A2(n14), .B1(n3591), .B2(\registers[24][14] ), 
        .ZN(n1194) );
  INV_X1 U2992 ( .A(n1195), .ZN(n4124) );
  AOI22_X1 U2993 ( .A1(n210), .A2(n3590), .B1(n3592), .B2(\registers[24][15] ), 
        .ZN(n1195) );
  INV_X1 U2994 ( .A(n1196), .ZN(n4125) );
  AOI22_X1 U2995 ( .A1(n890), .A2(n171), .B1(n3592), .B2(\registers[24][16] ), 
        .ZN(n1196) );
  INV_X1 U2996 ( .A(n1197), .ZN(n4126) );
  AOI22_X1 U2997 ( .A1(n250), .A2(n3589), .B1(n3591), .B2(\registers[24][17] ), 
        .ZN(n1197) );
  INV_X1 U2998 ( .A(n1198), .ZN(n4127) );
  AOI22_X1 U2999 ( .A1(n886), .A2(n603), .B1(n3592), .B2(\registers[24][18] ), 
        .ZN(n1198) );
  INV_X1 U3000 ( .A(n1199), .ZN(n4128) );
  AOI22_X1 U3001 ( .A1(n883), .A2(n3590), .B1(n3593), .B2(\registers[24][19] ), 
        .ZN(n1199) );
  INV_X1 U3002 ( .A(n1200), .ZN(n4129) );
  AOI22_X1 U3003 ( .A1(n161), .A2(n3589), .B1(n3592), .B2(\registers[24][20] ), 
        .ZN(n1200) );
  INV_X1 U3004 ( .A(n1202), .ZN(n4130) );
  AOI22_X1 U3005 ( .A1(n245), .A2(n171), .B1(n3592), .B2(\registers[24][22] ), 
        .ZN(n1202) );
  INV_X1 U3006 ( .A(n1203), .ZN(n4131) );
  AOI22_X1 U3007 ( .A1(n265), .A2(n3589), .B1(n3592), .B2(\registers[24][23] ), 
        .ZN(n1203) );
  INV_X1 U3008 ( .A(n1205), .ZN(n4132) );
  AOI22_X1 U3009 ( .A1(n872), .A2(n603), .B1(n3593), .B2(\registers[24][25] ), 
        .ZN(n1205) );
  INV_X1 U3010 ( .A(n1206), .ZN(n4133) );
  AOI22_X1 U3011 ( .A1(n559), .A2(n168), .B1(n3592), .B2(\registers[24][26] ), 
        .ZN(n1206) );
  INV_X1 U3012 ( .A(n1207), .ZN(n4134) );
  AOI22_X1 U3013 ( .A1(n556), .A2(n3589), .B1(n3592), .B2(\registers[24][27] ), 
        .ZN(n1207) );
  INV_X1 U3014 ( .A(n1208), .ZN(n4135) );
  AOI22_X1 U3015 ( .A1(net28529), .A2(n3590), .B1(n3591), .B2(
        \registers[24][28] ), .ZN(n1208) );
  INV_X1 U3016 ( .A(n1209), .ZN(n4136) );
  AOI22_X1 U3017 ( .A1(n230), .A2(n168), .B1(n3592), .B2(\registers[24][29] ), 
        .ZN(n1209) );
  INV_X1 U3018 ( .A(n1210), .ZN(n4137) );
  AOI22_X1 U3019 ( .A1(n395), .A2(n603), .B1(n3593), .B2(\registers[24][30] ), 
        .ZN(n1210) );
  INV_X1 U3020 ( .A(n1225), .ZN(n4087) );
  AOI22_X1 U3021 ( .A1(n283), .A2(n684), .B1(n3584), .B2(\registers[23][10] ), 
        .ZN(n1225) );
  INV_X1 U3022 ( .A(n1226), .ZN(n4088) );
  AOI22_X1 U3023 ( .A1(n548), .A2(n766), .B1(n3583), .B2(\registers[23][11] ), 
        .ZN(n1226) );
  INV_X1 U3024 ( .A(n1227), .ZN(n4089) );
  AOI22_X1 U3025 ( .A1(n898), .A2(n206), .B1(n3586), .B2(\registers[23][12] ), 
        .ZN(n1227) );
  INV_X1 U3026 ( .A(n1228), .ZN(n4090) );
  AOI22_X1 U3027 ( .A1(n284), .A2(n3582), .B1(n3585), .B2(\registers[23][13] ), 
        .ZN(n1228) );
  INV_X1 U3028 ( .A(n1229), .ZN(n4091) );
  AOI22_X1 U3029 ( .A1(n223), .A2(n766), .B1(n3584), .B2(\registers[23][14] ), 
        .ZN(n1229) );
  INV_X1 U3030 ( .A(n1230), .ZN(n4092) );
  AOI22_X1 U3031 ( .A1(n209), .A2(n684), .B1(n3585), .B2(\registers[23][15] ), 
        .ZN(n1230) );
  INV_X1 U3032 ( .A(n1231), .ZN(n4093) );
  AOI22_X1 U3033 ( .A1(n262), .A2(n3580), .B1(n3583), .B2(\registers[23][16] ), 
        .ZN(n1231) );
  INV_X1 U3034 ( .A(n1232), .ZN(n4094) );
  AOI22_X1 U3035 ( .A1(n250), .A2(n765), .B1(n3584), .B2(\registers[23][17] ), 
        .ZN(n1232) );
  INV_X1 U3036 ( .A(n1233), .ZN(n4095) );
  AOI22_X1 U3037 ( .A1(n886), .A2(n3581), .B1(n3583), .B2(\registers[23][18] ), 
        .ZN(n1233) );
  INV_X1 U3038 ( .A(n1234), .ZN(n4096) );
  AOI22_X1 U3039 ( .A1(n416), .A2(n3581), .B1(n3586), .B2(\registers[23][19] ), 
        .ZN(n1234) );
  INV_X1 U3040 ( .A(n1235), .ZN(n4097) );
  AOI22_X1 U3041 ( .A1(n882), .A2(n3582), .B1(n3584), .B2(\registers[23][20] ), 
        .ZN(n1235) );
  INV_X1 U3042 ( .A(n1236), .ZN(n4098) );
  AOI22_X1 U3043 ( .A1(n880), .A2(n3582), .B1(n3586), .B2(\registers[23][21] ), 
        .ZN(n1236) );
  INV_X1 U3044 ( .A(n1237), .ZN(n4099) );
  AOI22_X1 U3045 ( .A1(n245), .A2(n684), .B1(n3585), .B2(\registers[23][22] ), 
        .ZN(n1237) );
  INV_X1 U3046 ( .A(n1238), .ZN(n4100) );
  AOI22_X1 U3047 ( .A1(n265), .A2(n684), .B1(n3583), .B2(\registers[23][23] ), 
        .ZN(n1238) );
  INV_X1 U3048 ( .A(n1239), .ZN(n4101) );
  AOI22_X1 U3049 ( .A1(n398), .A2(n3581), .B1(n3583), .B2(\registers[23][24] ), 
        .ZN(n1239) );
  INV_X1 U3050 ( .A(n1240), .ZN(n4102) );
  AOI22_X1 U3051 ( .A1(n200), .A2(n766), .B1(n3586), .B2(\registers[23][25] ), 
        .ZN(n1240) );
  INV_X1 U3052 ( .A(n1241), .ZN(n4103) );
  AOI22_X1 U3053 ( .A1(n870), .A2(n206), .B1(n3586), .B2(\registers[23][26] ), 
        .ZN(n1241) );
  INV_X1 U3054 ( .A(n1242), .ZN(n4104) );
  AOI22_X1 U3055 ( .A1(n868), .A2(n3580), .B1(n3584), .B2(\registers[23][27] ), 
        .ZN(n1242) );
  INV_X1 U3056 ( .A(n1243), .ZN(n4105) );
  AOI22_X1 U3057 ( .A1(net28529), .A2(n3580), .B1(n3585), .B2(
        \registers[23][28] ), .ZN(n1243) );
  INV_X1 U3058 ( .A(n1244), .ZN(n4106) );
  AOI22_X1 U3059 ( .A1(n866), .A2(n766), .B1(n3586), .B2(\registers[23][29] ), 
        .ZN(n1244) );
  INV_X1 U3060 ( .A(n1245), .ZN(n4107) );
  AOI22_X1 U3061 ( .A1(n394), .A2(n206), .B1(n3584), .B2(\registers[23][30] ), 
        .ZN(n1245) );
  INV_X1 U3062 ( .A(n1259), .ZN(n4060) );
  AOI22_X1 U3063 ( .A1(n283), .A2(net26245), .B1(n241), .B2(
        \registers[22][10] ), .ZN(n1259) );
  INV_X1 U3064 ( .A(n1260), .ZN(n4061) );
  AOI22_X1 U3065 ( .A1(n796), .A2(net26243), .B1(net44604), .B2(
        \registers[22][11] ), .ZN(n1260) );
  INV_X1 U3066 ( .A(n1262), .ZN(n4062) );
  AOI22_X1 U3067 ( .A1(n284), .A2(net26245), .B1(net26249), .B2(
        \registers[22][13] ), .ZN(n1262) );
  INV_X1 U3068 ( .A(n1263), .ZN(n4063) );
  AOI22_X1 U3069 ( .A1(n894), .A2(net26245), .B1(net44604), .B2(
        \registers[22][14] ), .ZN(n1263) );
  INV_X1 U3070 ( .A(n1264), .ZN(n4064) );
  AOI22_X1 U3071 ( .A1(n209), .A2(n25), .B1(net44604), .B2(\registers[22][15] ), .ZN(n1264) );
  INV_X1 U3072 ( .A(n1265), .ZN(n4065) );
  AOI22_X1 U3073 ( .A1(n262), .A2(n25), .B1(net44322), .B2(\registers[22][16] ), .ZN(n1265) );
  INV_X1 U3074 ( .A(n1266), .ZN(n4066) );
  AOI22_X1 U3075 ( .A1(n250), .A2(net26247), .B1(net38912), .B2(
        \registers[22][17] ), .ZN(n1266) );
  INV_X1 U3076 ( .A(n1267), .ZN(n4067) );
  AOI22_X1 U3077 ( .A1(n886), .A2(net26245), .B1(net44322), .B2(
        \registers[22][18] ), .ZN(n1267) );
  INV_X1 U3078 ( .A(n1268), .ZN(n4068) );
  AOI22_X1 U3079 ( .A1(n416), .A2(net44303), .B1(net26249), .B2(
        \registers[22][19] ), .ZN(n1268) );
  INV_X1 U3080 ( .A(n1270), .ZN(n4069) );
  AOI22_X1 U3081 ( .A1(n880), .A2(net44304), .B1(net44860), .B2(
        \registers[22][21] ), .ZN(n1270) );
  INV_X1 U3082 ( .A(n1272), .ZN(n4070) );
  AOI22_X1 U3083 ( .A1(n265), .A2(net26247), .B1(n20), .B2(\registers[22][23] ), .ZN(n1272) );
  INV_X1 U3084 ( .A(n1273), .ZN(n4071) );
  AOI22_X1 U3085 ( .A1(n409), .A2(net26243), .B1(n241), .B2(
        \registers[22][24] ), .ZN(n1273) );
  INV_X1 U3086 ( .A(n1274), .ZN(n4072) );
  AOI22_X1 U3087 ( .A1(n200), .A2(net44303), .B1(net38912), .B2(
        \registers[22][25] ), .ZN(n1274) );
  INV_X1 U3088 ( .A(n1275), .ZN(n4073) );
  AOI22_X1 U3089 ( .A1(n870), .A2(n25), .B1(net38912), .B2(\registers[22][26] ), .ZN(n1275) );
  INV_X1 U3090 ( .A(n1276), .ZN(n4074) );
  AOI22_X1 U3091 ( .A1(n557), .A2(net44303), .B1(net26249), .B2(
        \registers[22][27] ), .ZN(n1276) );
  INV_X1 U3092 ( .A(n1278), .ZN(n4075) );
  AOI22_X1 U3093 ( .A1(n866), .A2(net26243), .B1(net38912), .B2(
        \registers[22][29] ), .ZN(n1278) );
  INV_X1 U3094 ( .A(n1279), .ZN(n4076) );
  AOI22_X1 U3095 ( .A1(n394), .A2(net44304), .B1(n241), .B2(
        \registers[22][30] ), .ZN(n1279) );
  INV_X1 U3096 ( .A(n1294), .ZN(n4028) );
  AOI22_X1 U3097 ( .A1(n283), .A2(n3570), .B1(n3572), .B2(\registers[19][10] ), 
        .ZN(n1294) );
  INV_X1 U3098 ( .A(n1295), .ZN(n4029) );
  AOI22_X1 U3099 ( .A1(n796), .A2(n244), .B1(n3572), .B2(\registers[19][11] ), 
        .ZN(n1295) );
  INV_X1 U3100 ( .A(n1296), .ZN(n4030) );
  AOI22_X1 U3101 ( .A1(n898), .A2(n3570), .B1(n3572), .B2(\registers[19][12] ), 
        .ZN(n1296) );
  INV_X1 U3102 ( .A(n1297), .ZN(n4031) );
  AOI22_X1 U3103 ( .A1(n284), .A2(n243), .B1(n3572), .B2(\registers[19][13] ), 
        .ZN(n1297) );
  INV_X1 U3104 ( .A(n1298), .ZN(n4032) );
  AOI22_X1 U3105 ( .A1(n894), .A2(n760), .B1(n3573), .B2(\registers[19][14] ), 
        .ZN(n1298) );
  INV_X1 U3106 ( .A(n1299), .ZN(n4033) );
  AOI22_X1 U3107 ( .A1(n209), .A2(n244), .B1(n3571), .B2(\registers[19][15] ), 
        .ZN(n1299) );
  INV_X1 U3108 ( .A(n1300), .ZN(n4034) );
  AOI22_X1 U3109 ( .A1(n261), .A2(n3568), .B1(n3573), .B2(\registers[19][16] ), 
        .ZN(n1300) );
  INV_X1 U3110 ( .A(n1301), .ZN(n4035) );
  AOI22_X1 U3111 ( .A1(n888), .A2(n243), .B1(n3571), .B2(\registers[19][17] ), 
        .ZN(n1301) );
  INV_X1 U3112 ( .A(n1302), .ZN(n4036) );
  AOI22_X1 U3113 ( .A1(n259), .A2(n243), .B1(n3571), .B2(\registers[19][18] ), 
        .ZN(n1302) );
  INV_X1 U3114 ( .A(n1303), .ZN(n4037) );
  AOI22_X1 U3115 ( .A1(n416), .A2(n760), .B1(n3572), .B2(\registers[19][19] ), 
        .ZN(n1303) );
  INV_X1 U3116 ( .A(n1304), .ZN(n4038) );
  AOI22_X1 U3117 ( .A1(n207), .A2(n761), .B1(n3573), .B2(\registers[19][20] ), 
        .ZN(n1304) );
  INV_X1 U3118 ( .A(n1305), .ZN(n4039) );
  AOI22_X1 U3119 ( .A1(n880), .A2(n3569), .B1(n3), .B2(\registers[19][21] ), 
        .ZN(n1305) );
  INV_X1 U3120 ( .A(n1306), .ZN(n4040) );
  AOI22_X1 U3121 ( .A1(n245), .A2(n577), .B1(n3572), .B2(\registers[19][22] ), 
        .ZN(n1306) );
  INV_X1 U3122 ( .A(n1307), .ZN(n4041) );
  AOI22_X1 U3123 ( .A1(n264), .A2(n577), .B1(n3571), .B2(\registers[19][23] ), 
        .ZN(n1307) );
  INV_X1 U3124 ( .A(n1308), .ZN(n4042) );
  AOI22_X1 U3125 ( .A1(n398), .A2(n3569), .B1(n3572), .B2(\registers[19][24] ), 
        .ZN(n1308) );
  INV_X1 U3126 ( .A(n1309), .ZN(n4043) );
  AOI22_X1 U3127 ( .A1(n199), .A2(n761), .B1(n3572), .B2(\registers[19][25] ), 
        .ZN(n1309) );
  INV_X1 U3128 ( .A(n1310), .ZN(n4044) );
  AOI22_X1 U3129 ( .A1(n870), .A2(n243), .B1(n3571), .B2(\registers[19][26] ), 
        .ZN(n1310) );
  INV_X1 U3130 ( .A(n1311), .ZN(n4045) );
  AOI22_X1 U3131 ( .A1(n556), .A2(n244), .B1(n3571), .B2(\registers[19][27] ), 
        .ZN(n1311) );
  INV_X1 U3132 ( .A(n1312), .ZN(n4046) );
  AOI22_X1 U3133 ( .A1(n246), .A2(n243), .B1(n3573), .B2(\registers[19][28] ), 
        .ZN(n1312) );
  INV_X1 U3134 ( .A(n1313), .ZN(n4047) );
  AOI22_X1 U3135 ( .A1(n231), .A2(n3568), .B1(n31), .B2(\registers[19][29] ), 
        .ZN(n1313) );
  INV_X1 U3136 ( .A(n1314), .ZN(n4048) );
  AOI22_X1 U3137 ( .A1(n800), .A2(n3568), .B1(n3573), .B2(\registers[19][30] ), 
        .ZN(n1314) );
  INV_X1 U3138 ( .A(n1327), .ZN(n3996) );
  AOI22_X1 U3139 ( .A1(n799), .A2(n595), .B1(n3565), .B2(\registers[18][10] ), 
        .ZN(n1327) );
  INV_X1 U3140 ( .A(n1328), .ZN(n3997) );
  AOI22_X1 U3141 ( .A1(n549), .A2(n758), .B1(n3566), .B2(\registers[18][11] ), 
        .ZN(n1328) );
  INV_X1 U3142 ( .A(n1329), .ZN(n3998) );
  AOI22_X1 U3143 ( .A1(n166), .A2(n759), .B1(n3566), .B2(\registers[18][12] ), 
        .ZN(n1329) );
  INV_X1 U3144 ( .A(n1330), .ZN(n3999) );
  AOI22_X1 U3145 ( .A1(n896), .A2(n3562), .B1(n3565), .B2(\registers[18][13] ), 
        .ZN(n1330) );
  INV_X1 U3146 ( .A(n1331), .ZN(n4000) );
  AOI22_X1 U3147 ( .A1(n223), .A2(n3564), .B1(n3565), .B2(\registers[18][14] ), 
        .ZN(n1331) );
  INV_X1 U3148 ( .A(n1332), .ZN(n4001) );
  AOI22_X1 U3149 ( .A1(n210), .A2(n3563), .B1(n3565), .B2(\registers[18][15] ), 
        .ZN(n1332) );
  INV_X1 U3150 ( .A(n1333), .ZN(n4002) );
  AOI22_X1 U3151 ( .A1(n890), .A2(n3562), .B1(n3566), .B2(\registers[18][16] ), 
        .ZN(n1333) );
  INV_X1 U3152 ( .A(n1334), .ZN(n4003) );
  AOI22_X1 U3153 ( .A1(n888), .A2(n3562), .B1(n3565), .B2(\registers[18][17] ), 
        .ZN(n1334) );
  INV_X1 U3154 ( .A(n1335), .ZN(n4004) );
  AOI22_X1 U3155 ( .A1(n259), .A2(n758), .B1(n3565), .B2(\registers[18][18] ), 
        .ZN(n1335) );
  INV_X1 U3156 ( .A(n1336), .ZN(n4005) );
  AOI22_X1 U3157 ( .A1(n883), .A2(n3563), .B1(n3565), .B2(\registers[18][19] ), 
        .ZN(n1336) );
  INV_X1 U3158 ( .A(n1337), .ZN(n4006) );
  AOI22_X1 U3159 ( .A1(n207), .A2(n759), .B1(n3565), .B2(\registers[18][20] ), 
        .ZN(n1337) );
  INV_X1 U3160 ( .A(n1338), .ZN(n4007) );
  AOI22_X1 U3161 ( .A1(n242), .A2(n759), .B1(n3565), .B2(\registers[18][21] ), 
        .ZN(n1338) );
  INV_X1 U3162 ( .A(n1339), .ZN(n4008) );
  AOI22_X1 U3163 ( .A1(n877), .A2(n759), .B1(n3565), .B2(\registers[18][22] ), 
        .ZN(n1339) );
  INV_X1 U3164 ( .A(n1340), .ZN(n4009) );
  AOI22_X1 U3165 ( .A1(n876), .A2(n595), .B1(n3566), .B2(\registers[18][23] ), 
        .ZN(n1340) );
  INV_X1 U3166 ( .A(n1341), .ZN(n4010) );
  AOI22_X1 U3167 ( .A1(n397), .A2(n758), .B1(n3566), .B2(\registers[18][24] ), 
        .ZN(n1341) );
  INV_X1 U3168 ( .A(n1342), .ZN(n4011) );
  AOI22_X1 U3169 ( .A1(n199), .A2(n758), .B1(n3565), .B2(\registers[18][25] ), 
        .ZN(n1342) );
  INV_X1 U3170 ( .A(n1343), .ZN(n4012) );
  AOI22_X1 U3171 ( .A1(n558), .A2(n758), .B1(n3565), .B2(\registers[18][26] ), 
        .ZN(n1343) );
  INV_X1 U3172 ( .A(n1344), .ZN(n4013) );
  AOI22_X1 U3173 ( .A1(n556), .A2(n3564), .B1(n3565), .B2(\registers[18][27] ), 
        .ZN(n1344) );
  INV_X1 U3174 ( .A(n1345), .ZN(n4014) );
  AOI22_X1 U3175 ( .A1(n246), .A2(n758), .B1(n3566), .B2(\registers[18][28] ), 
        .ZN(n1345) );
  INV_X1 U3176 ( .A(n1346), .ZN(n4015) );
  AOI22_X1 U3177 ( .A1(n230), .A2(n3563), .B1(n3565), .B2(\registers[18][29] ), 
        .ZN(n1346) );
  INV_X1 U3178 ( .A(n1347), .ZN(n4016) );
  AOI22_X1 U3179 ( .A1(n395), .A2(n595), .B1(n3565), .B2(\registers[18][30] ), 
        .ZN(n1347) );
  INV_X1 U3180 ( .A(n1365), .ZN(n3869) );
  AOI22_X1 U3181 ( .A1(n799), .A2(n687), .B1(n217), .B2(\registers[13][10] ), 
        .ZN(n1365) );
  INV_X1 U3182 ( .A(n1366), .ZN(n3870) );
  AOI22_X1 U3183 ( .A1(n796), .A2(n3544), .B1(n217), .B2(\registers[13][11] ), 
        .ZN(n1366) );
  INV_X1 U3184 ( .A(n1367), .ZN(n3871) );
  AOI22_X1 U3185 ( .A1(n165), .A2(n3545), .B1(n218), .B2(\registers[13][12] ), 
        .ZN(n1367) );
  INV_X1 U3186 ( .A(n1368), .ZN(n3872) );
  AOI22_X1 U3187 ( .A1(n284), .A2(n3546), .B1(n218), .B2(\registers[13][13] ), 
        .ZN(n1368) );
  INV_X1 U3188 ( .A(n1369), .ZN(n3873) );
  AOI22_X1 U3189 ( .A1(n894), .A2(n3546), .B1(n217), .B2(\registers[13][14] ), 
        .ZN(n1369) );
  INV_X1 U3190 ( .A(n1371), .ZN(n3874) );
  AOI22_X1 U3191 ( .A1(n262), .A2(n775), .B1(n220), .B2(\registers[13][16] ), 
        .ZN(n1371) );
  INV_X1 U3192 ( .A(n1372), .ZN(n3875) );
  AOI22_X1 U3193 ( .A1(n888), .A2(n687), .B1(n216), .B2(\registers[13][17] ), 
        .ZN(n1372) );
  INV_X1 U3194 ( .A(n1373), .ZN(n3876) );
  AOI22_X1 U3195 ( .A1(n886), .A2(n408), .B1(n3550), .B2(\registers[13][18] ), 
        .ZN(n1373) );
  INV_X1 U3196 ( .A(n1374), .ZN(n3877) );
  AOI22_X1 U3197 ( .A1(n545), .A2(n3544), .B1(n220), .B2(\registers[13][19] ), 
        .ZN(n1374) );
  INV_X1 U3198 ( .A(n1375), .ZN(n3878) );
  AOI22_X1 U3199 ( .A1(n207), .A2(n687), .B1(n215), .B2(\registers[13][20] ), 
        .ZN(n1375) );
  INV_X1 U3200 ( .A(n1376), .ZN(n3879) );
  AOI22_X1 U3201 ( .A1(n242), .A2(n408), .B1(n17), .B2(\registers[13][21] ), 
        .ZN(n1376) );
  INV_X1 U3202 ( .A(n1377), .ZN(n3880) );
  AOI22_X1 U3203 ( .A1(n19), .A2(n775), .B1(n219), .B2(\registers[13][22] ), 
        .ZN(n1377) );
  INV_X1 U3204 ( .A(n1378), .ZN(n3881) );
  AOI22_X1 U3205 ( .A1(n265), .A2(n775), .B1(n3548), .B2(\registers[13][23] ), 
        .ZN(n1378) );
  INV_X1 U3206 ( .A(n1379), .ZN(n3882) );
  AOI22_X1 U3207 ( .A1(n411), .A2(n408), .B1(n218), .B2(\registers[13][24] ), 
        .ZN(n1379) );
  INV_X1 U3208 ( .A(n1380), .ZN(n3883) );
  AOI22_X1 U3209 ( .A1(n200), .A2(n3545), .B1(n3550), .B2(\registers[13][25] ), 
        .ZN(n1380) );
  INV_X1 U3210 ( .A(n1381), .ZN(n3884) );
  AOI22_X1 U3211 ( .A1(n559), .A2(n687), .B1(n3549), .B2(\registers[13][26] ), 
        .ZN(n1381) );
  INV_X1 U3212 ( .A(n1382), .ZN(n3885) );
  AOI22_X1 U3213 ( .A1(n868), .A2(n3544), .B1(n3549), .B2(\registers[13][27] ), 
        .ZN(n1382) );
  INV_X1 U3214 ( .A(n1383), .ZN(n3886) );
  AOI22_X1 U3215 ( .A1(net28529), .A2(n3546), .B1(n218), .B2(
        \registers[13][28] ), .ZN(n1383) );
  INV_X1 U3216 ( .A(n1384), .ZN(n3887) );
  AOI22_X1 U3217 ( .A1(n866), .A2(n3545), .B1(n3548), .B2(\registers[13][29] ), 
        .ZN(n1384) );
  INV_X1 U3218 ( .A(n1385), .ZN(n3888) );
  AOI22_X1 U3219 ( .A1(n394), .A2(n408), .B1(n218), .B2(\registers[13][30] ), 
        .ZN(n1385) );
  INV_X1 U3220 ( .A(n1398), .ZN(n3838) );
  AOI22_X1 U3221 ( .A1(n283), .A2(n693), .B1(n3541), .B2(\registers[12][10] ), 
        .ZN(n1398) );
  INV_X1 U3222 ( .A(n1399), .ZN(n3839) );
  AOI22_X1 U3223 ( .A1(n796), .A2(n3538), .B1(n3539), .B2(\registers[12][11] ), 
        .ZN(n1399) );
  INV_X1 U3224 ( .A(n1401), .ZN(n3840) );
  AOI22_X1 U3225 ( .A1(n284), .A2(n693), .B1(n3540), .B2(\registers[12][13] ), 
        .ZN(n1401) );
  INV_X1 U3226 ( .A(n1402), .ZN(n3841) );
  AOI22_X1 U3227 ( .A1(n894), .A2(n693), .B1(n3541), .B2(\registers[12][14] ), 
        .ZN(n1402) );
  INV_X1 U3228 ( .A(n1403), .ZN(n3842) );
  AOI22_X1 U3229 ( .A1(n210), .A2(n3537), .B1(n3542), .B2(\registers[12][15] ), 
        .ZN(n1403) );
  INV_X1 U3230 ( .A(n1404), .ZN(n3843) );
  AOI22_X1 U3231 ( .A1(n261), .A2(n3537), .B1(n3540), .B2(\registers[12][16] ), 
        .ZN(n1404) );
  INV_X1 U3232 ( .A(n1405), .ZN(n3844) );
  AOI22_X1 U3233 ( .A1(n250), .A2(n769), .B1(n3542), .B2(\registers[12][17] ), 
        .ZN(n1405) );
  INV_X1 U3234 ( .A(n1406), .ZN(n3845) );
  AOI22_X1 U3235 ( .A1(n259), .A2(n692), .B1(n3540), .B2(\registers[12][18] ), 
        .ZN(n1406) );
  INV_X1 U3236 ( .A(n1407), .ZN(n3846) );
  AOI22_X1 U3237 ( .A1(n545), .A2(n770), .B1(n3542), .B2(\registers[12][19] ), 
        .ZN(n1407) );
  INV_X1 U3238 ( .A(n1408), .ZN(n3847) );
  AOI22_X1 U3239 ( .A1(n882), .A2(n203), .B1(n3540), .B2(\registers[12][20] ), 
        .ZN(n1408) );
  INV_X1 U3240 ( .A(n1409), .ZN(n3848) );
  AOI22_X1 U3241 ( .A1(n242), .A2(n3538), .B1(n3540), .B2(\registers[12][21] ), 
        .ZN(n1409) );
  INV_X1 U3242 ( .A(n1410), .ZN(n3849) );
  AOI22_X1 U3243 ( .A1(n19), .A2(n770), .B1(n3542), .B2(\registers[12][22] ), 
        .ZN(n1410) );
  INV_X1 U3244 ( .A(n1411), .ZN(n3850) );
  AOI22_X1 U3245 ( .A1(n264), .A2(n3537), .B1(n3542), .B2(\registers[12][23] ), 
        .ZN(n1411) );
  INV_X1 U3246 ( .A(n1412), .ZN(n3851) );
  AOI22_X1 U3247 ( .A1(n411), .A2(n3538), .B1(n3539), .B2(\registers[12][24] ), 
        .ZN(n1412) );
  INV_X1 U3248 ( .A(n1413), .ZN(n3852) );
  AOI22_X1 U3249 ( .A1(n199), .A2(n692), .B1(n3541), .B2(\registers[12][25] ), 
        .ZN(n1413) );
  INV_X1 U3250 ( .A(n1414), .ZN(n3853) );
  AOI22_X1 U3251 ( .A1(n559), .A2(n204), .B1(n3539), .B2(\registers[12][26] ), 
        .ZN(n1414) );
  INV_X1 U3252 ( .A(n1415), .ZN(n3854) );
  AOI22_X1 U3253 ( .A1(n556), .A2(n769), .B1(n3540), .B2(\registers[12][27] ), 
        .ZN(n1415) );
  INV_X1 U3254 ( .A(n1416), .ZN(n3855) );
  AOI22_X1 U3255 ( .A1(n246), .A2(n769), .B1(n3541), .B2(\registers[12][28] ), 
        .ZN(n1416) );
  INV_X1 U3256 ( .A(n1417), .ZN(n3856) );
  AOI22_X1 U3257 ( .A1(n231), .A2(n203), .B1(n3539), .B2(\registers[12][29] ), 
        .ZN(n1417) );
  INV_X1 U3258 ( .A(n1418), .ZN(n3857) );
  AOI22_X1 U3259 ( .A1(n800), .A2(n769), .B1(n3541), .B2(\registers[12][30] ), 
        .ZN(n1418) );
  INV_X1 U3260 ( .A(n1433), .ZN(n3807) );
  AOI22_X1 U3261 ( .A1(n799), .A2(n679), .B1(n3521), .B2(\registers[9][10] ), 
        .ZN(n1433) );
  INV_X1 U3262 ( .A(n1434), .ZN(n3808) );
  AOI22_X1 U3263 ( .A1(n548), .A2(n774), .B1(n3525), .B2(\registers[9][11] ), 
        .ZN(n1434) );
  INV_X1 U3264 ( .A(n1435), .ZN(n3809) );
  AOI22_X1 U3265 ( .A1(n898), .A2(n3519), .B1(n3522), .B2(\registers[9][12] ), 
        .ZN(n1435) );
  INV_X1 U3266 ( .A(n1436), .ZN(n3810) );
  AOI22_X1 U3267 ( .A1(n284), .A2(n774), .B1(n3526), .B2(\registers[9][13] ), 
        .ZN(n1436) );
  INV_X1 U3268 ( .A(n1438), .ZN(n3811) );
  AOI22_X1 U3269 ( .A1(n892), .A2(n3518), .B1(n3522), .B2(\registers[9][15] ), 
        .ZN(n1438) );
  INV_X1 U3270 ( .A(n1439), .ZN(n3812) );
  AOI22_X1 U3271 ( .A1(n890), .A2(n3519), .B1(n3523), .B2(\registers[9][16] ), 
        .ZN(n1439) );
  INV_X1 U3272 ( .A(n1440), .ZN(n3813) );
  AOI22_X1 U3273 ( .A1(n887), .A2(n3520), .B1(n3525), .B2(\registers[9][17] ), 
        .ZN(n1440) );
  INV_X1 U3274 ( .A(n1441), .ZN(n3814) );
  AOI22_X1 U3275 ( .A1(n886), .A2(n3520), .B1(n3522), .B2(\registers[9][18] ), 
        .ZN(n1441) );
  INV_X1 U3276 ( .A(n1442), .ZN(n3815) );
  AOI22_X1 U3277 ( .A1(n545), .A2(n3518), .B1(n3523), .B2(\registers[9][19] ), 
        .ZN(n1442) );
  INV_X1 U3278 ( .A(n1443), .ZN(n3816) );
  AOI22_X1 U3279 ( .A1(n207), .A2(n3520), .B1(n3526), .B2(\registers[9][20] ), 
        .ZN(n1443) );
  INV_X1 U3280 ( .A(n1444), .ZN(n3817) );
  AOI22_X1 U3281 ( .A1(n242), .A2(n3519), .B1(n3524), .B2(\registers[9][21] ), 
        .ZN(n1444) );
  INV_X1 U3282 ( .A(n1445), .ZN(n3818) );
  AOI22_X1 U3283 ( .A1(n245), .A2(n774), .B1(n3521), .B2(\registers[9][22] ), 
        .ZN(n1445) );
  INV_X1 U3284 ( .A(n1446), .ZN(n3819) );
  AOI22_X1 U3285 ( .A1(n876), .A2(n773), .B1(n3525), .B2(\registers[9][23] ), 
        .ZN(n1446) );
  INV_X1 U3286 ( .A(n1447), .ZN(n3820) );
  AOI22_X1 U3287 ( .A1(n409), .A2(n680), .B1(n3522), .B2(\registers[9][24] ), 
        .ZN(n1447) );
  INV_X1 U3288 ( .A(n1448), .ZN(n3821) );
  AOI22_X1 U3289 ( .A1(n872), .A2(n773), .B1(n3521), .B2(\registers[9][25] ), 
        .ZN(n1448) );
  INV_X1 U3290 ( .A(n1449), .ZN(n3822) );
  AOI22_X1 U3291 ( .A1(n559), .A2(n680), .B1(n3524), .B2(\registers[9][26] ), 
        .ZN(n1449) );
  INV_X1 U3292 ( .A(n1450), .ZN(n3823) );
  AOI22_X1 U3293 ( .A1(n868), .A2(n3518), .B1(n3524), .B2(\registers[9][27] ), 
        .ZN(n1450) );
  INV_X1 U3294 ( .A(n1451), .ZN(n3824) );
  AOI22_X1 U3295 ( .A1(n246), .A2(n679), .B1(n3526), .B2(\registers[9][28] ), 
        .ZN(n1451) );
  INV_X1 U3296 ( .A(n1452), .ZN(n3825) );
  AOI22_X1 U3297 ( .A1(n231), .A2(n680), .B1(n3523), .B2(\registers[9][29] ), 
        .ZN(n1452) );
  INV_X1 U3298 ( .A(n1453), .ZN(n3826) );
  AOI22_X1 U3299 ( .A1(n395), .A2(n773), .B1(n3527), .B2(\registers[9][30] ), 
        .ZN(n1453) );
  INV_X1 U3300 ( .A(n1466), .ZN(n3776) );
  AOI22_X1 U3301 ( .A1(n799), .A2(n389), .B1(n3515), .B2(\registers[8][10] ), 
        .ZN(n1466) );
  INV_X1 U3302 ( .A(n1467), .ZN(n3777) );
  AOI22_X1 U3303 ( .A1(n548), .A2(n276), .B1(n3514), .B2(\registers[8][11] ), 
        .ZN(n1467) );
  INV_X1 U3304 ( .A(n1468), .ZN(n3778) );
  AOI22_X1 U3305 ( .A1(n898), .A2(n3512), .B1(n3516), .B2(\registers[8][12] ), 
        .ZN(n1468) );
  INV_X1 U3306 ( .A(n1469), .ZN(n3779) );
  AOI22_X1 U3307 ( .A1(n896), .A2(n3513), .B1(n3516), .B2(\registers[8][13] ), 
        .ZN(n1469) );
  INV_X1 U3308 ( .A(n1470), .ZN(n3780) );
  AOI22_X1 U3309 ( .A1(n894), .A2(n3512), .B1(n3515), .B2(\registers[8][14] ), 
        .ZN(n1470) );
  INV_X1 U3310 ( .A(n1471), .ZN(n3781) );
  AOI22_X1 U3311 ( .A1(n209), .A2(n276), .B1(n3516), .B2(\registers[8][15] ), 
        .ZN(n1471) );
  INV_X1 U3312 ( .A(n1472), .ZN(n3782) );
  AOI22_X1 U3313 ( .A1(n262), .A2(n277), .B1(n3515), .B2(\registers[8][16] ), 
        .ZN(n1472) );
  INV_X1 U3314 ( .A(n1473), .ZN(n3783) );
  AOI22_X1 U3315 ( .A1(n888), .A2(n277), .B1(n3515), .B2(\registers[8][17] ), 
        .ZN(n1473) );
  INV_X1 U3316 ( .A(n1475), .ZN(n3784) );
  AOI22_X1 U3317 ( .A1(n545), .A2(n276), .B1(n3516), .B2(\registers[8][19] ), 
        .ZN(n1475) );
  INV_X1 U3318 ( .A(n1476), .ZN(n3785) );
  AOI22_X1 U3319 ( .A1(n882), .A2(n389), .B1(n3514), .B2(\registers[8][20] ), 
        .ZN(n1476) );
  INV_X1 U3320 ( .A(n1477), .ZN(n3786) );
  AOI22_X1 U3321 ( .A1(n880), .A2(n277), .B1(n3516), .B2(\registers[8][21] ), 
        .ZN(n1477) );
  INV_X1 U3322 ( .A(n1478), .ZN(n3787) );
  AOI22_X1 U3323 ( .A1(n19), .A2(n3512), .B1(n3516), .B2(\registers[8][22] ), 
        .ZN(n1478) );
  INV_X1 U3324 ( .A(n1479), .ZN(n3788) );
  AOI22_X1 U3325 ( .A1(n876), .A2(n390), .B1(n3515), .B2(\registers[8][23] ), 
        .ZN(n1479) );
  INV_X1 U3326 ( .A(n1480), .ZN(n3789) );
  AOI22_X1 U3327 ( .A1(n409), .A2(n276), .B1(n3514), .B2(\registers[8][24] ), 
        .ZN(n1480) );
  INV_X1 U3328 ( .A(n1481), .ZN(n3790) );
  AOI22_X1 U3329 ( .A1(n872), .A2(n276), .B1(n3514), .B2(\registers[8][25] ), 
        .ZN(n1481) );
  INV_X1 U3330 ( .A(n1482), .ZN(n3791) );
  AOI22_X1 U3331 ( .A1(n558), .A2(n276), .B1(n3516), .B2(\registers[8][26] ), 
        .ZN(n1482) );
  INV_X1 U3332 ( .A(n1483), .ZN(n3792) );
  AOI22_X1 U3333 ( .A1(n557), .A2(n3513), .B1(n3515), .B2(\registers[8][27] ), 
        .ZN(n1483) );
  INV_X1 U3334 ( .A(n1484), .ZN(n3793) );
  AOI22_X1 U3335 ( .A1(net28529), .A2(n277), .B1(n3516), .B2(
        \registers[8][28] ), .ZN(n1484) );
  INV_X1 U3336 ( .A(n1485), .ZN(n3794) );
  AOI22_X1 U3337 ( .A1(n230), .A2(n3513), .B1(n3516), .B2(\registers[8][29] ), 
        .ZN(n1485) );
  INV_X1 U3338 ( .A(n1486), .ZN(n3795) );
  AOI22_X1 U3339 ( .A1(n394), .A2(n390), .B1(n3516), .B2(\registers[8][30] ), 
        .ZN(n1486) );
  INV_X1 U3340 ( .A(n1499), .ZN(n3963) );
  AOI22_X1 U3341 ( .A1(n799), .A2(n3505), .B1(n3509), .B2(\registers[7][10] ), 
        .ZN(n1499) );
  INV_X1 U3342 ( .A(n1500), .ZN(n3964) );
  AOI22_X1 U3343 ( .A1(n549), .A2(n764), .B1(n3510), .B2(\registers[7][11] ), 
        .ZN(n1500) );
  INV_X1 U3344 ( .A(n1501), .ZN(n3965) );
  AOI22_X1 U3345 ( .A1(n166), .A2(n214), .B1(n3507), .B2(\registers[7][12] ), 
        .ZN(n1501) );
  INV_X1 U3346 ( .A(n1502), .ZN(n3966) );
  AOI22_X1 U3347 ( .A1(n896), .A2(n682), .B1(n3510), .B2(\registers[7][13] ), 
        .ZN(n1502) );
  INV_X1 U3348 ( .A(n1503), .ZN(n3967) );
  AOI22_X1 U3349 ( .A1(n223), .A2(n3506), .B1(n3510), .B2(\registers[7][14] ), 
        .ZN(n1503) );
  INV_X1 U3350 ( .A(n1504), .ZN(n3968) );
  AOI22_X1 U3351 ( .A1(n892), .A2(n683), .B1(n3508), .B2(\registers[7][15] ), 
        .ZN(n1504) );
  INV_X1 U3352 ( .A(n1505), .ZN(n3969) );
  AOI22_X1 U3353 ( .A1(n261), .A2(n213), .B1(n3509), .B2(\registers[7][16] ), 
        .ZN(n1505) );
  INV_X1 U3354 ( .A(n1506), .ZN(n3970) );
  AOI22_X1 U3355 ( .A1(n250), .A2(n3506), .B1(n3510), .B2(\registers[7][17] ), 
        .ZN(n1506) );
  INV_X1 U3356 ( .A(n1507), .ZN(n3971) );
  AOI22_X1 U3357 ( .A1(n259), .A2(n213), .B1(n3509), .B2(\registers[7][18] ), 
        .ZN(n1507) );
  INV_X1 U3358 ( .A(n1508), .ZN(n3972) );
  AOI22_X1 U3359 ( .A1(n883), .A2(n214), .B1(n3508), .B2(\registers[7][19] ), 
        .ZN(n1508) );
  INV_X1 U3360 ( .A(n1509), .ZN(n3973) );
  AOI22_X1 U3361 ( .A1(n207), .A2(n3505), .B1(n3509), .B2(\registers[7][20] ), 
        .ZN(n1509) );
  INV_X1 U3362 ( .A(n1510), .ZN(n3974) );
  AOI22_X1 U3363 ( .A1(n880), .A2(n3505), .B1(n3508), .B2(\registers[7][21] ), 
        .ZN(n1510) );
  INV_X1 U3364 ( .A(n1511), .ZN(n3975) );
  AOI22_X1 U3365 ( .A1(n245), .A2(n764), .B1(n3510), .B2(\registers[7][22] ), 
        .ZN(n1511) );
  INV_X1 U3366 ( .A(n1512), .ZN(n3976) );
  AOI22_X1 U3367 ( .A1(n264), .A2(n682), .B1(n3507), .B2(\registers[7][23] ), 
        .ZN(n1512) );
  INV_X1 U3368 ( .A(n1513), .ZN(n3977) );
  AOI22_X1 U3369 ( .A1(n410), .A2(n764), .B1(n3508), .B2(\registers[7][24] ), 
        .ZN(n1513) );
  INV_X1 U3370 ( .A(n1514), .ZN(n3978) );
  AOI22_X1 U3371 ( .A1(n200), .A2(n682), .B1(n3507), .B2(\registers[7][25] ), 
        .ZN(n1514) );
  INV_X1 U3372 ( .A(n1515), .ZN(n3979) );
  AOI22_X1 U3373 ( .A1(n870), .A2(n683), .B1(n3507), .B2(\registers[7][26] ), 
        .ZN(n1515) );
  INV_X1 U3374 ( .A(n1516), .ZN(n3980) );
  AOI22_X1 U3375 ( .A1(n557), .A2(n3506), .B1(n3507), .B2(\registers[7][27] ), 
        .ZN(n1516) );
  INV_X1 U3376 ( .A(n1517), .ZN(n3981) );
  AOI22_X1 U3377 ( .A1(net28529), .A2(n213), .B1(n3509), .B2(
        \registers[7][28] ), .ZN(n1517) );
  INV_X1 U3378 ( .A(n1518), .ZN(n3982) );
  AOI22_X1 U3379 ( .A1(n866), .A2(n213), .B1(n3508), .B2(\registers[7][29] ), 
        .ZN(n1518) );
  INV_X1 U3380 ( .A(n1519), .ZN(n3983) );
  AOI22_X1 U3381 ( .A1(n395), .A2(n682), .B1(n3509), .B2(\registers[7][30] ), 
        .ZN(n1519) );
  INV_X1 U3382 ( .A(n1533), .ZN(n3932) );
  AOI22_X1 U3383 ( .A1(n283), .A2(n229), .B1(net26585), .B2(\registers[6][10] ), .ZN(n1533) );
  INV_X1 U3384 ( .A(n1534), .ZN(n3933) );
  AOI22_X1 U3385 ( .A1(n548), .A2(net39089), .B1(net26595), .B2(
        \registers[6][11] ), .ZN(n1534) );
  INV_X1 U3386 ( .A(n1535), .ZN(n3934) );
  AOI22_X1 U3387 ( .A1(n165), .A2(net38992), .B1(net26595), .B2(
        \registers[6][12] ), .ZN(n1535) );
  INV_X1 U3388 ( .A(n1536), .ZN(n3935) );
  AOI22_X1 U3389 ( .A1(n896), .A2(net26581), .B1(net26597), .B2(
        \registers[6][13] ), .ZN(n1536) );
  INV_X1 U3390 ( .A(n1537), .ZN(n3936) );
  AOI22_X1 U3391 ( .A1(n228), .A2(n223), .B1(net26595), .B2(\registers[6][14] ), .ZN(n1537) );
  INV_X1 U3392 ( .A(n1539), .ZN(n3937) );
  AOI22_X1 U3393 ( .A1(n261), .A2(net39090), .B1(net26597), .B2(
        \registers[6][16] ), .ZN(n1539) );
  INV_X1 U3394 ( .A(n1540), .ZN(n3938) );
  AOI22_X1 U3395 ( .A1(n888), .A2(net38993), .B1(net26589), .B2(
        \registers[6][17] ), .ZN(n1540) );
  INV_X1 U3396 ( .A(n1541), .ZN(n3939) );
  AOI22_X1 U3397 ( .A1(n259), .A2(net26579), .B1(net26585), .B2(
        \registers[6][18] ), .ZN(n1541) );
  INV_X1 U3398 ( .A(n1542), .ZN(n3940) );
  AOI22_X1 U3399 ( .A1(n545), .A2(net39089), .B1(net26589), .B2(
        \registers[6][19] ), .ZN(n1542) );
  INV_X1 U3400 ( .A(n1543), .ZN(n3941) );
  AOI22_X1 U3401 ( .A1(n882), .A2(n32), .B1(net26589), .B2(\registers[6][20] ), 
        .ZN(n1543) );
  INV_X1 U3402 ( .A(n1544), .ZN(n3942) );
  AOI22_X1 U3403 ( .A1(n880), .A2(net26583), .B1(net26585), .B2(
        \registers[6][21] ), .ZN(n1544) );
  INV_X1 U3404 ( .A(n1545), .ZN(n3943) );
  AOI22_X1 U3405 ( .A1(n245), .A2(n229), .B1(net26597), .B2(\registers[6][22] ), .ZN(n1545) );
  INV_X1 U3406 ( .A(n1546), .ZN(n3944) );
  AOI22_X1 U3407 ( .A1(n876), .A2(net39090), .B1(net26591), .B2(
        \registers[6][23] ), .ZN(n1546) );
  INV_X1 U3408 ( .A(n1547), .ZN(n3945) );
  AOI22_X1 U3409 ( .A1(n397), .A2(net26581), .B1(net26595), .B2(
        \registers[6][24] ), .ZN(n1547) );
  INV_X1 U3410 ( .A(n1548), .ZN(n3946) );
  AOI22_X1 U3411 ( .A1(n872), .A2(net26579), .B1(net26589), .B2(
        \registers[6][25] ), .ZN(n1548) );
  INV_X1 U3412 ( .A(n1549), .ZN(n3947) );
  AOI22_X1 U3413 ( .A1(n559), .A2(net38992), .B1(net26585), .B2(
        \registers[6][26] ), .ZN(n1549) );
  INV_X1 U3414 ( .A(n1550), .ZN(n3948) );
  AOI22_X1 U3415 ( .A1(n556), .A2(n228), .B1(net26591), .B2(\registers[6][27] ), .ZN(n1550) );
  INV_X1 U3416 ( .A(n1551), .ZN(n3949) );
  AOI22_X1 U3417 ( .A1(net28529), .A2(net38992), .B1(net26591), .B2(
        \registers[6][28] ), .ZN(n1551) );
  INV_X1 U3418 ( .A(n1552), .ZN(n3950) );
  AOI22_X1 U3419 ( .A1(n230), .A2(n32), .B1(net26595), .B2(\registers[6][29] ), 
        .ZN(n1552) );
  INV_X1 U3420 ( .A(n1553), .ZN(n3951) );
  AOI22_X1 U3421 ( .A1(n800), .A2(n32), .B1(net26585), .B2(\registers[6][30] ), 
        .ZN(n1553) );
  INV_X1 U3422 ( .A(n1570), .ZN(n3900) );
  AOI22_X1 U3423 ( .A1(n799), .A2(n3494), .B1(n3497), .B2(\registers[1][10] ), 
        .ZN(n1570) );
  INV_X1 U3424 ( .A(n1571), .ZN(n3901) );
  AOI22_X1 U3425 ( .A1(n796), .A2(n678), .B1(n3498), .B2(\registers[1][11] ), 
        .ZN(n1571) );
  INV_X1 U3426 ( .A(n1572), .ZN(n3902) );
  AOI22_X1 U3427 ( .A1(n898), .A2(n677), .B1(n3499), .B2(\registers[1][12] ), 
        .ZN(n1572) );
  INV_X1 U3428 ( .A(n1573), .ZN(n3903) );
  AOI22_X1 U3429 ( .A1(n896), .A2(n3494), .B1(n3499), .B2(\registers[1][13] ), 
        .ZN(n1573) );
  INV_X1 U3430 ( .A(n1574), .ZN(n3904) );
  AOI22_X1 U3431 ( .A1(n223), .A2(n771), .B1(n3498), .B2(\registers[1][14] ), 
        .ZN(n1574) );
  INV_X1 U3432 ( .A(n1575), .ZN(n3905) );
  AOI22_X1 U3433 ( .A1(n210), .A2(n3492), .B1(n3498), .B2(\registers[1][15] ), 
        .ZN(n1575) );
  INV_X1 U3434 ( .A(n1576), .ZN(n3906) );
  AOI22_X1 U3435 ( .A1(n890), .A2(n3493), .B1(n3496), .B2(\registers[1][16] ), 
        .ZN(n1576) );
  INV_X1 U3436 ( .A(n1577), .ZN(n3907) );
  AOI22_X1 U3437 ( .A1(n888), .A2(n3493), .B1(n3499), .B2(\registers[1][17] ), 
        .ZN(n1577) );
  INV_X1 U3438 ( .A(n1578), .ZN(n3908) );
  AOI22_X1 U3439 ( .A1(n886), .A2(n678), .B1(n3499), .B2(\registers[1][18] ), 
        .ZN(n1578) );
  INV_X1 U3440 ( .A(n1579), .ZN(n3909) );
  AOI22_X1 U3441 ( .A1(n883), .A2(n3492), .B1(n3498), .B2(\registers[1][19] ), 
        .ZN(n1579) );
  INV_X1 U3442 ( .A(n1580), .ZN(n3910) );
  AOI22_X1 U3443 ( .A1(n161), .A2(n772), .B1(n3495), .B2(\registers[1][20] ), 
        .ZN(n1580) );
  INV_X1 U3444 ( .A(n1581), .ZN(n3911) );
  AOI22_X1 U3445 ( .A1(n242), .A2(n772), .B1(n3495), .B2(\registers[1][21] ), 
        .ZN(n1581) );
  INV_X1 U3446 ( .A(n1582), .ZN(n3912) );
  AOI22_X1 U3447 ( .A1(n877), .A2(n772), .B1(n3497), .B2(\registers[1][22] ), 
        .ZN(n1582) );
  INV_X1 U3448 ( .A(n1583), .ZN(n3913) );
  AOI22_X1 U3449 ( .A1(n265), .A2(n772), .B1(n3496), .B2(\registers[1][23] ), 
        .ZN(n1583) );
  INV_X1 U3450 ( .A(n1584), .ZN(n3914) );
  AOI22_X1 U3451 ( .A1(n411), .A2(n678), .B1(n3499), .B2(\registers[1][24] ), 
        .ZN(n1584) );
  INV_X1 U3452 ( .A(n1585), .ZN(n3915) );
  AOI22_X1 U3453 ( .A1(n199), .A2(n771), .B1(n3496), .B2(\registers[1][25] ), 
        .ZN(n1585) );
  INV_X1 U3454 ( .A(n1586), .ZN(n3916) );
  AOI22_X1 U3455 ( .A1(n870), .A2(n771), .B1(n3500), .B2(\registers[1][26] ), 
        .ZN(n1586) );
  INV_X1 U3456 ( .A(n1587), .ZN(n3917) );
  AOI22_X1 U3457 ( .A1(n556), .A2(n3492), .B1(n3501), .B2(\registers[1][27] ), 
        .ZN(n1587) );
  INV_X1 U3458 ( .A(n1588), .ZN(n3918) );
  AOI22_X1 U3459 ( .A1(n246), .A2(n771), .B1(n3497), .B2(\registers[1][28] ), 
        .ZN(n1588) );
  INV_X1 U3460 ( .A(n1589), .ZN(n3919) );
  AOI22_X1 U3461 ( .A1(n231), .A2(n678), .B1(n3495), .B2(\registers[1][29] ), 
        .ZN(n1589) );
  INV_X1 U3462 ( .A(n1590), .ZN(n3920) );
  AOI22_X1 U3463 ( .A1(n394), .A2(n677), .B1(n3501), .B2(\registers[1][30] ), 
        .ZN(n1590) );
  INV_X1 U3464 ( .A(n1348), .ZN(n4017) );
  AOI22_X1 U3465 ( .A1(n785), .A2(n759), .B1(n3565), .B2(\registers[18][31] ), 
        .ZN(n1348) );
  INV_X1 U3466 ( .A(n1315), .ZN(n4049) );
  AOI22_X1 U3467 ( .A1(n785), .A2(n760), .B1(n3), .B2(\registers[19][31] ), 
        .ZN(n1315) );
  INV_X1 U3468 ( .A(n1177), .ZN(n4170) );
  AOI22_X1 U3469 ( .A1(n550), .A2(n778), .B1(n597), .B2(\registers[25][31] ), 
        .ZN(n1177) );
  INV_X1 U3470 ( .A(n1386), .ZN(n3889) );
  AOI22_X1 U3471 ( .A1(n785), .A2(n3544), .B1(n215), .B2(\registers[13][31] ), 
        .ZN(n1386) );
  INV_X1 U3472 ( .A(n1419), .ZN(n3858) );
  AOI22_X1 U3473 ( .A1(n550), .A2(n3538), .B1(n3540), .B2(\registers[12][31] ), 
        .ZN(n1419) );
  INV_X1 U3474 ( .A(n1105), .ZN(n4232) );
  AOI22_X1 U3475 ( .A1(n550), .A2(n3634), .B1(n3637), .B2(\registers[29][31] ), 
        .ZN(n1105) );
  INV_X1 U3476 ( .A(n1139), .ZN(n4201) );
  AOI22_X1 U3477 ( .A1(n550), .A2(n767), .B1(n3631), .B2(\registers[28][31] ), 
        .ZN(n1139) );
  INV_X1 U3478 ( .A(n1246), .ZN(n4108) );
  AOI22_X1 U3479 ( .A1(n550), .A2(n3580), .B1(n3586), .B2(\registers[23][31] ), 
        .ZN(n1246) );
  INV_X1 U3480 ( .A(n1520), .ZN(n3984) );
  AOI22_X1 U3481 ( .A1(n785), .A2(n683), .B1(n3510), .B2(\registers[7][31] ), 
        .ZN(n1520) );
  INV_X1 U3482 ( .A(n1454), .ZN(n3827) );
  AOI22_X1 U3483 ( .A1(n550), .A2(n773), .B1(n3527), .B2(\registers[9][31] ), 
        .ZN(n1454) );
  INV_X1 U3484 ( .A(n1591), .ZN(n3921) );
  AOI22_X1 U3485 ( .A1(n785), .A2(n772), .B1(n3501), .B2(\registers[1][31] ), 
        .ZN(n1591) );
  INV_X1 U3486 ( .A(n1280), .ZN(n4077) );
  AOI22_X1 U3487 ( .A1(n550), .A2(net44304), .B1(net44605), .B2(
        \registers[22][31] ), .ZN(n1280) );
  INV_X1 U3488 ( .A(n1554), .ZN(n3952) );
  AOI22_X1 U3489 ( .A1(n550), .A2(net38993), .B1(net26595), .B2(
        \registers[6][31] ), .ZN(n1554) );
  INV_X1 U3490 ( .A(n1487), .ZN(n3796) );
  AOI22_X1 U3491 ( .A1(n785), .A2(n389), .B1(n3516), .B2(\registers[8][31] ), 
        .ZN(n1487) );
  INV_X1 U3492 ( .A(n1211), .ZN(n4138) );
  AOI22_X1 U3493 ( .A1(n785), .A2(n171), .B1(n3592), .B2(\registers[24][31] ), 
        .ZN(n1211) );
  AND2_X1 U3494 ( .A1(RD2), .A2(ENABLE), .ZN(N218) );
  AND2_X1 U3495 ( .A1(RD1), .A2(ENABLE), .ZN(N83) );
  INV_X1 U3496 ( .A(n1003), .ZN(n905) );
  INV_X1 U3497 ( .A(n926), .ZN(n906) );
  INV_X1 U3498 ( .A(n1000), .ZN(n907) );
  INV_X1 U3499 ( .A(n1002), .ZN(n908) );
  INV_X1 U3500 ( .A(n1001), .ZN(n909) );
  INV_X1 U3501 ( .A(n999), .ZN(n910) );
  INV_X1 U3502 ( .A(n997), .ZN(n911) );
  INV_X1 U3503 ( .A(n993), .ZN(n912) );
  INV_X1 U3504 ( .A(n925), .ZN(n913) );
  INV_X1 U3505 ( .A(n927), .ZN(n914) );
  INV_X1 U3506 ( .A(n998), .ZN(n915) );
  INV_X1 U3507 ( .A(n924), .ZN(n916) );
  INV_X1 U3508 ( .A(n995), .ZN(n917) );
  INV_X1 U3509 ( .A(n926), .ZN(n918) );
  INV_X1 U3510 ( .A(n996), .ZN(n919) );
  INV_X1 U3511 ( .A(n928), .ZN(n920) );
  INV_X1 U3512 ( .A(n1350), .ZN(n921) );
  INV_X1 U3513 ( .A(n1350), .ZN(n922) );
  INV_X1 U3514 ( .A(n1350), .ZN(n923) );
  INV_X1 U3515 ( .A(n921), .ZN(n924) );
  INV_X1 U3516 ( .A(n921), .ZN(n925) );
  INV_X1 U3517 ( .A(n923), .ZN(n926) );
  INV_X1 U3518 ( .A(n922), .ZN(n927) );
  INV_X1 U3519 ( .A(n923), .ZN(n928) );
  INV_X1 U3520 ( .A(n921), .ZN(n993) );
  INV_X1 U3521 ( .A(n3556), .ZN(n994) );
  INV_X1 U3522 ( .A(n923), .ZN(n995) );
  INV_X1 U3523 ( .A(n922), .ZN(n996) );
  INV_X1 U3524 ( .A(n3556), .ZN(n997) );
  INV_X1 U3525 ( .A(n922), .ZN(n998) );
  INV_X1 U3526 ( .A(n922), .ZN(n999) );
  INV_X1 U3527 ( .A(n921), .ZN(n1000) );
  INV_X1 U3528 ( .A(n921), .ZN(n1001) );
  INV_X1 U3529 ( .A(n922), .ZN(n1002) );
  INV_X1 U3530 ( .A(n3556), .ZN(n1003) );
  INV_X1 U3531 ( .A(n3559), .ZN(n1004) );
  INV_X1 U3532 ( .A(n1004), .ZN(n1005) );
  INV_X1 U3533 ( .A(n1004), .ZN(n1006) );
  INV_X1 U3534 ( .A(n1004), .ZN(n1007) );
  INV_X1 U3535 ( .A(n3557), .ZN(n1008) );
  INV_X1 U3536 ( .A(n1008), .ZN(n1009) );
  INV_X1 U3537 ( .A(n1008), .ZN(n1010) );
  INV_X1 U3538 ( .A(n1008), .ZN(n1011) );
  INV_X1 U3539 ( .A(n3558), .ZN(n1012) );
  INV_X1 U3540 ( .A(n1012), .ZN(n1013) );
  INV_X1 U3541 ( .A(n1012), .ZN(n1014) );
  INV_X1 U3542 ( .A(n3559), .ZN(n1015) );
  INV_X1 U3543 ( .A(n1015), .ZN(n1016) );
  INV_X1 U3544 ( .A(n1026), .ZN(n1017) );
  INV_X1 U3545 ( .A(n1027), .ZN(n1018) );
  INV_X1 U3546 ( .A(n1012), .ZN(n1019) );
  INV_X1 U3547 ( .A(n1028), .ZN(n1020) );
  INV_X1 U3548 ( .A(n3558), .ZN(n1021) );
  INV_X1 U3549 ( .A(n3561), .ZN(n1022) );
  INV_X1 U3550 ( .A(n3557), .ZN(n1023) );
  INV_X1 U3551 ( .A(n3560), .ZN(n1024) );
  INV_X1 U3552 ( .A(n3561), .ZN(n1025) );
  INV_X1 U3553 ( .A(n3560), .ZN(n1026) );
  INV_X1 U3554 ( .A(n3560), .ZN(n1027) );
  INV_X1 U3555 ( .A(n3561), .ZN(n1028) );
  CLKBUF_X1 U3556 ( .A(n187), .Z(n3557) );
  CLKBUF_X1 U3557 ( .A(n187), .Z(n3558) );
  INV_X1 U3558 ( .A(n1047), .ZN(n1029) );
  INV_X1 U3559 ( .A(n3555), .ZN(n1030) );
  INV_X1 U3560 ( .A(n1046), .ZN(n1031) );
  INV_X1 U3561 ( .A(n3554), .ZN(n1032) );
  INV_X1 U3562 ( .A(n3554), .ZN(n1033) );
  INV_X1 U3563 ( .A(n3553), .ZN(n1034) );
  INV_X1 U3564 ( .A(n3553), .ZN(n1035) );
  INV_X1 U3565 ( .A(n3553), .ZN(n1036) );
  INV_X1 U3566 ( .A(n3552), .ZN(n1037) );
  INV_X1 U3567 ( .A(n3552), .ZN(n1038) );
  INV_X1 U3568 ( .A(n3551), .ZN(n1039) );
  INV_X1 U3569 ( .A(n3552), .ZN(n1040) );
  INV_X1 U3570 ( .A(n3554), .ZN(n1041) );
  INV_X1 U3571 ( .A(n3551), .ZN(n1042) );
  INV_X1 U3572 ( .A(n3551), .ZN(n1043) );
  INV_X1 U3573 ( .A(n266), .ZN(n1044) );
  INV_X1 U3574 ( .A(n266), .ZN(n1045) );
  INV_X1 U3575 ( .A(n1351), .ZN(n1046) );
  INV_X1 U3576 ( .A(n266), .ZN(n1047) );
  BUF_X1 U3577 ( .A(n3555), .Z(n3553) );
  OAI22_X1 U3578 ( .A1(n554), .A2(n1021), .B1(n1009), .B2(n539), .ZN(n2971) );
  OAI22_X1 U3579 ( .A1(n193), .A2(n1028), .B1(n1020), .B2(n540), .ZN(n2970) );
  OAI22_X1 U3580 ( .A1(n400), .A2(n1027), .B1(n1019), .B2(n541), .ZN(n2969) );
  OAI22_X1 U3581 ( .A1(n194), .A2(n1027), .B1(n1018), .B2(n542), .ZN(n2968) );
  OAI22_X1 U3582 ( .A1(n191), .A2(n1026), .B1(n1019), .B2(n543), .ZN(n2967) );
  OAI22_X1 U3583 ( .A1(n607), .A2(n1022), .B1(n1018), .B2(n544), .ZN(n2966) );
  OAI22_X1 U3584 ( .A1(n9), .A2(n1025), .B1(n1014), .B2(n537), .ZN(n2973) );
  OAI22_X1 U3585 ( .A1(n546), .A2(n1024), .B1(n1013), .B2(n538), .ZN(n2972) );
  OAI22_X1 U3586 ( .A1(n23), .A2(net38966), .B1(n12), .B2(n934), .ZN(n2832) );
  OAI22_X1 U3587 ( .A1(n29), .A2(net38964), .B1(net38969), .B2(n933), .ZN(
        n2833) );
  OAI22_X1 U3588 ( .A1(net17879), .A2(net38964), .B1(net38974), .B2(n932), 
        .ZN(n2834) );
  OAI22_X1 U3589 ( .A1(n271), .A2(net38965), .B1(net38974), .B2(n931), .ZN(
        n2835) );
  OAI22_X1 U3590 ( .A1(n221), .A2(net38964), .B1(net38968), .B2(n930), .ZN(
        n2836) );
  OAI22_X1 U3591 ( .A1(n605), .A2(net38965), .B1(net38970), .B2(n929), .ZN(
        n2837) );
  INV_X1 U3592 ( .A(n590), .ZN(n1048) );
  INV_X1 U3593 ( .A(n1048), .ZN(n1049) );
  INV_X1 U3594 ( .A(n1048), .ZN(n1050) );
  INV_X1 U3595 ( .A(n1048), .ZN(n1051) );
  INV_X1 U3596 ( .A(n1269), .ZN(n1052) );
  INV_X1 U3597 ( .A(n1201), .ZN(n1053) );
  INV_X1 U3598 ( .A(n1271), .ZN(n1054) );
  INV_X1 U3599 ( .A(n1204), .ZN(n1055) );
  INV_X1 U3600 ( .A(n3529), .ZN(n1056) );
  INV_X1 U3601 ( .A(n1056), .ZN(n1057) );
  INV_X1 U3602 ( .A(n3529), .ZN(n1058) );
  INV_X1 U3603 ( .A(n1058), .ZN(n1059) );
  INV_X1 U3604 ( .A(n1058), .ZN(n1060) );
  INV_X1 U3605 ( .A(n1058), .ZN(n1061) );
  INV_X1 U3606 ( .A(n1218), .ZN(n1062) );
  INV_X1 U3607 ( .A(n1370), .ZN(n1063) );
  INV_X1 U3608 ( .A(n3531), .ZN(n1064) );
  INV_X1 U3609 ( .A(n1064), .ZN(n1065) );
  INV_X1 U3610 ( .A(n1064), .ZN(n1066) );
  INV_X1 U3611 ( .A(n1064), .ZN(n1067) );
  INV_X1 U3612 ( .A(n3532), .ZN(n1071) );
  INV_X1 U3613 ( .A(n1071), .ZN(n1098) );
  INV_X1 U3614 ( .A(n1071), .ZN(n1115) );
  INV_X1 U3615 ( .A(n1071), .ZN(n1141) );
  INV_X1 U3616 ( .A(n3532), .ZN(n1143) );
  INV_X1 U3617 ( .A(n3533), .ZN(n1201) );
  INV_X1 U3618 ( .A(n3528), .ZN(n1204) );
  INV_X1 U3619 ( .A(n3530), .ZN(n1218) );
  INV_X1 U3620 ( .A(n3531), .ZN(n1261) );
  INV_X1 U3621 ( .A(n3533), .ZN(n1269) );
  INV_X1 U3622 ( .A(n3528), .ZN(n1271) );
  INV_X1 U3623 ( .A(n3531), .ZN(n1281) );
  INV_X1 U3624 ( .A(n3529), .ZN(n1349) );
  INV_X1 U3625 ( .A(n1051), .ZN(n1353) );
  INV_X1 U3626 ( .A(n3530), .ZN(n1370) );
  INV_X1 U3627 ( .A(n1049), .ZN(n1400) );
  BUF_X1 U3628 ( .A(n590), .Z(n3533) );
  BUF_X1 U3629 ( .A(n590), .Z(n3528) );
  CLKBUF_X1 U3630 ( .A(n590), .Z(n3530) );
  CLKBUF_X1 U3631 ( .A(n590), .Z(n3532) );
  INV_X1 U3632 ( .A(n3305), .ZN(n1421) );
  INV_X1 U3633 ( .A(n3315), .ZN(n1437) );
  INV_X1 U3634 ( .A(n3307), .ZN(n1474) );
  INV_X1 U3635 ( .A(n3307), .ZN(n1538) );
  INV_X1 U3636 ( .A(n3305), .ZN(n3286) );
  INV_X1 U3637 ( .A(n3315), .ZN(n3287) );
  INV_X1 U3638 ( .A(n3314), .ZN(n3288) );
  INV_X1 U3639 ( .A(n3307), .ZN(n3289) );
  INV_X1 U3640 ( .A(n3313), .ZN(n3290) );
  INV_X1 U3641 ( .A(n3304), .ZN(n3291) );
  INV_X1 U3642 ( .A(n3311), .ZN(n3292) );
  INV_X1 U3643 ( .A(n3304), .ZN(n3293) );
  INV_X1 U3644 ( .A(n3312), .ZN(n3294) );
  INV_X1 U3645 ( .A(n3305), .ZN(n3295) );
  INV_X1 U3646 ( .A(n3314), .ZN(n3296) );
  INV_X1 U3647 ( .A(n3311), .ZN(n3297) );
  INV_X1 U3648 ( .A(n3312), .ZN(n3298) );
  INV_X1 U3649 ( .A(n3310), .ZN(n3299) );
  INV_X1 U3650 ( .A(n1420), .ZN(n3300) );
  INV_X1 U3651 ( .A(n1420), .ZN(n3301) );
  INV_X1 U3652 ( .A(n3536), .ZN(n3302) );
  INV_X1 U3653 ( .A(n3534), .ZN(n3303) );
  INV_X1 U3654 ( .A(n3301), .ZN(n3304) );
  INV_X1 U3655 ( .A(n3300), .ZN(n3305) );
  INV_X1 U3656 ( .A(n3536), .ZN(n3306) );
  INV_X1 U3657 ( .A(n3300), .ZN(n3307) );
  INV_X1 U3658 ( .A(n3535), .ZN(n3308) );
  INV_X1 U3659 ( .A(n3536), .ZN(n3309) );
  INV_X1 U3660 ( .A(n3536), .ZN(n3310) );
  INV_X1 U3661 ( .A(n3301), .ZN(n3311) );
  INV_X1 U3662 ( .A(n3301), .ZN(n3312) );
  INV_X1 U3663 ( .A(n3536), .ZN(n3313) );
  INV_X1 U3664 ( .A(n3301), .ZN(n3314) );
  INV_X1 U3665 ( .A(n3300), .ZN(n3315) );
  INV_X1 U3666 ( .A(n3300), .ZN(n3316) );
  INV_X1 U3667 ( .A(n1420), .ZN(n3536) );
  BUF_X1 U3668 ( .A(n3536), .Z(n3535) );
  NAND2_X1 U3669 ( .A1(n1521), .A2(n414), .ZN(n1556) );
  OAI22_X1 U3670 ( .A1(n182), .A2(n751), .B1(n3502), .B2(n106), .ZN(n3212) );
  OAI22_X1 U3671 ( .A1(n4250), .A2(n750), .B1(n8), .B2(n105), .ZN(n3213) );
  OAI22_X1 U3672 ( .A1(n744), .A2(n750), .B1(n3502), .B2(n104), .ZN(n3214) );
  OAI22_X1 U3673 ( .A1(n4248), .A2(n749), .B1(n746), .B2(n103), .ZN(n3215) );
  OAI22_X1 U3674 ( .A1(n703), .A2(n750), .B1(n746), .B2(n117), .ZN(n3201) );
  OAI22_X1 U3675 ( .A1(n4261), .A2(n750), .B1(n3503), .B2(n118), .ZN(n3200) );
  OAI22_X1 U3676 ( .A1(n600), .A2(n749), .B1(n3502), .B2(n119), .ZN(n3199) );
  OAI22_X1 U3677 ( .A1(n4263), .A2(n749), .B1(n3504), .B2(n120), .ZN(n3198) );
  OAI22_X1 U3678 ( .A1(n260), .A2(n751), .B1(n3503), .B2(n109), .ZN(n3209) );
  OAI22_X1 U3679 ( .A1(n602), .A2(n750), .B1(n8), .B2(n110), .ZN(n3208) );
  OAI22_X1 U3680 ( .A1(n402), .A2(n751), .B1(n3502), .B2(n111), .ZN(n3207) );
  OAI22_X1 U3681 ( .A1(n553), .A2(n749), .B1(n748), .B2(n112), .ZN(n3206) );
  OAI22_X1 U3682 ( .A1(n281), .A2(n751), .B1(n8), .B2(n113), .ZN(n3205) );
  OAI22_X1 U3683 ( .A1(n4257), .A2(n750), .B1(n8), .B2(n114), .ZN(n3204) );
  OAI22_X1 U3684 ( .A1(n598), .A2(n750), .B1(n8), .B2(n115), .ZN(n3203) );
  OAI22_X1 U3685 ( .A1(n274), .A2(n749), .B1(n3502), .B2(n116), .ZN(n3202) );
  NAND2_X1 U3686 ( .A1(n1106), .A2(n1521), .ZN(n1555) );
  OAI22_X1 U3687 ( .A1(n730), .A2(n288), .B1(n369), .B2(n152), .ZN(n3166) );
  OAI22_X1 U3688 ( .A1(n600), .A2(n353), .B1(n366), .B2(n151), .ZN(n3167) );
  OAI22_X1 U3689 ( .A1(n178), .A2(n288), .B1(n359), .B2(n150), .ZN(n3168) );
  OAI22_X1 U3690 ( .A1(n703), .A2(n353), .B1(n359), .B2(n149), .ZN(n3169) );
  OAI22_X1 U3691 ( .A1(n555), .A2(net38964), .B1(net38974), .B2(n955), .ZN(
        n2811) );
  OAI22_X1 U3692 ( .A1(n275), .A2(net38966), .B1(net38970), .B2(n956), .ZN(
        n2810) );
  OAI22_X1 U3693 ( .A1(n239), .A2(net38966), .B1(net38972), .B2(n957), .ZN(
        n2809) );
  OAI22_X1 U3694 ( .A1(n170), .A2(net38964), .B1(n12), .B2(n958), .ZN(n2808)
         );
  OAI22_X1 U3695 ( .A1(n673), .A2(net38964), .B1(n12), .B2(n959), .ZN(n2807)
         );
  OAI22_X1 U3696 ( .A1(n198), .A2(net38964), .B1(n2), .B2(n960), .ZN(n2806) );
  OAI22_X1 U3697 ( .A1(n705), .A2(net38966), .B1(net38973), .B2(n953), .ZN(
        n2813) );
  OAI22_X1 U3698 ( .A1(n4265), .A2(net38965), .B1(net38968), .B2(n954), .ZN(
        n2812) );
  OAI22_X1 U3699 ( .A1(n607), .A2(net26415), .B1(net26419), .B2(n448), .ZN(
        n3062) );
  OAI22_X1 U3700 ( .A1(n608), .A2(net44473), .B1(net26419), .B2(n447), .ZN(
        n3063) );
  OAI22_X1 U3701 ( .A1(n4269), .A2(net44474), .B1(net26419), .B2(n446), .ZN(
        n3064) );
  OAI22_X1 U3702 ( .A1(n4268), .A2(net44473), .B1(net26419), .B2(n445), .ZN(
        n3065) );
  OAI22_X1 U3703 ( .A1(n4267), .A2(net26413), .B1(net26419), .B2(n444), .ZN(
        n3066) );
  OAI22_X1 U3704 ( .A1(n27), .A2(net26415), .B1(net26421), .B2(n443), .ZN(
        n3067) );
  NAND2_X1 U3705 ( .A1(n1247), .A2(n1144), .ZN(n1317) );
  OAI22_X1 U3706 ( .A1(n263), .A2(n3605), .B1(n3611), .B2(n801), .ZN(n2901) );
  OAI22_X1 U3707 ( .A1(net44818), .A2(n3605), .B1(n3613), .B2(n804), .ZN(n2898) );
  OAI22_X1 U3708 ( .A1(n706), .A2(n3605), .B1(n3613), .B2(n807), .ZN(n2895) );
  OAI22_X1 U3709 ( .A1(n10), .A2(n3605), .B1(n3612), .B2(n810), .ZN(n2892) );
  OAI22_X1 U3710 ( .A1(n708), .A2(n3605), .B1(n3612), .B2(n811), .ZN(n2891) );
  OAI22_X1 U3711 ( .A1(n6), .A2(n3605), .B1(n3612), .B2(n812), .ZN(n2890) );
  OAI22_X1 U3712 ( .A1(n399), .A2(n3605), .B1(n3608), .B2(n802), .ZN(n2900) );
  OAI22_X1 U3713 ( .A1(n742), .A2(n3605), .B1(n3613), .B2(n803), .ZN(n2899) );
  OAI22_X1 U3714 ( .A1(n4246), .A2(n3605), .B1(n3613), .B2(n805), .ZN(n2897)
         );
  OAI22_X1 U3715 ( .A1(n4247), .A2(n3605), .B1(n3613), .B2(n806), .ZN(n2896)
         );
  OAI22_X1 U3716 ( .A1(n4249), .A2(n3605), .B1(n3612), .B2(n808), .ZN(n2894)
         );
  OAI22_X1 U3717 ( .A1(n4250), .A2(n3605), .B1(n3612), .B2(n809), .ZN(n2893)
         );
  CLKBUF_X1 U3718 ( .A(n783), .Z(n3612) );
  CLKBUF_X1 U3719 ( .A(n783), .Z(n3613) );
  AND2_X1 U3720 ( .A1(n1142), .A2(n1070), .ZN(n3317) );
  OAI22_X1 U3721 ( .A1(n4253), .A2(n1026), .B1(n1014), .B2(n525), .ZN(n2985)
         );
  OAI22_X1 U3722 ( .A1(n602), .A2(n1025), .B1(n1013), .B2(n526), .ZN(n2984) );
  OAI22_X1 U3723 ( .A1(n403), .A2(n1025), .B1(n1006), .B2(n527), .ZN(n2983) );
  OAI22_X1 U3724 ( .A1(n553), .A2(n1021), .B1(n1005), .B2(n528), .ZN(n2982) );
  OAI22_X1 U3725 ( .A1(n180), .A2(n1028), .B1(n1020), .B2(n529), .ZN(n2981) );
  OAI22_X1 U3726 ( .A1(n269), .A2(n1022), .B1(n1011), .B2(n530), .ZN(n2980) );
  OAI22_X1 U3727 ( .A1(n598), .A2(n1025), .B1(n1010), .B2(n531), .ZN(n2979) );
  OAI22_X1 U3728 ( .A1(n15), .A2(n1024), .B1(n1009), .B2(n532), .ZN(n2978) );
  OAI22_X1 U3729 ( .A1(n574), .A2(n1023), .B1(n1007), .B2(n533), .ZN(n2977) );
  OAI22_X1 U3730 ( .A1(n4261), .A2(n1024), .B1(n1006), .B2(n534), .ZN(n2976)
         );
  OAI22_X1 U3731 ( .A1(n601), .A2(n1023), .B1(n1011), .B2(n535), .ZN(n2975) );
  OAI22_X1 U3732 ( .A1(n201), .A2(n1022), .B1(n1010), .B2(n536), .ZN(n2974) );
  NAND2_X1 U3733 ( .A1(n1178), .A2(n1352), .ZN(n1423) );
  NAND2_X1 U3734 ( .A1(n1178), .A2(n1521), .ZN(n1560) );
  NAND2_X1 U3735 ( .A1(n1178), .A2(n1070), .ZN(n1146) );
  OAI22_X1 U3736 ( .A1(n186), .A2(n1029), .B1(n192), .B2(n459), .ZN(n3051) );
  OAI22_X1 U3737 ( .A1(n4252), .A2(n1032), .B1(n233), .B2(n460), .ZN(n3050) );
  OAI22_X1 U3738 ( .A1(n172), .A2(n1031), .B1(n1044), .B2(n449), .ZN(n3061) );
  OAI22_X1 U3739 ( .A1(n270), .A2(n1043), .B1(n232), .B2(n450), .ZN(n3060) );
  OAI22_X1 U3740 ( .A1(n4245), .A2(n1030), .B1(n1044), .B2(n451), .ZN(n3059)
         );
  OAI22_X1 U3741 ( .A1(n197), .A2(n1031), .B1(n232), .B2(n452), .ZN(n3058) );
  OAI22_X1 U3742 ( .A1(n593), .A2(n1042), .B1(n233), .B2(n453), .ZN(n3057) );
  OAI22_X1 U3743 ( .A1(n1042), .A2(n591), .B1(n1045), .B2(n454), .ZN(n3056) );
  OAI22_X1 U3744 ( .A1(n707), .A2(n1029), .B1(n232), .B2(n455), .ZN(n3055) );
  OAI22_X1 U3745 ( .A1(n4249), .A2(n1043), .B1(n232), .B2(n456), .ZN(n3054) );
  OAI22_X1 U3746 ( .A1(n4250), .A2(n1030), .B1(n1045), .B2(n457), .ZN(n3053)
         );
  OAI22_X1 U3747 ( .A1(n700), .A2(n1030), .B1(n1046), .B2(n458), .ZN(n3052) );
  NAND2_X1 U3748 ( .A1(n676), .A2(n1070), .ZN(n1068) );
  NAND2_X1 U3749 ( .A1(n1247), .A2(n676), .ZN(n1215) );
  NAND2_X1 U3750 ( .A1(n1521), .A2(n1069), .ZN(n1489) );
  OAI22_X1 U3751 ( .A1(n185), .A2(n757), .B1(n3578), .B2(n619), .ZN(n2955) );
  NAND2_X1 U3752 ( .A1(n1247), .A2(n1140), .ZN(n1282) );
  OAI22_X1 U3753 ( .A1(n396), .A2(n370), .B1(n374), .B2(n652), .ZN(n2922) );
  OAI22_X1 U3754 ( .A1(n560), .A2(net38965), .B1(net38972), .B2(n941), .ZN(
        n2825) );
  OAI22_X1 U3755 ( .A1(n415), .A2(net38966), .B1(net38970), .B2(n942), .ZN(
        n2824) );
  OAI22_X1 U3756 ( .A1(n402), .A2(net38964), .B1(net38972), .B2(n943), .ZN(
        n2823) );
  OAI22_X1 U3757 ( .A1(n552), .A2(net38966), .B1(n12), .B2(n944), .ZN(n2822)
         );
  OAI22_X1 U3758 ( .A1(n728), .A2(net38964), .B1(n2), .B2(n945), .ZN(n2821) );
  OAI22_X1 U3759 ( .A1(n269), .A2(net38965), .B1(net38974), .B2(n946), .ZN(
        n2820) );
  OAI22_X1 U3760 ( .A1(n177), .A2(net38964), .B1(net38973), .B2(n947), .ZN(
        n2819) );
  OAI22_X1 U3761 ( .A1(n740), .A2(net38965), .B1(net38972), .B2(n948), .ZN(
        n2818) );
  OAI22_X1 U3762 ( .A1(n604), .A2(net38965), .B1(net38969), .B2(n949), .ZN(
        n2817) );
  OAI22_X1 U3763 ( .A1(n675), .A2(net38966), .B1(net38972), .B2(n950), .ZN(
        n2816) );
  OAI22_X1 U3764 ( .A1(n179), .A2(net38965), .B1(n2), .B2(n951), .ZN(n2815) );
  OAI22_X1 U3765 ( .A1(n201), .A2(net38965), .B1(net38969), .B2(n952), .ZN(
        n2814) );
  INV_X1 U3766 ( .A(n3501), .ZN(n3494) );
  INV_X1 U3767 ( .A(net26591), .ZN(net26583) );
  INV_X1 U3768 ( .A(n3527), .ZN(n3520) );
  INV_X1 U3769 ( .A(n3543), .ZN(n3538) );
  INV_X1 U3770 ( .A(n3548), .ZN(n3546) );
  INV_X1 U3771 ( .A(net33812), .ZN(net26417) );
  INV_X1 U3772 ( .A(n3567), .ZN(n3564) );
  INV_X1 U3773 ( .A(n3575), .ZN(n3570) );
  INV_X1 U3774 ( .A(n3587), .ZN(n3582) );
  INV_X1 U3775 ( .A(n3594), .ZN(n3590) );
  INV_X1 U3776 ( .A(n597), .ZN(n3597) );
  INV_X1 U3777 ( .A(n783), .ZN(n3607) );
  INV_X1 U3778 ( .A(n3622), .ZN(n3616) );
  INV_X1 U3779 ( .A(n3631), .ZN(n3625) );
  INV_X1 U3780 ( .A(n3639), .ZN(n3634) );
  CLKBUF_X1 U3781 ( .A(N218), .Z(n3640) );
  CLKBUF_X1 U3782 ( .A(N218), .Z(n3641) );
  CLKBUF_X1 U3783 ( .A(N218), .Z(n3642) );
  CLKBUF_X1 U3784 ( .A(N218), .Z(n3643) );
  CLKBUF_X1 U3785 ( .A(N83), .Z(n3644) );
  CLKBUF_X1 U3786 ( .A(N83), .Z(n3645) );
  CLKBUF_X1 U3787 ( .A(N83), .Z(n3646) );
  CLKBUF_X1 U3788 ( .A(N83), .Z(n3647) );
  CLKBUF_X1 U3789 ( .A(n3765), .Z(n3659) );
  CLKBUF_X1 U3790 ( .A(n3764), .Z(n3660) );
  CLKBUF_X1 U3791 ( .A(n3764), .Z(n3661) );
  CLKBUF_X1 U3792 ( .A(n3764), .Z(n3662) );
  CLKBUF_X1 U3793 ( .A(n3764), .Z(n3663) );
  CLKBUF_X1 U3794 ( .A(n3764), .Z(n3664) );
  CLKBUF_X1 U3795 ( .A(n3764), .Z(n3665) );
  CLKBUF_X1 U3796 ( .A(n3763), .Z(n3666) );
  CLKBUF_X1 U3797 ( .A(n3763), .Z(n3667) );
  CLKBUF_X1 U3798 ( .A(n3763), .Z(n3668) );
  CLKBUF_X1 U3799 ( .A(n3763), .Z(n3669) );
  CLKBUF_X1 U3800 ( .A(n3763), .Z(n3670) );
  CLKBUF_X1 U3801 ( .A(n3763), .Z(n3671) );
  CLKBUF_X1 U3802 ( .A(n3762), .Z(n3672) );
  CLKBUF_X1 U3803 ( .A(n3762), .Z(n3673) );
  CLKBUF_X1 U3804 ( .A(n3762), .Z(n3674) );
  CLKBUF_X1 U3805 ( .A(n3762), .Z(n3675) );
  CLKBUF_X1 U3806 ( .A(n3762), .Z(n3676) );
  CLKBUF_X1 U3807 ( .A(n3762), .Z(n3677) );
  CLKBUF_X1 U3808 ( .A(n3761), .Z(n3678) );
  CLKBUF_X1 U3809 ( .A(n3761), .Z(n3679) );
  CLKBUF_X1 U3810 ( .A(n3761), .Z(n3680) );
  CLKBUF_X1 U3811 ( .A(n3761), .Z(n3681) );
  CLKBUF_X1 U3812 ( .A(n3761), .Z(n3682) );
  CLKBUF_X1 U3813 ( .A(n3761), .Z(n3683) );
  CLKBUF_X1 U3814 ( .A(n3760), .Z(n3684) );
  CLKBUF_X1 U3815 ( .A(n3760), .Z(n3685) );
  CLKBUF_X1 U3816 ( .A(n3760), .Z(n3686) );
  CLKBUF_X1 U3817 ( .A(n3760), .Z(n3687) );
  CLKBUF_X1 U3818 ( .A(n3760), .Z(n3688) );
  CLKBUF_X1 U3819 ( .A(n3760), .Z(n3689) );
  CLKBUF_X1 U3820 ( .A(n3759), .Z(n3690) );
  CLKBUF_X1 U3821 ( .A(n3759), .Z(n3691) );
  CLKBUF_X1 U3822 ( .A(n3759), .Z(n3692) );
  CLKBUF_X1 U3823 ( .A(n3759), .Z(n3693) );
  CLKBUF_X1 U3824 ( .A(n3759), .Z(n3694) );
  CLKBUF_X1 U3825 ( .A(n3759), .Z(n3695) );
  CLKBUF_X1 U3826 ( .A(n3758), .Z(n3696) );
  CLKBUF_X1 U3827 ( .A(n3758), .Z(n3697) );
  CLKBUF_X1 U3828 ( .A(n3758), .Z(n3698) );
  CLKBUF_X1 U3829 ( .A(n3758), .Z(n3699) );
  CLKBUF_X1 U3830 ( .A(n3758), .Z(n3700) );
  CLKBUF_X1 U3831 ( .A(n3758), .Z(n3701) );
  CLKBUF_X1 U3832 ( .A(n3757), .Z(n3702) );
  CLKBUF_X1 U3833 ( .A(n3757), .Z(n3703) );
  CLKBUF_X1 U3834 ( .A(n3757), .Z(n3704) );
  CLKBUF_X1 U3835 ( .A(n3757), .Z(n3705) );
  CLKBUF_X1 U3836 ( .A(n3757), .Z(n3706) );
  CLKBUF_X1 U3837 ( .A(n3757), .Z(n3707) );
  CLKBUF_X1 U3838 ( .A(n3756), .Z(n3708) );
  CLKBUF_X1 U3839 ( .A(n3756), .Z(n3709) );
  CLKBUF_X1 U3840 ( .A(n3756), .Z(n3710) );
  CLKBUF_X1 U3841 ( .A(n3756), .Z(n3711) );
  CLKBUF_X1 U3842 ( .A(n3756), .Z(n3712) );
  CLKBUF_X1 U3843 ( .A(n3756), .Z(n3713) );
  CLKBUF_X1 U3844 ( .A(n3755), .Z(n3714) );
  CLKBUF_X1 U3845 ( .A(n3755), .Z(n3715) );
  CLKBUF_X1 U3846 ( .A(n3755), .Z(n3716) );
  CLKBUF_X1 U3847 ( .A(n3755), .Z(n3717) );
  CLKBUF_X1 U3848 ( .A(n3755), .Z(n3718) );
  CLKBUF_X1 U3849 ( .A(n3755), .Z(n3719) );
  CLKBUF_X1 U3850 ( .A(n3754), .Z(n3720) );
  CLKBUF_X1 U3851 ( .A(n3754), .Z(n3721) );
  CLKBUF_X1 U3852 ( .A(n3754), .Z(n3722) );
  CLKBUF_X1 U3853 ( .A(n3754), .Z(n3723) );
  CLKBUF_X1 U3854 ( .A(n3754), .Z(n3724) );
  CLKBUF_X1 U3855 ( .A(n3754), .Z(n3725) );
  CLKBUF_X1 U3856 ( .A(n3753), .Z(n3726) );
  CLKBUF_X1 U3857 ( .A(n3753), .Z(n3727) );
  CLKBUF_X1 U3858 ( .A(n3753), .Z(n3728) );
  CLKBUF_X1 U3859 ( .A(n3753), .Z(n3729) );
  CLKBUF_X1 U3860 ( .A(n3753), .Z(n3730) );
  CLKBUF_X1 U3861 ( .A(n3753), .Z(n3731) );
  CLKBUF_X1 U3862 ( .A(n3752), .Z(n3732) );
  CLKBUF_X1 U3863 ( .A(n3752), .Z(n3733) );
  CLKBUF_X1 U3864 ( .A(n3752), .Z(n3734) );
  CLKBUF_X1 U3865 ( .A(n3752), .Z(n3735) );
  CLKBUF_X1 U3866 ( .A(n3752), .Z(n3736) );
  CLKBUF_X1 U3867 ( .A(n3752), .Z(n3737) );
  CLKBUF_X1 U3868 ( .A(n3751), .Z(n3738) );
  CLKBUF_X1 U3869 ( .A(n3751), .Z(n3739) );
  CLKBUF_X1 U3870 ( .A(n3751), .Z(n3740) );
  CLKBUF_X1 U3871 ( .A(n3751), .Z(n3741) );
  CLKBUF_X1 U3872 ( .A(n3751), .Z(n3742) );
  CLKBUF_X1 U3873 ( .A(n3751), .Z(n3743) );
  CLKBUF_X1 U3874 ( .A(n3750), .Z(n3744) );
  CLKBUF_X1 U3875 ( .A(n3750), .Z(n3745) );
  CLKBUF_X1 U3876 ( .A(n3750), .Z(n3746) );
  CLKBUF_X1 U3877 ( .A(n3750), .Z(n3747) );
  CLKBUF_X1 U3878 ( .A(n3750), .Z(n3748) );
  CLKBUF_X1 U3879 ( .A(n3750), .Z(n3749) );
  INV_X2 U3880 ( .A(CLK), .ZN(n4272) );
endmodule


module REG_PIPO_6_00_00_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n4, n5, n6, n7, n8, n3, n9, n10, n11, n12, n13, n14;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n14), .ZN(n2) );
  INV_X1 U3 ( .A(n1), .ZN(n13) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n2), .B1(n14), .B2(DOUT[0]), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(n12) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n2), .B1(n14), .B2(DOUT[1]), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n11) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n2), .B1(n14), .B2(DOUT[2]), .ZN(n5) );
  INV_X1 U9 ( .A(n6), .ZN(n10) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n2), .B1(n14), .B2(DOUT[3]), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n9) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n2), .B1(n14), .B2(DOUT[4]), .ZN(n7) );
  INV_X1 U13 ( .A(n8), .ZN(n3) );
  AOI22_X1 U14 ( .A1(DIN[5]), .A2(n2), .B1(n14), .B2(DOUT[5]), .ZN(n8) );
  INV_X1 U15 ( .A(EN), .ZN(n14) );
endmodule


module REG_PIPO_32_00000000_00000000_10 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_9 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_8 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_7 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n3) );
  BUF_X1 U4 ( .A(n169), .Z(n2) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n9), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n9) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n10), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n10) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n11), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n11) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n13), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n13) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n14), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n14) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n15), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U29 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U30 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U31 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U32 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U33 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U35 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U37 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U38 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U39 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U40 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U41 ( .A(DIN[21]), .ZN(n19) );
  OAI22_X1 U42 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U43 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U44 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U45 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U46 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U47 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U48 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U49 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U50 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U51 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U52 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U53 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U54 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U55 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U56 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U57 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U58 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U59 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U60 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U61 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U62 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U63 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U64 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U65 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U66 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U67 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U68 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U69 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U70 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U71 ( .A(DIN[10]), .ZN(n30) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_5_00_00_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n2, n4, n5, n6, n7, n3, n8, n9, n10, n11, n12;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n12), .ZN(n2) );
  INV_X1 U3 ( .A(n1), .ZN(n11) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n2), .B1(n12), .B2(DOUT[0]), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(n10) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n2), .B1(n12), .B2(DOUT[1]), .ZN(n4) );
  INV_X1 U7 ( .A(n5), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n2), .B1(n12), .B2(DOUT[2]), .ZN(n5) );
  INV_X1 U9 ( .A(n6), .ZN(n8) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n2), .B1(n12), .B2(DOUT[3]), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n3) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n2), .B1(n12), .B2(DOUT[4]), .ZN(n7) );
  INV_X1 U13 ( .A(EN), .ZN(n12) );
endmodule


module REG_PIPO_5_00_00_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(n11) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  INV_X1 U5 ( .A(n16), .ZN(n10) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  INV_X1 U9 ( .A(n14), .ZN(n8) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  INV_X1 U11 ( .A(n13), .ZN(n3) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  INV_X1 U13 ( .A(EN), .ZN(n12) );
endmodule


module ALU_DATA_W32_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   net21771, net21770, net21751, net21743, net21739, net21736, net21735,
         net21734, net21732, net21729, net21728, net21724, net21720, net21718,
         net21715, net21712, net21710, net21709, net21708, net21702, net21695,
         net21694, net21692, net21690, net21687, net21684, net21682, net21673,
         net21670, net21669, net21668, net21665, net21663, net21660, net21659,
         net21658, net21657, net21656, net21653, net21651, net21650, net21649,
         net21648, net21646, net21644, net21632, net21627, net21624, net21623,
         net21616, net21613, net21612, net21611, net21610, net21609, net21608,
         net21607, net21606, net21605, net21604, net21602, net21601, net21596,
         net21594, net21587, net21584, net21582, net21581, net21579, net21578,
         net21576, net21566, net21537, net21530, net21527, net21526, net21522,
         net21520, net21517, net21513, net21511, net21506, net21500, net21498,
         net21495, net27471, net27508, net28036, net34301, net34352, net34468,
         net34470, net34481, net34559, net34572, net34592, net34610, net34647,
         net34649, net34660, net34670, net34669, net34711, net34734, net34761,
         net34823, net34828, net34839, net34841, net34845, net34851, net34952,
         net35034, net35222, net36957, net37090, net38513, net38998, net39083,
         net38525, net36964, net41309, net21580, net21574, net21571, net21568,
         net21600, net21599, net37054, net21643, net21641, net21639, net21638,
         net21637, net21635, net21629, net21628, net21598, net33827, net21654,
         net38526, net35166, net34853, net34782, net34658, net34496, net21689,
         net21677, net21676, net41055, net41052, net28037, net21782, net21781,
         net21777, net21776, net21775, net21704, net21703, net21696, net21683,
         net21675, net37086, net37084, net37070, net37069, net37068, net37066,
         net37033, net21567, net21564, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161;

  CLKBUF_X1 U3 ( .A(net21665), .Z(n1) );
  NOR2_X1 U4 ( .A1(net21566), .A2(n38), .ZN(net37069) );
  INV_X1 U5 ( .A(net21594), .ZN(n38) );
  NAND2_X1 U6 ( .A1(A[28]), .A2(n39), .ZN(net37084) );
  INV_X1 U7 ( .A(B[28]), .ZN(n39) );
  INV_X1 U8 ( .A(B[30]), .ZN(n66) );
  NAND2_X1 U9 ( .A1(B[29]), .A2(n31), .ZN(n27) );
  INV_X1 U10 ( .A(A[29]), .ZN(n31) );
  INV_X1 U11 ( .A(B[29]), .ZN(n30) );
  NAND2_X1 U12 ( .A1(B[30]), .A2(n67), .ZN(net37054) );
  INV_X1 U13 ( .A(A[30]), .ZN(n67) );
  INV_X1 U14 ( .A(n20), .ZN(net21735) );
  INV_X1 U15 ( .A(n18), .ZN(n100) );
  INV_X1 U16 ( .A(net38998), .ZN(net21695) );
  INV_X1 U17 ( .A(n17), .ZN(net21694) );
  OAI21_X1 U18 ( .B1(net34669), .B2(net21566), .A(net37090), .ZN(net27471) );
  NOR2_X1 U19 ( .A1(net37033), .A2(n3), .ZN(net34352) );
  INV_X1 U20 ( .A(net37084), .ZN(net37033) );
  NOR2_X1 U21 ( .A1(n2), .A2(n65), .ZN(net21537) );
  NOR2_X1 U22 ( .A1(n66), .A2(A[30]), .ZN(n65) );
  AND2_X1 U23 ( .A1(A[30]), .A2(n66), .ZN(n2) );
  AND2_X1 U24 ( .A1(B[28]), .A2(net21564), .ZN(n3) );
  AND2_X1 U25 ( .A1(n30), .A2(A[29]), .ZN(n4) );
  AND2_X1 U26 ( .A1(net21735), .A2(net34572), .ZN(n5) );
  XOR2_X1 U27 ( .A(B[29]), .B(A[29]), .Z(n6) );
  AND2_X1 U28 ( .A1(net21594), .A2(net21576), .ZN(n7) );
  INV_X1 U29 ( .A(n9), .ZN(n8) );
  AND2_X1 U30 ( .A1(net36957), .A2(net21682), .ZN(n9) );
  NAND2_X1 U31 ( .A1(n82), .A2(n10), .ZN(net21584) );
  AND2_X1 U32 ( .A1(n83), .A2(net21578), .ZN(n10) );
  AND2_X1 U33 ( .A1(n82), .A2(n11), .ZN(net38525) );
  AND2_X1 U34 ( .A1(n83), .A2(net21578), .ZN(n11) );
  CLKBUF_X1 U35 ( .A(n106), .Z(n12) );
  AOI21_X1 U36 ( .B1(net21781), .B2(net21770), .A(net21782), .ZN(n13) );
  OAI21_X1 U37 ( .B1(net37068), .B2(n3), .A(net37084), .ZN(n14) );
  AND3_X1 U38 ( .A1(net21771), .A2(net21770), .A3(net21530), .ZN(net34649) );
  XNOR2_X1 U39 ( .A(n16), .B(n15), .ZN(DIFF[22]) );
  AND2_X1 U40 ( .A1(net21607), .A2(net21613), .ZN(n15) );
  AND2_X1 U41 ( .A1(net21623), .A2(net21611), .ZN(n16) );
  AND2_X1 U42 ( .A1(A[13]), .A2(net21724), .ZN(n17) );
  AND2_X1 U43 ( .A1(A[7]), .A2(n156), .ZN(n18) );
  INV_X1 U44 ( .A(n140), .ZN(n19) );
  NOR2_X1 U45 ( .A1(n92), .A2(B[10]), .ZN(n20) );
  NAND2_X1 U46 ( .A1(net27508), .A2(n23), .ZN(n21) );
  NAND2_X1 U47 ( .A1(n21), .A2(n22), .ZN(n80) );
  OR2_X1 U48 ( .A1(net21610), .A2(net21609), .ZN(n22) );
  AND2_X1 U49 ( .A1(net21612), .A2(net21611), .ZN(n23) );
  XNOR2_X1 U50 ( .A(n24), .B(n25), .ZN(DIFF[31]) );
  NAND2_X1 U51 ( .A1(n29), .A2(n28), .ZN(n24) );
  XOR2_X1 U52 ( .A(B[31]), .B(A[31]), .Z(n25) );
  BUF_X1 U53 ( .A(net21598), .Z(net27508) );
  AOI21_X1 U54 ( .B1(n20), .B2(net21732), .A(n77), .ZN(n26) );
  AOI21_X2 U55 ( .B1(n4), .B2(net37054), .A(n2), .ZN(n28) );
  NAND3_X1 U56 ( .A1(net37086), .A2(net37054), .A3(n27), .ZN(n29) );
  AOI21_X1 U57 ( .B1(n14), .B2(n27), .A(n4), .ZN(net39083) );
  OAI21_X1 U58 ( .B1(net37068), .B2(n3), .A(net37084), .ZN(net37086) );
  INV_X1 U59 ( .A(A[28]), .ZN(net21564) );
  AOI21_X1 U60 ( .B1(net37070), .B2(net37069), .A(net37066), .ZN(net37068) );
  INV_X1 U61 ( .A(net21567), .ZN(net37066) );
  INV_X1 U62 ( .A(net37066), .ZN(net37090) );
  AOI21_X1 U63 ( .B1(net21568), .B2(n32), .A(n33), .ZN(net21567) );
  INV_X1 U64 ( .A(net21571), .ZN(n33) );
  OAI21_X1 U65 ( .B1(n34), .B2(n35), .A(net21574), .ZN(n32) );
  INV_X1 U66 ( .A(net21580), .ZN(n35) );
  OAI21_X1 U67 ( .B1(net38525), .B2(n35), .A(net21574), .ZN(net21582) );
  AOI21_X1 U68 ( .B1(n36), .B2(net21576), .A(n37), .ZN(n34) );
  INV_X1 U69 ( .A(net21578), .ZN(n37) );
  INV_X1 U70 ( .A(net21579), .ZN(n36) );
  OAI21_X1 U71 ( .B1(net21599), .B2(net21598), .A(net21600), .ZN(net37070) );
  NAND3_X1 U72 ( .A1(net21580), .A2(net21568), .A3(net21576), .ZN(net21566) );
  NAND3_X1 U73 ( .A1(net21696), .A2(net28037), .A3(n45), .ZN(net21675) );
  CLKBUF_X1 U74 ( .A(net21675), .Z(net34782) );
  AND4_X1 U75 ( .A1(net38526), .A2(net21675), .A3(net21677), .A4(net21676), 
        .ZN(net34496) );
  NOR2_X1 U76 ( .A1(n40), .A2(net21683), .ZN(n45) );
  NAND2_X1 U77 ( .A1(net21776), .A2(n13), .ZN(net21696) );
  NAND4_X1 U78 ( .A1(net21777), .A2(net33827), .A3(net21530), .A4(net21770), 
        .ZN(net21776) );
  NAND2_X1 U79 ( .A1(net41055), .A2(net21654), .ZN(net21777) );
  AND4_X2 U80 ( .A1(net21520), .A2(net21513), .A3(net21506), .A4(net35034), 
        .ZN(net28037) );
  AOI21_X1 U81 ( .B1(net21522), .B2(net28037), .A(net34851), .ZN(net34468) );
  NAND4_X1 U82 ( .A1(net34853), .A2(net34649), .A3(net28036), .A4(net28037), 
        .ZN(net21677) );
  NAND4_X1 U83 ( .A1(net21732), .A2(net21736), .A3(net21495), .A4(net21500), 
        .ZN(net21683) );
  NAND2_X1 U84 ( .A1(B[15]), .A2(n41), .ZN(net21684) );
  INV_X1 U85 ( .A(A[15]), .ZN(n41) );
  NAND2_X1 U86 ( .A1(B[13]), .A2(n43), .ZN(net21692) );
  INV_X1 U87 ( .A(A[13]), .ZN(n43) );
  NAND2_X1 U88 ( .A1(B[14]), .A2(n42), .ZN(net21704) );
  INV_X1 U89 ( .A(net21704), .ZN(net21689) );
  NAND4_X1 U90 ( .A1(net21703), .A2(net21692), .A3(net21704), .A4(net21684), 
        .ZN(n40) );
  AND4_X1 U91 ( .A1(net21703), .A2(net21692), .A3(net21704), .A4(net21684), 
        .ZN(net34853) );
  INV_X1 U92 ( .A(A[14]), .ZN(n42) );
  NAND2_X1 U93 ( .A1(B[12]), .A2(n44), .ZN(net21703) );
  INV_X1 U94 ( .A(net21703), .ZN(net21720) );
  INV_X1 U95 ( .A(A[12]), .ZN(n44) );
  AOI21_X1 U96 ( .B1(net21781), .B2(net21770), .A(net21782), .ZN(net21775) );
  AND2_X1 U97 ( .A1(net36964), .A2(net21775), .ZN(net36957) );
  INV_X1 U98 ( .A(net21526), .ZN(net21782) );
  INV_X1 U99 ( .A(net21527), .ZN(net21781) );
  NAND2_X1 U100 ( .A1(B[1]), .A2(net41052), .ZN(net33827) );
  OR2_X1 U101 ( .A1(B[1]), .A2(net41052), .ZN(net41055) );
  CLKBUF_X1 U102 ( .A(net41055), .Z(net34559) );
  INV_X1 U103 ( .A(A[1]), .ZN(net41052) );
  CLKBUF_X1 U104 ( .A(net34496), .Z(net34711) );
  OAI21_X1 U105 ( .B1(net34496), .B2(net21635), .A(net21637), .ZN(net21628) );
  AOI22_X1 U106 ( .A1(n49), .A2(net34853), .B1(net21702), .B2(n45), .ZN(
        net38526) );
  CLKBUF_X1 U107 ( .A(net38526), .Z(net34658) );
  OAI21_X1 U108 ( .B1(net21728), .B2(net21729), .A(n26), .ZN(n49) );
  AOI21_X1 U109 ( .B1(n46), .B2(net21684), .A(n47), .ZN(net21676) );
  CLKBUF_X1 U110 ( .A(net21676), .Z(net35166) );
  INV_X1 U111 ( .A(net21687), .ZN(n47) );
  OAI21_X1 U112 ( .B1(n48), .B2(net21689), .A(net21690), .ZN(n46) );
  INV_X1 U113 ( .A(net21689), .ZN(net41309) );
  OAI21_X1 U114 ( .B1(net21709), .B2(net21689), .A(net21690), .ZN(net21708) );
  AOI21_X1 U115 ( .B1(net38998), .B2(net21692), .A(n17), .ZN(n48) );
  NAND4_X1 U116 ( .A1(net21677), .A2(net34658), .A3(net35166), .A4(net34782), 
        .ZN(net21670) );
  CLKBUF_X1 U117 ( .A(net21702), .Z(net34851) );
  CLKBUF_X1 U118 ( .A(net21728), .Z(net34841) );
  CLKBUF_X1 U119 ( .A(net33827), .Z(net34828) );
  NAND4_X1 U120 ( .A1(net21777), .A2(net33827), .A3(net21530), .A4(net21770), 
        .ZN(net36964) );
  AND2_X1 U121 ( .A1(net33827), .A2(net21656), .ZN(net21771) );
  NAND2_X1 U122 ( .A1(B[2]), .A2(n50), .ZN(net21530) );
  INV_X1 U123 ( .A(A[2]), .ZN(n50) );
  NAND2_X1 U124 ( .A1(n51), .A2(B[3]), .ZN(net21770) );
  INV_X1 U125 ( .A(A[3]), .ZN(n51) );
  NAND2_X1 U126 ( .A1(n54), .A2(A[0]), .ZN(net21654) );
  CLKBUF_X1 U127 ( .A(net21654), .Z(net34823) );
  INV_X1 U128 ( .A(B[0]), .ZN(n54) );
  INV_X1 U129 ( .A(B[2]), .ZN(n52) );
  NAND2_X1 U130 ( .A1(n52), .A2(A[2]), .ZN(net21527) );
  OR2_X1 U131 ( .A1(n51), .A2(B[3]), .ZN(net21526) );
  INV_X1 U132 ( .A(A[0]), .ZN(n53) );
  NAND2_X1 U133 ( .A1(B[0]), .A2(n53), .ZN(net21656) );
  NAND2_X1 U134 ( .A1(net21628), .A2(net21629), .ZN(net21598) );
  OAI21_X1 U135 ( .B1(net21598), .B2(net21599), .A(net21600), .ZN(net34761) );
  AOI21_X1 U136 ( .B1(net21638), .B2(net21639), .A(n57), .ZN(net21637) );
  INV_X1 U137 ( .A(net21641), .ZN(n57) );
  AOI21_X1 U138 ( .B1(net21638), .B2(net21639), .A(n57), .ZN(n64) );
  NAND2_X1 U139 ( .A1(B[20]), .A2(n55), .ZN(net21629) );
  NAND2_X1 U140 ( .A1(net21612), .A2(net21629), .ZN(net21632) );
  INV_X1 U141 ( .A(n63), .ZN(n55) );
  CLKBUF_X1 U142 ( .A(A[20]), .Z(n63) );
  NAND4_X1 U143 ( .A1(net21638), .A2(net21650), .A3(net21651), .A4(net21646), 
        .ZN(net21635) );
  OAI21_X1 U144 ( .B1(net21635), .B2(net34711), .A(n64), .ZN(net34660) );
  NAND2_X1 U145 ( .A1(B[19]), .A2(n61), .ZN(net21638) );
  NAND2_X1 U146 ( .A1(net21641), .A2(net21638), .ZN(net21657) );
  INV_X1 U147 ( .A(A[19]), .ZN(n61) );
  OAI21_X1 U148 ( .B1(n58), .B2(net21643), .A(net21644), .ZN(net21639) );
  INV_X1 U149 ( .A(net21650), .ZN(net21643) );
  OAI21_X1 U150 ( .B1(net21659), .B2(net21643), .A(net21644), .ZN(net21658) );
  AOI21_X1 U151 ( .B1(n59), .B2(net21646), .A(n60), .ZN(n58) );
  INV_X1 U152 ( .A(net21648), .ZN(n60) );
  INV_X1 U153 ( .A(net21649), .ZN(n59) );
  NAND2_X1 U154 ( .A1(A[19]), .A2(n62), .ZN(net21641) );
  INV_X1 U155 ( .A(B[19]), .ZN(n62) );
  INV_X1 U156 ( .A(B[20]), .ZN(n56) );
  NAND2_X1 U157 ( .A1(A[20]), .A2(n56), .ZN(net21612) );
  NAND3_X1 U158 ( .A1(net21613), .A2(net21601), .A3(net21609), .ZN(net21599)
         );
  OAI21_X1 U159 ( .B1(net27508), .B2(net21599), .A(n69), .ZN(net34301) );
  AOI21_X1 U160 ( .B1(net21601), .B2(net21602), .A(n68), .ZN(net21600) );
  INV_X1 U161 ( .A(net21604), .ZN(n68) );
  AOI21_X1 U162 ( .B1(net21601), .B2(net21602), .A(n68), .ZN(n69) );
  INV_X1 U163 ( .A(net21613), .ZN(net21606) );
  NAND2_X1 U164 ( .A1(net21604), .A2(net21601), .ZN(net21616) );
  NAND2_X1 U165 ( .A1(net21611), .A2(net21609), .ZN(net21627) );
  NAND2_X1 U166 ( .A1(net21624), .A2(net21609), .ZN(net21623) );
  AOI21_X1 U167 ( .B1(net21608), .B2(net21609), .A(net21610), .ZN(net21605) );
  NAND2_X1 U168 ( .A1(net21644), .A2(net21650), .ZN(net21663) );
  INV_X1 U169 ( .A(net21651), .ZN(net21669) );
  NAND2_X1 U170 ( .A1(net21649), .A2(net21651), .ZN(net21673) );
  NAND2_X1 U171 ( .A1(net21648), .A2(net21646), .ZN(net21668) );
  NAND2_X1 U172 ( .A1(net21646), .A2(net21665), .ZN(n70) );
  NAND2_X1 U173 ( .A1(n70), .A2(net21648), .ZN(net21660) );
  NAND2_X1 U174 ( .A1(B[27]), .A2(n71), .ZN(net21568) );
  NAND2_X1 U175 ( .A1(net21571), .A2(net21568), .ZN(net21581) );
  INV_X1 U176 ( .A(A[27]), .ZN(n71) );
  NAND2_X1 U177 ( .A1(A[27]), .A2(n72), .ZN(net21571) );
  INV_X1 U178 ( .A(B[27]), .ZN(n72) );
  NAND2_X1 U179 ( .A1(A[26]), .A2(n74), .ZN(net21574) );
  NAND2_X1 U180 ( .A1(net21574), .A2(net21580), .ZN(net21587) );
  INV_X1 U181 ( .A(B[26]), .ZN(n74) );
  NAND2_X1 U182 ( .A1(B[26]), .A2(n73), .ZN(net21580) );
  INV_X1 U183 ( .A(A[26]), .ZN(n73) );
  NAND2_X1 U184 ( .A1(B[25]), .A2(n75), .ZN(net21576) );
  INV_X1 U185 ( .A(A[25]), .ZN(n75) );
  NAND2_X1 U186 ( .A1(A[25]), .A2(net21596), .ZN(net21578) );
  CLKBUF_X1 U187 ( .A(n107), .Z(n76) );
  INV_X1 U188 ( .A(net21734), .ZN(n77) );
  AND2_X1 U189 ( .A1(A[12]), .A2(net21739), .ZN(net38998) );
  OAI21_X1 U190 ( .B1(net21720), .B2(n139), .A(net21695), .ZN(n78) );
  INV_X1 U191 ( .A(n139), .ZN(n79) );
  INV_X1 U192 ( .A(net21715), .ZN(net38513) );
  NAND2_X1 U193 ( .A1(net34761), .A2(net21594), .ZN(net34669) );
  CLKBUF_X1 U194 ( .A(n96), .Z(n81) );
  INV_X1 U195 ( .A(net34649), .ZN(net21682) );
  NAND2_X1 U196 ( .A1(net34761), .A2(n7), .ZN(n82) );
  OR2_X1 U197 ( .A1(net35222), .A2(net21579), .ZN(n83) );
  INV_X1 U198 ( .A(net21576), .ZN(net35222) );
  CLKBUF_X1 U199 ( .A(B[4]), .Z(n84) );
  OR2_X1 U200 ( .A1(n156), .A2(A[7]), .ZN(net35034) );
  CLKBUF_X1 U201 ( .A(n26), .Z(net34952) );
  OR2_X1 U202 ( .A1(n160), .A2(B[4]), .ZN(n107) );
  OR2_X1 U203 ( .A1(n156), .A2(A[7]), .ZN(n99) );
  CLKBUF_X1 U204 ( .A(net21495), .Z(net34845) );
  CLKBUF_X1 U205 ( .A(A[14]), .Z(net34839) );
  CLKBUF_X1 U206 ( .A(n94), .Z(n85) );
  INV_X1 U207 ( .A(net21653), .ZN(net34734) );
  CLKBUF_X1 U208 ( .A(net21684), .Z(net34670) );
  OAI21_X1 U209 ( .B1(net34841), .B2(net21729), .A(net34952), .ZN(n86) );
  INV_X1 U210 ( .A(net21720), .ZN(net34647) );
  INV_X1 U211 ( .A(net28036), .ZN(net34610) );
  CLKBUF_X1 U212 ( .A(net21500), .Z(net34592) );
  OR2_X1 U213 ( .A1(n161), .A2(B[9]), .ZN(n94) );
  OR2_X1 U214 ( .A1(n147), .A2(B[11]), .ZN(net21734) );
  INV_X1 U215 ( .A(net21743), .ZN(net34572) );
  CLKBUF_X1 U216 ( .A(n104), .Z(n87) );
  INV_X1 U217 ( .A(net34468), .ZN(net21498) );
  CLKBUF_X1 U218 ( .A(net21513), .Z(net34481) );
  INV_X1 U219 ( .A(net21709), .ZN(net34470) );
  XOR2_X1 U220 ( .A(n88), .B(n8), .Z(DIFF[4]) );
  AND2_X1 U221 ( .A1(n76), .A2(net21520), .ZN(n88) );
  XOR2_X1 U222 ( .A(n89), .B(n101), .Z(DIFF[6]) );
  AND2_X1 U223 ( .A1(net21506), .A2(n12), .ZN(n89) );
  XOR2_X1 U224 ( .A(n97), .B(n98), .Z(DIFF[7]) );
  XNOR2_X1 U225 ( .A(n93), .B(n90), .ZN(DIFF[9]) );
  AND2_X1 U226 ( .A1(net34845), .A2(n85), .ZN(n90) );
  XOR2_X1 U227 ( .A(net27471), .B(net34352), .Z(DIFF[28]) );
  XNOR2_X1 U228 ( .A(net21624), .B(net21627), .ZN(DIFF[21]) );
  XNOR2_X1 U229 ( .A(net21663), .B(net21660), .ZN(DIFF[18]) );
  XNOR2_X1 U230 ( .A(net21668), .B(n1), .ZN(DIFF[17]) );
  XNOR2_X1 U231 ( .A(net21658), .B(net21657), .ZN(DIFF[19]) );
  XNOR2_X1 U232 ( .A(net21584), .B(net21587), .ZN(DIFF[26]) );
  NAND2_X1 U233 ( .A1(net21687), .A2(net34670), .ZN(n134) );
  XNOR2_X1 U234 ( .A(n135), .B(net34470), .ZN(DIFF[14]) );
  NAND2_X1 U235 ( .A1(net21690), .A2(net41309), .ZN(n135) );
  AOI21_X1 U236 ( .B1(net21506), .B2(n101), .A(n102), .ZN(n97) );
  XOR2_X1 U237 ( .A(n91), .B(n105), .Z(DIFF[5]) );
  AND2_X1 U238 ( .A1(net34481), .A2(n87), .ZN(n91) );
  XNOR2_X1 U239 ( .A(n141), .B(n79), .ZN(DIFF[12]) );
  NAND2_X1 U240 ( .A1(net21695), .A2(net34647), .ZN(n141) );
  XNOR2_X1 U241 ( .A(n6), .B(n14), .ZN(DIFF[29]) );
  OAI21_X1 U242 ( .B1(n103), .B2(net21511), .A(n87), .ZN(n101) );
  OAI21_X1 U243 ( .B1(n136), .B2(net21715), .A(net21694), .ZN(net21710) );
  XNOR2_X1 U244 ( .A(n112), .B(n111), .ZN(DIFF[2]) );
  NAND2_X1 U245 ( .A1(net21530), .A2(net21527), .ZN(n112) );
  XNOR2_X1 U246 ( .A(n108), .B(n109), .ZN(DIFF[3]) );
  XNOR2_X1 U247 ( .A(n127), .B(n114), .ZN(DIFF[1]) );
  OAI21_X1 U248 ( .B1(net21720), .B2(n19), .A(net21695), .ZN(n137) );
  OAI21_X1 U249 ( .B1(n146), .B2(net21743), .A(net21735), .ZN(n145) );
  OAI21_X1 U250 ( .B1(net21605), .B2(net21606), .A(net21607), .ZN(net21602) );
  NAND2_X1 U251 ( .A1(net27508), .A2(net21612), .ZN(net21624) );
  AOI21_X1 U252 ( .B1(n102), .B2(n99), .A(n18), .ZN(n152) );
  OAI21_X1 U253 ( .B1(net21751), .B2(n93), .A(n85), .ZN(n148) );
  XNOR2_X1 U254 ( .A(net39083), .B(net21537), .ZN(DIFF[30]) );
  NAND2_X1 U255 ( .A1(net21578), .A2(net21576), .ZN(n116) );
  NAND2_X1 U256 ( .A1(net21579), .A2(net21594), .ZN(n117) );
  NAND2_X1 U257 ( .A1(net21527), .A2(n110), .ZN(n108) );
  NAND2_X1 U258 ( .A1(n111), .A2(net21530), .ZN(n110) );
  NAND2_X1 U259 ( .A1(net35034), .A2(n100), .ZN(n98) );
  NAND2_X1 U260 ( .A1(net21653), .A2(net34823), .ZN(n114) );
  INV_X1 U261 ( .A(net21656), .ZN(net21653) );
  INV_X1 U262 ( .A(B[18]), .ZN(n129) );
  INV_X1 U263 ( .A(B[25]), .ZN(net21596) );
  NAND2_X1 U264 ( .A1(A[24]), .A2(n119), .ZN(net21579) );
  INV_X1 U265 ( .A(B[24]), .ZN(n119) );
  NAND2_X1 U266 ( .A1(A[21]), .A2(n126), .ZN(net21611) );
  NAND2_X1 U267 ( .A1(A[22]), .A2(n124), .ZN(net21607) );
  NAND2_X1 U268 ( .A1(A[16]), .A2(n133), .ZN(net21649) );
  INV_X1 U269 ( .A(B[16]), .ZN(n133) );
  NAND2_X1 U270 ( .A1(A[23]), .A2(n122), .ZN(net21604) );
  INV_X1 U271 ( .A(B[23]), .ZN(n122) );
  NAND2_X1 U272 ( .A1(B[16]), .A2(n132), .ZN(net21651) );
  INV_X1 U273 ( .A(A[16]), .ZN(n132) );
  NAND2_X1 U274 ( .A1(B[23]), .A2(n121), .ZN(net21601) );
  INV_X1 U275 ( .A(A[23]), .ZN(n121) );
  INV_X1 U276 ( .A(A[10]), .ZN(n92) );
  NAND2_X1 U277 ( .A1(B[24]), .A2(n118), .ZN(net21594) );
  INV_X1 U278 ( .A(A[24]), .ZN(n118) );
  NAND2_X1 U279 ( .A1(B[17]), .A2(n130), .ZN(net21646) );
  INV_X1 U280 ( .A(A[21]), .ZN(n125) );
  INV_X1 U281 ( .A(A[22]), .ZN(n123) );
  INV_X1 U282 ( .A(B[17]), .ZN(n131) );
  OAI21_X1 U283 ( .B1(net34468), .B2(net34610), .A(n142), .ZN(n140) );
  AND2_X1 U284 ( .A1(n149), .A2(n81), .ZN(n93) );
  NAND2_X1 U285 ( .A1(n94), .A2(n96), .ZN(n143) );
  XNOR2_X1 U286 ( .A(net21708), .B(n134), .ZN(DIFF[15]) );
  NAND2_X1 U287 ( .A1(B[22]), .A2(n123), .ZN(net21613) );
  INV_X1 U288 ( .A(B[22]), .ZN(n124) );
  NAND2_X1 U289 ( .A1(A[6]), .A2(n157), .ZN(n106) );
  NAND2_X1 U290 ( .A1(net36957), .A2(net21682), .ZN(net21522) );
  NAND2_X1 U291 ( .A1(B[21]), .A2(n125), .ZN(net21609) );
  INV_X1 U292 ( .A(B[21]), .ZN(n126) );
  NAND2_X1 U293 ( .A1(A[17]), .A2(n131), .ZN(net21648) );
  INV_X1 U294 ( .A(A[17]), .ZN(n130) );
  NAND4_X1 U295 ( .A1(n154), .A2(net21513), .A3(net21506), .A4(n99), .ZN(n153)
         );
  OAI21_X1 U296 ( .B1(net21669), .B2(net34711), .A(net21649), .ZN(net21665) );
  INV_X1 U297 ( .A(B[13]), .ZN(net21724) );
  INV_X1 U298 ( .A(B[6]), .ZN(n157) );
  INV_X1 U299 ( .A(B[15]), .ZN(net21712) );
  INV_X1 U300 ( .A(B[5]), .ZN(n155) );
  NAND2_X1 U301 ( .A1(n84), .A2(n160), .ZN(net21520) );
  INV_X1 U302 ( .A(B[8]), .ZN(n150) );
  INV_X1 U303 ( .A(B[12]), .ZN(net21739) );
  NAND2_X1 U304 ( .A1(net34839), .A2(net21718), .ZN(net21690) );
  NAND2_X1 U305 ( .A1(B[11]), .A2(n147), .ZN(net21732) );
  XNOR2_X1 U306 ( .A(net34660), .B(net21632), .ZN(DIFF[20]) );
  INV_X1 U307 ( .A(B[14]), .ZN(net21718) );
  NAND2_X1 U308 ( .A1(n152), .A2(n153), .ZN(net21702) );
  OAI21_X1 U309 ( .B1(n80), .B2(net21606), .A(net21607), .ZN(n120) );
  NAND2_X1 U310 ( .A1(B[5]), .A2(n159), .ZN(net21513) );
  XNOR2_X1 U311 ( .A(n120), .B(net21616), .ZN(DIFF[23]) );
  NAND2_X1 U312 ( .A1(net38513), .A2(net21694), .ZN(n138) );
  AND4_X1 U313 ( .A1(net21732), .A2(net21736), .A3(net21495), .A4(net21500), 
        .ZN(net28036) );
  NAND2_X1 U314 ( .A1(n143), .A2(net21736), .ZN(net21728) );
  NAND2_X1 U315 ( .A1(B[10]), .A2(n92), .ZN(net21736) );
  NAND2_X1 U316 ( .A1(n113), .A2(net34559), .ZN(n111) );
  NAND2_X1 U317 ( .A1(net21734), .A2(net21732), .ZN(n144) );
  NAND2_X1 U318 ( .A1(net21732), .A2(net21495), .ZN(net21729) );
  NAND2_X1 U319 ( .A1(A[18]), .A2(n129), .ZN(net21644) );
  NAND2_X1 U320 ( .A1(A[8]), .A2(n150), .ZN(n96) );
  XNOR2_X1 U321 ( .A(n116), .B(n115), .ZN(DIFF[25]) );
  OAI21_X1 U322 ( .B1(net21517), .B2(n9), .A(n76), .ZN(n105) );
  NAND2_X1 U323 ( .A1(n104), .A2(n107), .ZN(n154) );
  INV_X1 U324 ( .A(B[7]), .ZN(n156) );
  NAND2_X1 U325 ( .A1(net34823), .A2(net34734), .ZN(DIFF[0]) );
  NAND2_X1 U326 ( .A1(net34828), .A2(net34559), .ZN(n127) );
  NAND2_X1 U327 ( .A1(net34828), .A2(n114), .ZN(n113) );
  NAND2_X1 U328 ( .A1(B[18]), .A2(n128), .ZN(net21650) );
  INV_X1 U329 ( .A(A[18]), .ZN(n128) );
  NAND2_X1 U330 ( .A1(net21498), .A2(net34592), .ZN(n149) );
  NAND2_X1 U331 ( .A1(n81), .A2(net34592), .ZN(n95) );
  NAND2_X1 U332 ( .A1(B[8]), .A2(n151), .ZN(net21500) );
  INV_X1 U333 ( .A(A[5]), .ZN(n159) );
  NAND2_X1 U334 ( .A1(A[5]), .A2(n155), .ZN(n104) );
  INV_X1 U335 ( .A(A[9]), .ZN(n161) );
  NAND2_X1 U336 ( .A1(B[6]), .A2(n158), .ZN(net21506) );
  INV_X1 U337 ( .A(A[6]), .ZN(n158) );
  NAND2_X1 U338 ( .A1(n161), .A2(B[9]), .ZN(net21495) );
  INV_X1 U339 ( .A(A[4]), .ZN(n160) );
  INV_X1 U340 ( .A(A[8]), .ZN(n151) );
  NAND2_X1 U341 ( .A1(A[15]), .A2(net21712), .ZN(net21687) );
  NAND2_X1 U342 ( .A1(net21770), .A2(net21526), .ZN(n109) );
  NAND2_X1 U343 ( .A1(net34669), .A2(net21579), .ZN(n115) );
  INV_X1 U344 ( .A(A[11]), .ZN(n147) );
  XNOR2_X1 U345 ( .A(n95), .B(net21498), .ZN(DIFF[8]) );
  INV_X1 U346 ( .A(net34481), .ZN(net21511) );
  INV_X1 U347 ( .A(n105), .ZN(n103) );
  INV_X1 U348 ( .A(net21520), .ZN(net21517) );
  XNOR2_X1 U349 ( .A(net21582), .B(net21581), .ZN(DIFF[27]) );
  XNOR2_X1 U350 ( .A(n117), .B(net34301), .ZN(DIFF[24]) );
  INV_X1 U351 ( .A(net21611), .ZN(net21610) );
  INV_X1 U352 ( .A(net21612), .ZN(net21608) );
  INV_X1 U353 ( .A(net21660), .ZN(net21659) );
  XNOR2_X1 U354 ( .A(net21673), .B(net21670), .ZN(DIFF[16]) );
  INV_X1 U355 ( .A(net21710), .ZN(net21709) );
  INV_X1 U356 ( .A(net21692), .ZN(net21715) );
  INV_X1 U357 ( .A(n137), .ZN(n136) );
  XNOR2_X1 U358 ( .A(n78), .B(n138), .ZN(DIFF[13]) );
  INV_X1 U359 ( .A(n140), .ZN(n139) );
  INV_X1 U360 ( .A(n86), .ZN(n142) );
  XNOR2_X1 U361 ( .A(n145), .B(n144), .ZN(DIFF[11]) );
  INV_X1 U362 ( .A(net21736), .ZN(net21743) );
  XNOR2_X1 U363 ( .A(n146), .B(n5), .ZN(DIFF[10]) );
  INV_X1 U364 ( .A(n148), .ZN(n146) );
  INV_X1 U365 ( .A(n106), .ZN(n102) );
  INV_X1 U366 ( .A(net34845), .ZN(net21751) );
endmodule


module ALU_DATA_W32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   net22688, net22680, net22672, net22671, net22669, net22666, net22663,
         net22661, net22658, net22657, net22656, net22655, net22647, net22641,
         net22640, net22638, net22631, net22628, net22610, net22600, net22599,
         net22595, net22589, net27463, net28033, net33637, net34472, net34522,
         net34521, net34713, net36853, net37671, net37670, net37669, net34690,
         net34666, net34455, net37913, net38000, net37985, net37967, net37948,
         net37947, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274;

  BUF_X1 U2 ( .A(n232), .Z(n108) );
  OR2_X1 U3 ( .A1(A[14]), .A2(B[14]), .ZN(n214) );
  NOR2_X1 U4 ( .A1(net22599), .A2(n46), .ZN(n45) );
  INV_X1 U5 ( .A(net22628), .ZN(n46) );
  INV_X1 U6 ( .A(net22672), .ZN(n39) );
  INV_X1 U7 ( .A(n80), .ZN(net37671) );
  INV_X1 U8 ( .A(net37670), .ZN(net37948) );
  INV_X1 U9 ( .A(B[20]), .ZN(n31) );
  INV_X1 U10 ( .A(B[22]), .ZN(n27) );
  INV_X1 U11 ( .A(B[23]), .ZN(n25) );
  NAND2_X1 U12 ( .A1(n33), .A2(n34), .ZN(net22628) );
  INV_X1 U13 ( .A(A[24]), .ZN(n34) );
  INV_X1 U14 ( .A(n105), .ZN(n159) );
  INV_X1 U15 ( .A(n74), .ZN(n162) );
  INV_X1 U16 ( .A(n96), .ZN(n252) );
  NAND2_X1 U17 ( .A1(net37947), .A2(net37948), .ZN(net37669) );
  NOR2_X1 U18 ( .A1(n80), .A2(n81), .ZN(n82) );
  AND2_X1 U19 ( .A1(B[21]), .A2(A[21]), .ZN(n1) );
  AND2_X1 U20 ( .A1(n47), .A2(n48), .ZN(n2) );
  AND2_X1 U21 ( .A1(A[20]), .A2(B[20]), .ZN(n3) );
  AND2_X1 U22 ( .A1(n121), .A2(n269), .ZN(SUM[0]) );
  CLKBUF_X1 U23 ( .A(n268), .Z(n5) );
  CLKBUF_X1 U24 ( .A(n245), .Z(n6) );
  XNOR2_X1 U25 ( .A(n7), .B(n10), .ZN(SUM[29]) );
  AND2_X1 U26 ( .A1(n90), .A2(n91), .ZN(n7) );
  NAND2_X1 U27 ( .A1(n82), .A2(n2), .ZN(n77) );
  NAND2_X1 U28 ( .A1(n2), .A2(n57), .ZN(n75) );
  NAND2_X1 U29 ( .A1(net22657), .A2(n58), .ZN(net22655) );
  CLKBUF_X1 U30 ( .A(n199), .Z(n8) );
  AND2_X1 U31 ( .A1(n206), .A2(n199), .ZN(n9) );
  AND2_X1 U32 ( .A1(n92), .A2(n93), .ZN(n10) );
  INV_X1 U33 ( .A(B[24]), .ZN(n33) );
  INV_X1 U34 ( .A(n69), .ZN(n240) );
  OAI21_X1 U35 ( .B1(n42), .B2(n35), .A(n45), .ZN(n11) );
  AND2_X1 U36 ( .A1(n92), .A2(n93), .ZN(net34521) );
  NAND2_X1 U37 ( .A1(net34713), .A2(n77), .ZN(net28033) );
  CLKBUF_X1 U38 ( .A(n249), .Z(n106) );
  AND4_X1 U39 ( .A1(n60), .A2(net37913), .A3(net22663), .A4(n24), .ZN(n51) );
  NAND2_X1 U40 ( .A1(n11), .A2(n15), .ZN(n12) );
  NAND2_X1 U41 ( .A1(n12), .A2(n13), .ZN(n89) );
  OR2_X1 U42 ( .A1(n14), .A2(n94), .ZN(n13) );
  INV_X1 U43 ( .A(n93), .ZN(n14) );
  AND2_X1 U44 ( .A1(net22600), .A2(n93), .ZN(n15) );
  OR2_X1 U45 ( .A1(B[5]), .A2(A[5]), .ZN(n147) );
  NAND2_X1 U46 ( .A1(n31), .A2(n32), .ZN(n16) );
  CLKBUF_X1 U47 ( .A(n51), .Z(net38000) );
  BUF_X1 U48 ( .A(n19), .Z(net34472) );
  CLKBUF_X1 U49 ( .A(A[21]), .Z(n52) );
  NAND2_X1 U50 ( .A1(n112), .A2(n113), .ZN(n17) );
  CLKBUF_X1 U51 ( .A(net34666), .Z(n18) );
  NAND2_X1 U52 ( .A1(n208), .A2(n209), .ZN(n19) );
  INV_X1 U53 ( .A(B[21]), .ZN(n29) );
  XNOR2_X1 U54 ( .A(n20), .B(n122), .ZN(SUM[19]) );
  AND2_X1 U55 ( .A1(n203), .A2(n195), .ZN(n20) );
  XNOR2_X1 U56 ( .A(n21), .B(n22), .ZN(SUM[23]) );
  AND2_X1 U57 ( .A1(net22638), .A2(n76), .ZN(n21) );
  AND2_X1 U58 ( .A1(net22647), .A2(n61), .ZN(n22) );
  OR2_X1 U59 ( .A1(B[2]), .A2(A[2]), .ZN(n168) );
  OR2_X1 U60 ( .A1(B[12]), .A2(A[12]), .ZN(n228) );
  NAND2_X1 U61 ( .A1(n18), .A2(net22628), .ZN(n23) );
  NAND3_X1 U62 ( .A1(n51), .A2(net22672), .A3(n19), .ZN(n43) );
  INV_X1 U63 ( .A(net22680), .ZN(n41) );
  INV_X1 U64 ( .A(A[23]), .ZN(n26) );
  INV_X1 U65 ( .A(A[22]), .ZN(n28) );
  CLKBUF_X1 U66 ( .A(A[23]), .Z(n62) );
  INV_X1 U67 ( .A(A[20]), .ZN(n32) );
  NAND2_X1 U68 ( .A1(n26), .A2(n25), .ZN(n24) );
  NAND2_X1 U69 ( .A1(n49), .A2(n61), .ZN(n36) );
  NAND2_X1 U70 ( .A1(net22688), .A2(n41), .ZN(n40) );
  OR2_X1 U71 ( .A1(net22671), .A2(n40), .ZN(n47) );
  INV_X1 U72 ( .A(n3), .ZN(n59) );
  INV_X1 U73 ( .A(n52), .ZN(n30) );
  CLKBUF_X1 U74 ( .A(A[22]), .Z(n63) );
  NAND2_X1 U75 ( .A1(n27), .A2(n28), .ZN(n60) );
  INV_X1 U76 ( .A(n60), .ZN(n50) );
  INV_X1 U77 ( .A(n50), .ZN(net22641) );
  INV_X1 U78 ( .A(n1), .ZN(n58) );
  AOI21_X1 U79 ( .B1(n55), .B2(n3), .A(n1), .ZN(n38) );
  OAI21_X1 U80 ( .B1(n38), .B2(n50), .A(net22638), .ZN(n49) );
  NAND2_X1 U81 ( .A1(n51), .A2(n40), .ZN(n44) );
  AND2_X1 U82 ( .A1(n41), .A2(net22688), .ZN(net22669) );
  NOR2_X1 U83 ( .A1(n40), .A2(net22671), .ZN(n53) );
  OAI21_X1 U84 ( .B1(n42), .B2(n35), .A(n45), .ZN(n37) );
  NAND2_X1 U85 ( .A1(n37), .A2(net22600), .ZN(net34455) );
  NAND2_X1 U86 ( .A1(n29), .A2(n30), .ZN(n55) );
  NAND2_X1 U87 ( .A1(n29), .A2(n30), .ZN(net37913) );
  AND2_X1 U88 ( .A1(net22669), .A2(n39), .ZN(n54) );
  NOR2_X1 U89 ( .A1(n54), .A2(n53), .ZN(n56) );
  INV_X1 U90 ( .A(n54), .ZN(n48) );
  NOR2_X1 U91 ( .A1(net37985), .A2(n35), .ZN(net37967) );
  NAND2_X1 U92 ( .A1(n43), .A2(n44), .ZN(n42) );
  NAND2_X1 U93 ( .A1(n31), .A2(n32), .ZN(net22663) );
  CLKBUF_X1 U94 ( .A(n16), .Z(n57) );
  NAND2_X1 U95 ( .A1(net22647), .A2(n36), .ZN(n35) );
  NAND2_X1 U96 ( .A1(n25), .A2(n26), .ZN(net22640) );
  NAND2_X1 U97 ( .A1(n25), .A2(n26), .ZN(n61) );
  AND2_X1 U98 ( .A1(net22647), .A2(n36), .ZN(net34713) );
  CLKBUF_X1 U99 ( .A(n248), .Z(n64) );
  OR2_X1 U100 ( .A1(A[11]), .A2(B[11]), .ZN(n65) );
  CLKBUF_X1 U101 ( .A(n161), .Z(n66) );
  CLKBUF_X1 U102 ( .A(n130), .Z(n67) );
  CLKBUF_X1 U103 ( .A(n142), .Z(n68) );
  NAND2_X1 U104 ( .A1(n59), .A2(n75), .ZN(net22658) );
  NAND2_X1 U105 ( .A1(n59), .A2(n57), .ZN(net22666) );
  INV_X1 U106 ( .A(n59), .ZN(net37947) );
  AND2_X1 U107 ( .A1(n242), .A2(n218), .ZN(n69) );
  AND4_X1 U108 ( .A1(n142), .A2(n153), .A3(n140), .A4(n147), .ZN(n118) );
  AND4_X1 U109 ( .A1(n251), .A2(n253), .A3(n130), .A4(n135), .ZN(n110) );
  OAI21_X1 U110 ( .B1(n6), .B2(n231), .A(n246), .ZN(n70) );
  OAI21_X1 U111 ( .B1(n268), .B2(n233), .A(n262), .ZN(n71) );
  OR2_X1 U112 ( .A1(n69), .A2(n217), .ZN(n72) );
  NAND2_X1 U113 ( .A1(n72), .A2(n219), .ZN(n237) );
  OAI21_X1 U114 ( .B1(n245), .B2(n231), .A(n246), .ZN(n243) );
  OAI21_X1 U115 ( .B1(n268), .B2(n233), .A(n262), .ZN(n133) );
  AND2_X1 U116 ( .A1(net22671), .A2(net22672), .ZN(n73) );
  AND2_X1 U117 ( .A1(B[3]), .A2(A[3]), .ZN(n74) );
  NAND4_X1 U118 ( .A1(net22663), .A2(n55), .A3(net22640), .A4(n60), .ZN(n79)
         );
  NAND2_X1 U119 ( .A1(net37913), .A2(n16), .ZN(n80) );
  NAND2_X1 U120 ( .A1(n58), .A2(net37913), .ZN(net22661) );
  NOR2_X1 U121 ( .A1(n79), .A2(net22669), .ZN(net37985) );
  NAND2_X1 U122 ( .A1(n73), .A2(net38000), .ZN(n78) );
  NAND2_X1 U123 ( .A1(net22655), .A2(net22641), .ZN(n76) );
  NAND2_X1 U124 ( .A1(net22640), .A2(net22641), .ZN(n81) );
  NAND2_X1 U125 ( .A1(net22638), .A2(net22641), .ZN(net22656) );
  NAND2_X1 U126 ( .A1(n78), .A2(net37967), .ZN(net34666) );
  AOI21_X1 U127 ( .B1(n84), .B2(n85), .A(n86), .ZN(n83) );
  XNOR2_X1 U128 ( .A(n83), .B(net33637), .ZN(SUM[31]) );
  INV_X1 U129 ( .A(n87), .ZN(n86) );
  OAI21_X1 U130 ( .B1(n89), .B2(n88), .A(n90), .ZN(n84) );
  INV_X1 U131 ( .A(n91), .ZN(n88) );
  OAI21_X1 U132 ( .B1(net34521), .B2(n88), .A(n90), .ZN(net27463) );
  OR2_X1 U133 ( .A1(B[30]), .A2(A[30]), .ZN(n85) );
  NAND2_X1 U134 ( .A1(n87), .A2(n85), .ZN(net36853) );
  NAND2_X1 U135 ( .A1(B[30]), .A2(A[30]), .ZN(n87) );
  NAND2_X1 U136 ( .A1(B[29]), .A2(A[29]), .ZN(n90) );
  OR2_X1 U137 ( .A1(B[29]), .A2(A[29]), .ZN(n91) );
  NAND2_X1 U138 ( .A1(net34455), .A2(n94), .ZN(n92) );
  NAND2_X1 U139 ( .A1(B[28]), .A2(A[28]), .ZN(n93) );
  NAND2_X1 U140 ( .A1(n93), .A2(n94), .ZN(net22595) );
  OAI21_X1 U141 ( .B1(n23), .B2(net22599), .A(net34690), .ZN(net22589) );
  CLKBUF_X1 U142 ( .A(net22600), .Z(net34690) );
  NAND2_X1 U143 ( .A1(net22610), .A2(net22628), .ZN(net22631) );
  NAND2_X1 U144 ( .A1(net34666), .A2(net22628), .ZN(net34522) );
  OR2_X1 U145 ( .A1(B[28]), .A2(A[28]), .ZN(n94) );
  NAND2_X1 U146 ( .A1(n56), .A2(net37671), .ZN(n95) );
  AND2_X1 U147 ( .A1(n95), .A2(net37669), .ZN(net22657) );
  INV_X1 U148 ( .A(net37913), .ZN(net37670) );
  AND2_X1 U149 ( .A1(B[10]), .A2(A[10]), .ZN(n96) );
  XNOR2_X1 U150 ( .A(net27463), .B(net36853), .ZN(SUM[30]) );
  INV_X1 U151 ( .A(n118), .ZN(n233) );
  CLKBUF_X1 U152 ( .A(n140), .Z(n97) );
  CLKBUF_X1 U153 ( .A(n247), .Z(n99) );
  INV_X1 U154 ( .A(n110), .ZN(n231) );
  AND4_X1 U155 ( .A1(n228), .A2(n229), .A3(n214), .A4(n230), .ZN(n98) );
  AND4_X1 U156 ( .A1(n230), .A2(n229), .A3(n214), .A4(n228), .ZN(n126) );
  CLKBUF_X1 U157 ( .A(n225), .Z(n100) );
  CLKBUF_X1 U158 ( .A(A[14]), .Z(n101) );
  CLKBUF_X1 U159 ( .A(B[0]), .Z(n102) );
  OR2_X1 U160 ( .A1(A[11]), .A2(B[11]), .ZN(n251) );
  INV_X1 U161 ( .A(n158), .ZN(n103) );
  CLKBUF_X1 U162 ( .A(n165), .Z(n104) );
  AND2_X1 U163 ( .A1(B[2]), .A2(A[2]), .ZN(n105) );
  CLKBUF_X1 U164 ( .A(n131), .Z(n107) );
  OR2_X1 U165 ( .A1(B[9]), .A2(A[9]), .ZN(n130) );
  CLKBUF_X1 U166 ( .A(n151), .Z(n109) );
  CLKBUF_X1 U167 ( .A(n253), .Z(n111) );
  NAND2_X1 U168 ( .A1(net34522), .A2(n115), .ZN(n112) );
  AND2_X1 U169 ( .A1(n112), .A2(n113), .ZN(n184) );
  OR2_X1 U170 ( .A1(n114), .A2(n179), .ZN(n113) );
  INV_X1 U171 ( .A(n178), .ZN(n114) );
  AND2_X1 U172 ( .A1(net22610), .A2(n178), .ZN(n115) );
  CLKBUF_X1 U173 ( .A(n65), .Z(n116) );
  CLKBUF_X1 U174 ( .A(n134), .Z(n117) );
  CLKBUF_X1 U175 ( .A(n146), .Z(n119) );
  OAI211_X1 U176 ( .C1(n247), .C2(n248), .A(n249), .B(n250), .ZN(n120) );
  CLKBUF_X1 U177 ( .A(n202), .Z(n121) );
  AND2_X1 U178 ( .A1(net22688), .A2(n190), .ZN(n122) );
  XOR2_X1 U179 ( .A(n123), .B(n204), .Z(SUM[18]) );
  AND2_X1 U180 ( .A1(n195), .A2(n191), .ZN(n123) );
  XOR2_X1 U181 ( .A(n124), .B(n205), .Z(SUM[17]) );
  AND2_X1 U182 ( .A1(n200), .A2(n193), .ZN(n124) );
  XOR2_X1 U183 ( .A(n255), .B(n125), .Z(SUM[11]) );
  AND2_X1 U184 ( .A1(n250), .A2(n116), .ZN(n125) );
  OR2_X1 U185 ( .A1(B[10]), .A2(A[10]), .ZN(n253) );
  NAND2_X1 U186 ( .A1(n273), .A2(n274), .ZN(n269) );
  INV_X1 U187 ( .A(n5), .ZN(n152) );
  INV_X1 U188 ( .A(n121), .ZN(n167) );
  NAND2_X1 U189 ( .A1(n180), .A2(n174), .ZN(n181) );
  XNOR2_X1 U190 ( .A(net22661), .B(net22658), .ZN(SUM[21]) );
  XNOR2_X1 U191 ( .A(n185), .B(n184), .ZN(SUM[26]) );
  NAND2_X1 U192 ( .A1(n172), .A2(n175), .ZN(n185) );
  XNOR2_X1 U193 ( .A(net22655), .B(net22656), .ZN(SUM[22]) );
  NAND2_X1 U194 ( .A1(n178), .A2(n179), .ZN(n187) );
  NAND2_X1 U195 ( .A1(n8), .A2(n192), .ZN(n207) );
  XNOR2_X1 U196 ( .A(n258), .B(n257), .ZN(SUM[10]) );
  XNOR2_X1 U197 ( .A(n241), .B(n240), .ZN(SUM[13]) );
  XNOR2_X1 U198 ( .A(n234), .B(n235), .ZN(SUM[15]) );
  XNOR2_X1 U199 ( .A(n239), .B(n237), .ZN(SUM[14]) );
  XNOR2_X1 U200 ( .A(n244), .B(n70), .ZN(SUM[12]) );
  OAI21_X1 U201 ( .B1(n144), .B2(n145), .A(n119), .ZN(n141) );
  OAI21_X1 U202 ( .B1(n9), .B2(n198), .A(n200), .ZN(n204) );
  OAI21_X1 U203 ( .B1(n259), .B2(n260), .A(n107), .ZN(n257) );
  NOR2_X1 U204 ( .A1(n169), .A2(n170), .ZN(net22600) );
  XNOR2_X1 U205 ( .A(n163), .B(n160), .ZN(SUM[2]) );
  XNOR2_X1 U206 ( .A(n155), .B(n156), .ZN(SUM[3]) );
  XNOR2_X1 U207 ( .A(n201), .B(n167), .ZN(SUM[1]) );
  AOI21_X1 U208 ( .B1(n214), .B2(n237), .A(n216), .ZN(n234) );
  OAI21_X1 U209 ( .B1(n217), .B2(n218), .A(n219), .ZN(n215) );
  XNOR2_X1 U210 ( .A(net22589), .B(net22595), .ZN(SUM[28]) );
  NOR2_X1 U211 ( .A1(n212), .A2(n236), .ZN(n235) );
  OAI21_X1 U212 ( .B1(n17), .B2(n183), .A(n172), .ZN(n182) );
  NAND2_X1 U213 ( .A1(n243), .A2(n228), .ZN(n242) );
  INV_X1 U214 ( .A(n210), .ZN(n209) );
  XNOR2_X1 U215 ( .A(n132), .B(n71), .ZN(SUM[8]) );
  NAND2_X1 U216 ( .A1(n206), .A2(n8), .ZN(n205) );
  NAND2_X1 U217 ( .A1(n204), .A2(n191), .ZN(n203) );
  NAND2_X1 U218 ( .A1(n252), .A2(n256), .ZN(n255) );
  NAND2_X1 U219 ( .A1(n257), .A2(n253), .ZN(n256) );
  NAND2_X1 U220 ( .A1(n164), .A2(n104), .ZN(n160) );
  NAND2_X1 U221 ( .A1(n166), .A2(n167), .ZN(n164) );
  XOR2_X1 U222 ( .A(n127), .B(n129), .Z(SUM[9]) );
  AND2_X1 U223 ( .A1(n67), .A2(n107), .ZN(n127) );
  XNOR2_X1 U224 ( .A(n149), .B(n148), .ZN(SUM[5]) );
  XNOR2_X1 U225 ( .A(n154), .B(n152), .ZN(SUM[4]) );
  XNOR2_X1 U226 ( .A(n136), .B(n137), .ZN(SUM[7]) );
  NAND2_X1 U227 ( .A1(n68), .A2(n143), .ZN(n136) );
  NAND2_X1 U228 ( .A1(n138), .A2(n139), .ZN(n137) );
  NAND2_X1 U229 ( .A1(n97), .A2(n141), .ZN(n138) );
  XOR2_X1 U230 ( .A(n128), .B(n141), .Z(SUM[6]) );
  AND2_X1 U231 ( .A1(n97), .A2(n139), .ZN(n128) );
  AOI21_X1 U232 ( .B1(n266), .B2(n142), .A(n267), .ZN(n263) );
  NAND2_X1 U233 ( .A1(n103), .A2(n159), .ZN(n163) );
  NAND2_X1 U234 ( .A1(n218), .A2(n228), .ZN(n244) );
  NAND2_X1 U235 ( .A1(n219), .A2(n229), .ZN(n241) );
  NAND2_X1 U236 ( .A1(n166), .A2(n104), .ZN(n201) );
  NAND2_X1 U237 ( .A1(n252), .A2(n111), .ZN(n258) );
  NAND2_X1 U238 ( .A1(n238), .A2(n214), .ZN(n239) );
  OAI21_X1 U239 ( .B1(n157), .B2(n158), .A(n159), .ZN(n156) );
  NOR2_X1 U240 ( .A1(n188), .A2(n189), .ZN(net22672) );
  NAND2_X1 U241 ( .A1(n192), .A2(n193), .ZN(n188) );
  NAND2_X1 U242 ( .A1(n190), .A2(n191), .ZN(n189) );
  AOI21_X1 U243 ( .B1(n194), .B2(n195), .A(n196), .ZN(net22680) );
  NAND2_X1 U244 ( .A1(n197), .A2(n191), .ZN(n194) );
  OAI21_X1 U245 ( .B1(n198), .B2(n199), .A(n200), .ZN(n197) );
  AOI21_X1 U246 ( .B1(n171), .B2(n172), .A(n173), .ZN(n170) );
  NAND2_X1 U247 ( .A1(n175), .A2(n176), .ZN(n171) );
  OAI21_X1 U248 ( .B1(n177), .B2(net22610), .A(n178), .ZN(n176) );
  OAI211_X1 U249 ( .C1(n99), .C2(n64), .A(n106), .B(n250), .ZN(n224) );
  NAND2_X1 U250 ( .A1(n65), .A2(n96), .ZN(n249) );
  NAND2_X1 U251 ( .A1(n254), .A2(n253), .ZN(n247) );
  INV_X1 U252 ( .A(n102), .ZN(n273) );
  NAND2_X1 U253 ( .A1(n108), .A2(n153), .ZN(n150) );
  OR2_X1 U254 ( .A1(B[7]), .A2(A[7]), .ZN(n142) );
  NAND2_X1 U255 ( .A1(B[26]), .A2(A[26]), .ZN(n172) );
  NAND2_X1 U256 ( .A1(B[25]), .A2(A[25]), .ZN(n178) );
  NAND2_X1 U257 ( .A1(B[16]), .A2(A[16]), .ZN(n199) );
  NAND2_X1 U258 ( .A1(B[24]), .A2(A[24]), .ZN(net22610) );
  OR2_X1 U259 ( .A1(B[18]), .A2(A[18]), .ZN(n191) );
  OR2_X1 U260 ( .A1(B[25]), .A2(A[25]), .ZN(n179) );
  OR2_X1 U261 ( .A1(B[27]), .A2(A[27]), .ZN(n174) );
  NAND2_X1 U262 ( .A1(B[27]), .A2(A[27]), .ZN(n180) );
  NAND2_X1 U263 ( .A1(B[23]), .A2(n62), .ZN(net22647) );
  OR2_X1 U264 ( .A1(B[26]), .A2(A[26]), .ZN(n175) );
  OR2_X1 U265 ( .A1(A[8]), .A2(B[8]), .ZN(n135) );
  OR2_X1 U266 ( .A1(A[17]), .A2(B[17]), .ZN(n193) );
  OR2_X1 U267 ( .A1(B[6]), .A2(A[6]), .ZN(n140) );
  OR2_X1 U268 ( .A1(B[19]), .A2(A[19]), .ZN(n190) );
  OR2_X1 U269 ( .A1(B[16]), .A2(A[16]), .ZN(n192) );
  OR2_X1 U270 ( .A1(B[1]), .A2(A[1]), .ZN(n166) );
  OR2_X1 U271 ( .A1(B[13]), .A2(A[13]), .ZN(n229) );
  OR2_X1 U272 ( .A1(B[4]), .A2(A[4]), .ZN(n153) );
  OR2_X1 U273 ( .A1(B[3]), .A2(A[3]), .ZN(n161) );
  XOR2_X1 U274 ( .A(B[31]), .B(A[31]), .Z(net33637) );
  OR2_X1 U275 ( .A1(B[15]), .A2(A[15]), .ZN(n230) );
  NOR2_X1 U276 ( .A1(n226), .A2(n227), .ZN(n220) );
  NAND2_X1 U277 ( .A1(n131), .A2(n134), .ZN(n254) );
  NAND2_X1 U278 ( .A1(n261), .A2(n117), .ZN(n129) );
  NAND2_X1 U279 ( .A1(B[19]), .A2(A[19]), .ZN(net22688) );
  NAND2_X1 U280 ( .A1(n130), .A2(n251), .ZN(n248) );
  NAND2_X1 U281 ( .A1(n147), .A2(n119), .ZN(n149) );
  NAND4_X1 U282 ( .A1(n142), .A2(n147), .A3(n140), .A4(n265), .ZN(n264) );
  NAND2_X1 U283 ( .A1(B[22]), .A2(n63), .ZN(net22638) );
  NAND2_X1 U284 ( .A1(A[17]), .A2(B[17]), .ZN(n200) );
  NAND2_X1 U285 ( .A1(n202), .A2(n165), .ZN(n272) );
  OAI21_X1 U286 ( .B1(n211), .B2(n212), .A(n213), .ZN(n210) );
  AOI21_X1 U287 ( .B1(n214), .B2(n215), .A(n216), .ZN(n211) );
  NAND2_X1 U288 ( .A1(B[6]), .A2(A[6]), .ZN(n139) );
  NAND2_X1 U289 ( .A1(B[14]), .A2(n101), .ZN(n238) );
  NAND2_X1 U290 ( .A1(n117), .A2(n135), .ZN(n132) );
  NAND2_X1 U291 ( .A1(n71), .A2(n135), .ZN(n261) );
  XNOR2_X1 U292 ( .A(n186), .B(n187), .ZN(SUM[25]) );
  NAND2_X1 U293 ( .A1(n271), .A2(n270), .ZN(n232) );
  NAND2_X1 U294 ( .A1(B[18]), .A2(A[18]), .ZN(n195) );
  NAND2_X1 U295 ( .A1(B[8]), .A2(A[8]), .ZN(n134) );
  XNOR2_X1 U296 ( .A(n2), .B(net22666), .ZN(SUM[20]) );
  NAND2_X1 U297 ( .A1(B[0]), .A2(A[0]), .ZN(n202) );
  INV_X1 U298 ( .A(A[0]), .ZN(n274) );
  NAND2_X1 U299 ( .A1(B[12]), .A2(A[12]), .ZN(n218) );
  NOR2_X1 U300 ( .A1(n221), .A2(n220), .ZN(n208) );
  NAND2_X1 U301 ( .A1(B[5]), .A2(A[5]), .ZN(n146) );
  NAND2_X1 U302 ( .A1(B[9]), .A2(A[9]), .ZN(n131) );
  NAND2_X1 U303 ( .A1(n109), .A2(n153), .ZN(n154) );
  NAND2_X1 U304 ( .A1(n150), .A2(n109), .ZN(n148) );
  NAND2_X1 U305 ( .A1(n208), .A2(n209), .ZN(net22671) );
  NAND2_X1 U306 ( .A1(n263), .A2(n264), .ZN(n225) );
  NAND2_X1 U307 ( .A1(n146), .A2(n151), .ZN(n265) );
  NAND2_X1 U308 ( .A1(B[4]), .A2(A[4]), .ZN(n151) );
  NAND2_X1 U309 ( .A1(n232), .A2(n118), .ZN(n226) );
  XNOR2_X1 U310 ( .A(net34472), .B(n207), .ZN(SUM[16]) );
  NAND2_X1 U311 ( .A1(n23), .A2(net22610), .ZN(n186) );
  NAND2_X1 U312 ( .A1(net34472), .A2(n192), .ZN(n206) );
  NAND2_X1 U313 ( .A1(n110), .A2(n126), .ZN(n227) );
  NAND2_X1 U314 ( .A1(B[15]), .A2(A[15]), .ZN(n213) );
  NAND2_X1 U315 ( .A1(n66), .A2(n162), .ZN(n155) );
  AOI21_X1 U316 ( .B1(n161), .B2(n105), .A(n74), .ZN(n270) );
  NAND4_X1 U317 ( .A1(n272), .A2(n166), .A3(n168), .A4(n161), .ZN(n271) );
  NAND2_X1 U318 ( .A1(B[13]), .A2(A[13]), .ZN(n219) );
  NAND2_X1 U319 ( .A1(B[11]), .A2(A[11]), .ZN(n250) );
  NAND2_X1 U320 ( .A1(A[7]), .A2(B[7]), .ZN(n143) );
  NAND2_X1 U321 ( .A1(B[1]), .A2(A[1]), .ZN(n165) );
  INV_X1 U322 ( .A(n147), .ZN(n145) );
  INV_X1 U323 ( .A(n148), .ZN(n144) );
  INV_X1 U324 ( .A(n160), .ZN(n157) );
  INV_X1 U325 ( .A(n174), .ZN(n173) );
  INV_X1 U326 ( .A(n179), .ZN(n177) );
  INV_X1 U327 ( .A(n180), .ZN(n169) );
  NAND3_X1 U328 ( .A1(n175), .A2(n174), .A3(n179), .ZN(net22599) );
  XNOR2_X1 U329 ( .A(n182), .B(n181), .ZN(SUM[27]) );
  INV_X1 U330 ( .A(n175), .ZN(n183) );
  XNOR2_X1 U331 ( .A(net22631), .B(net28033), .ZN(SUM[24]) );
  INV_X1 U332 ( .A(n190), .ZN(n196) );
  INV_X1 U333 ( .A(n193), .ZN(n198) );
  NAND2_X1 U334 ( .A1(n223), .A2(n222), .ZN(n221) );
  NAND2_X1 U335 ( .A1(n120), .A2(n98), .ZN(n223) );
  NAND3_X1 U336 ( .A1(n225), .A2(n110), .A3(n98), .ZN(n222) );
  INV_X1 U337 ( .A(n213), .ZN(n236) );
  INV_X1 U338 ( .A(n230), .ZN(n212) );
  INV_X1 U339 ( .A(n238), .ZN(n216) );
  INV_X1 U340 ( .A(n229), .ZN(n217) );
  INV_X1 U341 ( .A(n224), .ZN(n246) );
  INV_X1 U342 ( .A(n133), .ZN(n245) );
  INV_X1 U343 ( .A(n129), .ZN(n260) );
  INV_X1 U344 ( .A(n100), .ZN(n262) );
  INV_X1 U345 ( .A(n143), .ZN(n267) );
  INV_X1 U346 ( .A(n139), .ZN(n266) );
  INV_X1 U347 ( .A(n168), .ZN(n158) );
  INV_X1 U348 ( .A(n108), .ZN(n268) );
  INV_X1 U349 ( .A(n67), .ZN(n259) );
endmodule


module ALU_DATA_W32_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331;

  AND2_X1 U1 ( .A1(n106), .A2(n105), .ZN(n103) );
  AND2_X1 U2 ( .A1(n25), .A2(n26), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n269), .A2(n118), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n269), .A2(n118), .ZN(n129) );
  AND3_X1 U5 ( .A1(n3), .A2(n4), .A3(n5), .ZN(n18) );
  AND2_X1 U6 ( .A1(n22), .A2(n23), .ZN(n3) );
  OR2_X1 U7 ( .A1(n19), .A2(n21), .ZN(n4) );
  OR2_X1 U8 ( .A1(n19), .A2(n20), .ZN(n5) );
  NAND2_X1 U9 ( .A1(n243), .A2(n91), .ZN(n6) );
  AND2_X1 U10 ( .A1(n162), .A2(n163), .ZN(n7) );
  AND2_X1 U11 ( .A1(n8), .A2(n9), .ZN(n22) );
  OR2_X1 U12 ( .A1(n11), .A2(n30), .ZN(n8) );
  OR2_X1 U13 ( .A1(n11), .A2(n29), .ZN(n9) );
  AND2_X1 U14 ( .A1(n243), .A2(n91), .ZN(n10) );
  NAND2_X1 U15 ( .A1(n329), .A2(n26), .ZN(n11) );
  NAND2_X1 U16 ( .A1(n162), .A2(n163), .ZN(n19) );
  NAND2_X1 U17 ( .A1(n163), .A2(n325), .ZN(n172) );
  NAND2_X1 U18 ( .A1(n99), .A2(n100), .ZN(n98) );
  NAND2_X1 U19 ( .A1(n103), .A2(n104), .ZN(n99) );
  NAND2_X1 U20 ( .A1(n53), .A2(n54), .ZN(n52) );
  NAND2_X1 U21 ( .A1(n57), .A2(n58), .ZN(n53) );
  AOI21_X1 U22 ( .B1(n81), .B2(n82), .A(n83), .ZN(n69) );
  NOR2_X1 U23 ( .A1(n97), .A2(n98), .ZN(n82) );
  AOI21_X1 U24 ( .B1(n34), .B2(n35), .A(n36), .ZN(n17) );
  NOR2_X1 U25 ( .A1(n51), .A2(n52), .ZN(n35) );
  OAI21_X1 U26 ( .B1(n69), .B2(n68), .A(n70), .ZN(n34) );
  OAI21_X1 U27 ( .B1(n220), .B2(n219), .A(n221), .ZN(n187) );
  NAND4_X1 U28 ( .A1(n291), .A2(n292), .A3(n293), .A4(n294), .ZN(n219) );
  NOR3_X1 U29 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n221) );
  AOI21_X1 U30 ( .B1(n233), .B2(n234), .A(n235), .ZN(n220) );
  NOR2_X1 U31 ( .A1(n2), .A2(n130), .ZN(n266) );
  NOR2_X1 U32 ( .A1(n142), .A2(n73), .ZN(n291) );
  NOR2_X1 U33 ( .A1(n67), .A2(n45), .ZN(n204) );
  NOR2_X1 U34 ( .A1(n111), .A2(n6), .ZN(n249) );
  OAI21_X1 U35 ( .B1(n167), .B2(n166), .A(n168), .ZN(n165) );
  AOI21_X1 U36 ( .B1(n187), .B2(n188), .A(n189), .ZN(n167) );
  NAND2_X1 U37 ( .A1(n264), .A2(n265), .ZN(n233) );
  AOI21_X1 U38 ( .B1(n267), .B2(n266), .A(n268), .ZN(n265) );
  NOR2_X1 U39 ( .A1(n281), .A2(n282), .ZN(n264) );
  NOR2_X1 U40 ( .A1(n272), .A2(n273), .ZN(n267) );
  NAND2_X1 U41 ( .A1(n225), .A2(n80), .ZN(n73) );
  NOR2_X1 U42 ( .A1(n71), .A2(n72), .ZN(n70) );
  NAND4_X1 U43 ( .A1(n61), .A2(n79), .A3(n62), .A4(n80), .ZN(n71) );
  OAI22_X1 U44 ( .A1(n73), .A2(n74), .B1(n73), .B2(n75), .ZN(n72) );
  NOR3_X1 U45 ( .A1(n45), .A2(n194), .A3(n195), .ZN(n193) );
  NOR3_X1 U46 ( .A1(n6), .A2(n239), .A3(n240), .ZN(n238) );
  NOR3_X1 U47 ( .A1(n169), .A2(n170), .A3(n171), .ZN(n168) );
  NOR2_X1 U48 ( .A1(n172), .A2(n174), .ZN(n170) );
  NOR2_X1 U49 ( .A1(n172), .A2(n164), .ZN(n171) );
  NAND2_X1 U50 ( .A1(n198), .A2(n44), .ZN(n45) );
  NOR2_X1 U51 ( .A1(n28), .A2(n326), .ZN(n163) );
  NAND2_X1 U52 ( .A1(n33), .A2(n186), .ZN(n326) );
  NAND2_X1 U53 ( .A1(n243), .A2(n91), .ZN(n92) );
  NOR2_X1 U54 ( .A1(n142), .A2(n73), .ZN(n138) );
  OAI21_X1 U55 ( .B1(n129), .B2(n283), .A(n255), .ZN(n282) );
  OAI21_X1 U56 ( .B1(n73), .B2(n229), .A(n210), .ZN(n222) );
  NAND2_X1 U57 ( .A1(n207), .A2(n62), .ZN(n58) );
  NOR2_X1 U58 ( .A1(n73), .A2(n77), .ZN(n223) );
  NAND2_X1 U59 ( .A1(n199), .A2(n43), .ZN(n159) );
  NOR2_X1 U60 ( .A1(n2), .A2(n124), .ZN(n281) );
  NOR2_X1 U61 ( .A1(n181), .A2(n182), .ZN(n175) );
  NOR2_X1 U62 ( .A1(n11), .A2(n184), .ZN(n181) );
  NOR2_X1 U63 ( .A1(n11), .A2(n32), .ZN(n182) );
  NAND2_X1 U64 ( .A1(n244), .A2(n90), .ZN(n146) );
  NOR2_X1 U65 ( .A1(n45), .A2(n56), .ZN(n196) );
  NAND2_X1 U66 ( .A1(n252), .A2(n106), .ZN(n104) );
  NOR2_X1 U67 ( .A1(n92), .A2(n102), .ZN(n241) );
  NAND2_X1 U68 ( .A1(n279), .A2(n134), .ZN(n130) );
  AND2_X1 U69 ( .A1(n164), .A2(n32), .ZN(n162) );
  AND2_X1 U70 ( .A1(n20), .A2(n29), .ZN(n325) );
  NOR2_X1 U71 ( .A1(n276), .A2(n277), .ZN(n272) );
  NOR2_X1 U72 ( .A1(A[0]), .A2(n278), .ZN(n276) );
  NAND2_X1 U73 ( .A1(n232), .A2(n78), .ZN(n142) );
  NAND2_X1 U74 ( .A1(n174), .A2(n21), .ZN(n155) );
  NAND2_X1 U75 ( .A1(n157), .A2(n199), .ZN(n316) );
  NAND2_X1 U76 ( .A1(n195), .A2(n50), .ZN(n67) );
  NAND2_X1 U77 ( .A1(n156), .A2(n157), .ZN(n150) );
  NAND2_X1 U78 ( .A1(n158), .A2(n159), .ZN(n156) );
  NOR2_X1 U79 ( .A1(n121), .A2(n122), .ZN(n120) );
  NOR2_X1 U80 ( .A1(n2), .A2(n130), .ZN(n119) );
  NAND2_X1 U81 ( .A1(n123), .A2(n124), .ZN(n122) );
  NAND2_X1 U82 ( .A1(n240), .A2(n96), .ZN(n111) );
  NOR2_X1 U83 ( .A1(n150), .A2(n151), .ZN(n149) );
  OAI21_X1 U84 ( .B1(n152), .B2(n153), .A(n154), .ZN(n151) );
  NAND2_X1 U85 ( .A1(n41), .A2(n43), .ZN(n153) );
  NOR2_X1 U86 ( .A1(n115), .A2(n116), .ZN(n114) );
  NAND2_X1 U87 ( .A1(n106), .A2(n118), .ZN(n115) );
  NAND2_X1 U88 ( .A1(n105), .A2(n117), .ZN(n116) );
  NOR2_X1 U89 ( .A1(n39), .A2(n40), .ZN(n38) );
  NAND2_X1 U90 ( .A1(n41), .A2(n42), .ZN(n40) );
  NAND2_X1 U91 ( .A1(n43), .A2(n44), .ZN(n39) );
  NOR2_X1 U92 ( .A1(n132), .A2(n131), .ZN(n112) );
  NOR2_X1 U93 ( .A1(n129), .A2(n135), .ZN(n131) );
  NOR3_X1 U94 ( .A1(n129), .A2(n133), .A3(n134), .ZN(n132) );
  NOR2_X1 U95 ( .A1(n86), .A2(n87), .ZN(n85) );
  NAND2_X1 U96 ( .A1(n90), .A2(n91), .ZN(n86) );
  NAND2_X1 U97 ( .A1(n88), .A2(n89), .ZN(n87) );
  NAND2_X1 U98 ( .A1(n274), .A2(n135), .ZN(n273) );
  NAND2_X1 U99 ( .A1(n206), .A2(n58), .ZN(n205) );
  NAND2_X1 U100 ( .A1(n251), .A2(n104), .ZN(n250) );
  NAND2_X1 U101 ( .A1(n301), .A2(n146), .ZN(n292) );
  NOR2_X1 U102 ( .A1(n247), .A2(n248), .ZN(n234) );
  OAI211_X1 U103 ( .C1(n117), .C2(n260), .A(n105), .B(n93), .ZN(n247) );
  NAND2_X1 U104 ( .A1(n249), .A2(n250), .ZN(n248) );
  NAND2_X1 U105 ( .A1(n255), .A2(n252), .ZN(n260) );
  NOR2_X1 U106 ( .A1(n202), .A2(n203), .ZN(n188) );
  OAI211_X1 U107 ( .C1(n79), .C2(n215), .A(n61), .B(n46), .ZN(n202) );
  NAND2_X1 U108 ( .A1(n204), .A2(n205), .ZN(n203) );
  NAND2_X1 U109 ( .A1(n210), .A2(n207), .ZN(n215) );
  NAND2_X1 U110 ( .A1(n191), .A2(n190), .ZN(n189) );
  NOR2_X1 U111 ( .A1(n196), .A2(n197), .ZN(n190) );
  NOR2_X1 U112 ( .A1(n193), .A2(n192), .ZN(n191) );
  NAND2_X1 U113 ( .A1(n237), .A2(n236), .ZN(n235) );
  NOR2_X1 U114 ( .A1(n241), .A2(n242), .ZN(n236) );
  NOR2_X1 U115 ( .A1(n238), .A2(n143), .ZN(n237) );
  NAND2_X1 U116 ( .A1(n145), .A2(n146), .ZN(n136) );
  NAND2_X1 U117 ( .A1(n47), .A2(n48), .ZN(n37) );
  NOR2_X1 U118 ( .A1(n49), .A2(n50), .ZN(n47) );
  NAND2_X1 U119 ( .A1(n94), .A2(n10), .ZN(n84) );
  NOR2_X1 U120 ( .A1(n95), .A2(n96), .ZN(n94) );
  OR2_X1 U121 ( .A1(n45), .A2(n46), .ZN(n12) );
  OR2_X1 U122 ( .A1(n92), .A2(n93), .ZN(n13) );
  AND2_X1 U123 ( .A1(n312), .A2(n313), .ZN(n311) );
  NOR2_X1 U124 ( .A1(n314), .A2(n161), .ZN(n313) );
  AOI21_X1 U125 ( .B1(n318), .B2(n159), .A(n155), .ZN(n312) );
  NOR2_X1 U126 ( .A1(n42), .A2(n316), .ZN(n314) );
  INV_X1 U127 ( .A(A[18]), .ZN(n226) );
  XNOR2_X1 U128 ( .A(B[31]), .B(A[31]), .ZN(n26) );
  NAND2_X1 U129 ( .A1(B[24]), .A2(n324), .ZN(n199) );
  INV_X1 U130 ( .A(A[24]), .ZN(n324) );
  NAND2_X1 U131 ( .A1(B[25]), .A2(n323), .ZN(n157) );
  INV_X1 U132 ( .A(A[25]), .ZN(n323) );
  INV_X1 U133 ( .A(B[19]), .ZN(n217) );
  NAND2_X1 U134 ( .A1(B[26]), .A2(n320), .ZN(n174) );
  INV_X1 U135 ( .A(A[26]), .ZN(n320) );
  NAND2_X1 U136 ( .A1(B[19]), .A2(n230), .ZN(n210) );
  NAND2_X1 U137 ( .A1(n329), .A2(n26), .ZN(n28) );
  NAND2_X1 U138 ( .A1(B[27]), .A2(n173), .ZN(n164) );
  INV_X1 U139 ( .A(A[27]), .ZN(n173) );
  NAND2_X1 U140 ( .A1(B[20]), .A2(n214), .ZN(n195) );
  INV_X1 U141 ( .A(A[20]), .ZN(n214) );
  NAND2_X1 U142 ( .A1(A[24]), .A2(n321), .ZN(n43) );
  INV_X1 U143 ( .A(B[24]), .ZN(n321) );
  INV_X1 U144 ( .A(A[3]), .ZN(n288) );
  INV_X1 U145 ( .A(B[21]), .ZN(n216) );
  NAND2_X1 U146 ( .A1(B[23]), .A2(n200), .ZN(n152) );
  INV_X1 U147 ( .A(A[23]), .ZN(n200) );
  NAND2_X1 U148 ( .A1(B[21]), .A2(n201), .ZN(n56) );
  NAND2_X1 U149 ( .A1(B[29]), .A2(n183), .ZN(n32) );
  NAND2_X1 U150 ( .A1(B[22]), .A2(n212), .ZN(n198) );
  NAND2_X1 U151 ( .A1(B[16]), .A2(n307), .ZN(n225) );
  INV_X1 U152 ( .A(A[16]), .ZN(n307) );
  INV_X1 U153 ( .A(A[17]), .ZN(n227) );
  INV_X1 U154 ( .A(B[22]), .ZN(n211) );
  NAND2_X1 U155 ( .A1(B[28]), .A2(n327), .ZN(n186) );
  NAND2_X1 U156 ( .A1(A[23]), .A2(n317), .ZN(n42) );
  INV_X1 U157 ( .A(B[23]), .ZN(n317) );
  NAND2_X1 U158 ( .A1(A[26]), .A2(n319), .ZN(n21) );
  INV_X1 U159 ( .A(B[26]), .ZN(n319) );
  NAND2_X1 U160 ( .A1(A[20]), .A2(n213), .ZN(n50) );
  INV_X1 U161 ( .A(B[20]), .ZN(n213) );
  NAND2_X1 U162 ( .A1(A[25]), .A2(n315), .ZN(n41) );
  INV_X1 U163 ( .A(B[25]), .ZN(n315) );
  NAND2_X1 U164 ( .A1(A[17]), .A2(n218), .ZN(n79) );
  INV_X1 U165 ( .A(B[28]), .ZN(n328) );
  NAND2_X1 U166 ( .A1(A[27]), .A2(n331), .ZN(n20) );
  INV_X1 U167 ( .A(B[27]), .ZN(n331) );
  NAND2_X1 U168 ( .A1(A[16]), .A2(n306), .ZN(n80) );
  INV_X1 U169 ( .A(B[16]), .ZN(n306) );
  NAND2_X1 U170 ( .A1(A[18]), .A2(n208), .ZN(n62) );
  INV_X1 U171 ( .A(B[29]), .ZN(n330) );
  NOR2_X1 U172 ( .A1(n126), .A2(n127), .ZN(n121) );
  INV_X1 U173 ( .A(A[0]), .ZN(n128) );
  INV_X1 U174 ( .A(A[31]), .ZN(n180) );
  NOR2_X1 U175 ( .A1(B[30]), .A2(n27), .ZN(n25) );
  INV_X1 U176 ( .A(A[30]), .ZN(n27) );
  NOR2_X1 U177 ( .A1(A[30]), .A2(n179), .ZN(n178) );
  INV_X1 U178 ( .A(B[30]), .ZN(n179) );
  NAND2_X1 U179 ( .A1(A[3]), .A2(n286), .ZN(n135) );
  NOR2_X1 U180 ( .A1(n24), .A2(n1), .ZN(n23) );
  NOR2_X1 U181 ( .A1(B[31]), .A2(n180), .ZN(n24) );
  AND2_X1 U182 ( .A1(n14), .A2(n177), .ZN(n176) );
  NAND2_X1 U183 ( .A1(B[31]), .A2(n180), .ZN(n14) );
  OAI21_X1 U184 ( .B1(n17), .B2(n16), .A(n18), .ZN(n15) );
  NAND2_X1 U185 ( .A1(A[19]), .A2(n217), .ZN(n61) );
  INV_X1 U186 ( .A(A[19]), .ZN(n230) );
  INV_X1 U187 ( .A(A[29]), .ZN(n183) );
  NAND2_X1 U188 ( .A1(A[29]), .A2(n330), .ZN(n29) );
  NAND2_X1 U189 ( .A1(A[22]), .A2(n211), .ZN(n44) );
  INV_X1 U190 ( .A(A[22]), .ZN(n212) );
  INV_X1 U191 ( .A(B[6]), .ZN(n253) );
  NAND2_X1 U192 ( .A1(B[6]), .A2(n270), .ZN(n252) );
  NAND2_X1 U193 ( .A1(A[28]), .A2(n328), .ZN(n33) );
  INV_X1 U194 ( .A(A[28]), .ZN(n327) );
  NAND2_X1 U195 ( .A1(A[21]), .A2(n216), .ZN(n46) );
  INV_X1 U196 ( .A(A[21]), .ZN(n201) );
  NAND2_X1 U197 ( .A1(B[17]), .A2(n227), .ZN(n66) );
  INV_X1 U198 ( .A(B[17]), .ZN(n218) );
  NAND2_X1 U199 ( .A1(A[7]), .A2(n262), .ZN(n105) );
  INV_X1 U200 ( .A(A[7]), .ZN(n284) );
  NAND2_X1 U201 ( .A1(A[13]), .A2(n296), .ZN(n88) );
  INV_X1 U202 ( .A(A[13]), .ZN(n304) );
  NAND2_X1 U203 ( .A1(A[6]), .A2(n253), .ZN(n106) );
  INV_X1 U204 ( .A(A[6]), .ZN(n270) );
  NAND2_X1 U205 ( .A1(A[2]), .A2(n280), .ZN(n134) );
  INV_X1 U206 ( .A(A[2]), .ZN(n287) );
  NAND2_X1 U207 ( .A1(A[15]), .A2(n297), .ZN(n75) );
  INV_X1 U208 ( .A(A[15]), .ZN(n228) );
  NAND2_X1 U209 ( .A1(A[5]), .A2(n263), .ZN(n117) );
  INV_X1 U210 ( .A(A[5]), .ZN(n271) );
  NAND2_X1 U211 ( .A1(A[4]), .A2(n289), .ZN(n118) );
  INV_X1 U212 ( .A(A[4]), .ZN(n290) );
  NAND2_X1 U213 ( .A1(A[8]), .A2(n258), .ZN(n96) );
  INV_X1 U214 ( .A(A[8]), .ZN(n259) );
  NAND2_X1 U215 ( .A1(A[12]), .A2(n302), .ZN(n90) );
  INV_X1 U216 ( .A(A[12]), .ZN(n305) );
  INV_X1 U217 ( .A(B[14]), .ZN(n308) );
  NAND2_X1 U218 ( .A1(B[14]), .A2(n309), .ZN(n232) );
  NAND2_X1 U219 ( .A1(A[11]), .A2(n300), .ZN(n89) );
  INV_X1 U220 ( .A(A[11]), .ZN(n245) );
  NAND2_X1 U221 ( .A1(A[9]), .A2(n261), .ZN(n93) );
  INV_X1 U222 ( .A(A[9]), .ZN(n246) );
  NAND2_X1 U223 ( .A1(A[10]), .A2(n256), .ZN(n91) );
  INV_X1 U224 ( .A(A[10]), .ZN(n257) );
  NAND2_X1 U225 ( .A1(A[14]), .A2(n308), .ZN(n78) );
  INV_X1 U226 ( .A(A[14]), .ZN(n309) );
  NAND2_X1 U227 ( .A1(A[1]), .A2(n275), .ZN(n274) );
  NOR2_X1 U228 ( .A1(A[1]), .A2(n275), .ZN(n277) );
  INV_X1 U229 ( .A(A[1]), .ZN(n125) );
  NAND2_X1 U230 ( .A1(B[2]), .A2(n287), .ZN(n279) );
  INV_X1 U231 ( .A(B[2]), .ZN(n280) );
  NAND2_X1 U232 ( .A1(B[18]), .A2(n226), .ZN(n207) );
  INV_X1 U233 ( .A(B[18]), .ZN(n208) );
  NAND2_X1 U234 ( .A1(B[8]), .A2(n259), .ZN(n240) );
  INV_X1 U235 ( .A(B[8]), .ZN(n258) );
  INV_X1 U236 ( .A(B[0]), .ZN(n278) );
  NOR2_X1 U237 ( .A1(B[0]), .A2(n128), .ZN(n126) );
  NAND2_X1 U238 ( .A1(B[12]), .A2(n305), .ZN(n244) );
  INV_X1 U239 ( .A(B[12]), .ZN(n302) );
  NAND2_X1 U240 ( .A1(B[5]), .A2(n271), .ZN(n110) );
  INV_X1 U241 ( .A(B[5]), .ZN(n263) );
  INV_X1 U242 ( .A(B[10]), .ZN(n256) );
  NAND2_X1 U243 ( .A1(B[10]), .A2(n257), .ZN(n243) );
  INV_X1 U244 ( .A(B[9]), .ZN(n261) );
  NAND2_X1 U245 ( .A1(B[9]), .A2(n246), .ZN(n102) );
  NAND2_X1 U246 ( .A1(B[3]), .A2(n288), .ZN(n124) );
  INV_X1 U247 ( .A(B[3]), .ZN(n286) );
  NAND2_X1 U248 ( .A1(B[4]), .A2(n290), .ZN(n269) );
  INV_X1 U249 ( .A(B[4]), .ZN(n289) );
  NAND2_X1 U250 ( .A1(B[15]), .A2(n228), .ZN(n77) );
  INV_X1 U251 ( .A(B[15]), .ZN(n297) );
  NAND2_X1 U252 ( .A1(B[13]), .A2(n304), .ZN(n298) );
  INV_X1 U253 ( .A(B[13]), .ZN(n296) );
  NAND2_X1 U254 ( .A1(B[11]), .A2(n245), .ZN(n141) );
  INV_X1 U255 ( .A(B[11]), .ZN(n300) );
  NAND2_X1 U256 ( .A1(B[7]), .A2(n284), .ZN(n255) );
  INV_X1 U257 ( .A(B[7]), .ZN(n262) );
  NOR2_X1 U258 ( .A1(B[1]), .A2(n125), .ZN(n127) );
  NAND2_X1 U259 ( .A1(B[1]), .A2(n125), .ZN(n123) );
  INV_X1 U260 ( .A(B[1]), .ZN(n275) );
  NAND2_X1 U261 ( .A1(GE), .A2(LE), .ZN(NE) );
  INV_X1 U262 ( .A(n15), .ZN(LE) );
  NAND2_X1 U263 ( .A1(n31), .A2(n32), .ZN(n30) );
  INV_X1 U264 ( .A(n33), .ZN(n31) );
  NAND3_X1 U265 ( .A1(n37), .A2(n12), .A3(n38), .ZN(n36) );
  NOR2_X1 U266 ( .A1(n55), .A2(n49), .ZN(n54) );
  INV_X1 U267 ( .A(n56), .ZN(n49) );
  NOR2_X1 U268 ( .A1(n59), .A2(n60), .ZN(n57) );
  INV_X1 U269 ( .A(n61), .ZN(n60) );
  INV_X1 U270 ( .A(n62), .ZN(n59) );
  NAND3_X1 U271 ( .A1(n48), .A2(n63), .A3(n64), .ZN(n51) );
  NAND3_X1 U272 ( .A1(n61), .A2(n62), .A3(n65), .ZN(n64) );
  INV_X1 U273 ( .A(n66), .ZN(n65) );
  INV_X1 U274 ( .A(n67), .ZN(n63) );
  INV_X1 U275 ( .A(n45), .ZN(n48) );
  NAND2_X1 U276 ( .A1(n76), .A2(n77), .ZN(n74) );
  INV_X1 U277 ( .A(n78), .ZN(n76) );
  NAND3_X1 U278 ( .A1(n84), .A2(n13), .A3(n85), .ZN(n83) );
  NOR2_X1 U279 ( .A1(n101), .A2(n95), .ZN(n100) );
  INV_X1 U280 ( .A(n102), .ZN(n95) );
  NAND3_X1 U281 ( .A1(n10), .A2(n107), .A3(n108), .ZN(n97) );
  NAND3_X1 U282 ( .A1(n105), .A2(n106), .A3(n109), .ZN(n108) );
  INV_X1 U283 ( .A(n110), .ZN(n109) );
  INV_X1 U284 ( .A(n111), .ZN(n107) );
  NAND3_X1 U285 ( .A1(n112), .A2(n113), .A3(n114), .ZN(n81) );
  NAND2_X1 U286 ( .A1(n119), .A2(n120), .ZN(n113) );
  INV_X1 U287 ( .A(n124), .ZN(n133) );
  NAND4_X1 U288 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(n68) );
  NAND3_X1 U289 ( .A1(n88), .A2(n90), .A3(n140), .ZN(n139) );
  INV_X1 U290 ( .A(n141), .ZN(n140) );
  NOR2_X1 U291 ( .A1(n143), .A2(n144), .ZN(n137) );
  INV_X1 U292 ( .A(n77), .ZN(n144) );
  NOR2_X1 U293 ( .A1(n147), .A2(n148), .ZN(n145) );
  INV_X1 U294 ( .A(n90), .ZN(n147) );
  NAND2_X1 U295 ( .A1(n7), .A2(n149), .ZN(n16) );
  INV_X1 U296 ( .A(n155), .ZN(n154) );
  NOR2_X1 U297 ( .A1(n160), .A2(n161), .ZN(n158) );
  INV_X1 U298 ( .A(n43), .ZN(n160) );
  INV_X1 U299 ( .A(n165), .ZN(GE) );
  NAND2_X1 U300 ( .A1(n175), .A2(n176), .ZN(n169) );
  NAND2_X1 U301 ( .A1(n178), .A2(n26), .ZN(n177) );
  NAND2_X1 U302 ( .A1(n185), .A2(n29), .ZN(n184) );
  INV_X1 U303 ( .A(n186), .ZN(n185) );
  INV_X1 U304 ( .A(n46), .ZN(n194) );
  NAND3_X1 U305 ( .A1(n198), .A2(n152), .A3(n199), .ZN(n197) );
  NOR2_X1 U306 ( .A1(n209), .A2(n55), .ZN(n206) );
  INV_X1 U307 ( .A(n210), .ZN(n55) );
  INV_X1 U308 ( .A(n207), .ZN(n209) );
  NAND3_X1 U309 ( .A1(n225), .A2(n66), .A3(n207), .ZN(n224) );
  NAND2_X1 U310 ( .A1(n231), .A2(n75), .ZN(n229) );
  INV_X1 U311 ( .A(n232), .ZN(n231) );
  INV_X1 U312 ( .A(n93), .ZN(n239) );
  NAND3_X1 U313 ( .A1(n243), .A2(n141), .A3(n244), .ZN(n242) );
  NOR2_X1 U314 ( .A1(n254), .A2(n101), .ZN(n251) );
  INV_X1 U315 ( .A(n255), .ZN(n101) );
  INV_X1 U316 ( .A(n252), .ZN(n254) );
  NAND3_X1 U317 ( .A1(n269), .A2(n110), .A3(n252), .ZN(n268) );
  NAND2_X1 U318 ( .A1(n285), .A2(n135), .ZN(n283) );
  INV_X1 U319 ( .A(n279), .ZN(n285) );
  NOR2_X1 U320 ( .A1(n295), .A2(n148), .ZN(n294) );
  INV_X1 U321 ( .A(n88), .ZN(n148) );
  INV_X1 U322 ( .A(n75), .ZN(n295) );
  NAND3_X1 U323 ( .A1(n298), .A2(n244), .A3(n299), .ZN(n293) );
  INV_X1 U324 ( .A(n89), .ZN(n299) );
  NOR2_X1 U325 ( .A1(n303), .A2(n143), .ZN(n301) );
  INV_X1 U326 ( .A(n298), .ZN(n143) );
  INV_X1 U327 ( .A(n244), .ZN(n303) );
  NAND2_X1 U328 ( .A1(n310), .A2(n311), .ZN(n166) );
  INV_X1 U329 ( .A(n41), .ZN(n161) );
  NOR2_X1 U330 ( .A1(n322), .A2(n192), .ZN(n318) );
  INV_X1 U331 ( .A(n157), .ZN(n192) );
  INV_X1 U332 ( .A(n199), .ZN(n322) );
  INV_X1 U333 ( .A(n172), .ZN(n310) );
  XNOR2_X1 U334 ( .A(B[30]), .B(A[30]), .ZN(n329) );
endmodule


module ALU_DATA_W32 ( .FUNC({\FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), A, 
        B, RES );
  input [31:0] A;
  input [31:0] B;
  output [31:0] RES;
  input \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N794, N795, N796, n121, n123, n124, n127, n136, n146, n148, n151,
         n157, n159, n162, n163, n170, n172, n175, n176, n183, n184, n186,
         n192, n195, n196, n197, n198, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n214, n217, n219, n220, n232, n239, n247,
         n253, n254, n258, n259, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n279, n285, n295, n302, n338, n339, n378, n401,
         n402, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n454, n465, n474, n480, n482, n483, n484, n485, n487,
         n488, n489, n496, n497, n506, n507, n508, n509, n512, n513, n520,
         n521, n522, n523, n527, n528, n540, n541, n542, n543, n544, n545,
         n547, n549, n550, net18425, net18431, net18434, net20020, net20024,
         net20044, net20047, net20105, net20206, net25112, net25113, net25114,
         net25116, net25130, net25131, net25132, net25136, net25137, net25138,
         net25143, net25146, net25150, net25169, net25231, net25236, net25237,
         net25238, net25366, net25429, net25442, net25443, net25448, net25464,
         net25484, net25499, net25502, net25503, net25523, net25527, net25577,
         net25583, net25596, net25629, net27095, net27083, net27081, net27105,
         net27103, net27101, net27113, net27127, net27125, net27123, net27121,
         net27143, net27141, net27137, net27133, net27131, net27161, net27159,
         net27155, net27151, net27149, net27175, net27167, net27165, net27179,
         net27177, net27185, net27183, net27181, net27191, net27189, net27187,
         net27203, net27201, net27195, net27193, net27209, net27207, net27205,
         net27408, net27525, net27527, net28242, net28241, net28422, net28421,
         net28420, net33169, net33190, net33647, net33654, net33657, net33684,
         net33829, net33834, net34232, net34298, net34297, net34351, net34566,
         net34616, net34655, net34836, net34835, net34866, net34869, net34889,
         net34906, net34986, net35006, net35005, net35004, net35616, net35624,
         net35631, net35986, net35985, net35981, net35893, net35871, net38433,
         net39040, net41315, net25121, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n19, n20, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n122, n125, n126, n128, n129, n130, n131, n132, n133, n134, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n147, n149,
         n150, n152, n153, n154, n155, n156, n158, n160, n161, n164, n165,
         n166, n167, n168, n169, n171, n173, n174, n177, n178, n179, n180,
         n181, n182, n185, n187, n188, n189, n190, n191, n193, n194, n199,
         n200, n201, n212, n213, n215, n216, n218, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n233, n234, n235, n236,
         n237, n238, n240, n241, n242, n243, n244, n245, n246, n248, n249,
         n250, n251, n252, n255, n256, n257, n260, n261, n262, n273, n274,
         n275, n276, n277, n278, n280, n281, n282, n283, n284, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n296, n297, n298, n299,
         n300, n301, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n403, n404,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n466, n467, n468, n469, n470, n471, n472, n473,
         n475, n476, n477, n478, n479, n481, n486, n490, n491, n492, n493,
         n494, n495, n498, n499, n500, n501, n502, n503, n504, n505, n510,
         n511, n514, n515, n516, n517, n518, n519, n524, n525, n526, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n546,
         n548, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848;
  wire   [3:0] FUNC;

  ALU_DATA_W32_DW01_sub_2 sub_128 ( .A({net34616, n113, n181, A[28:26], n242, 
        A[24:22], n49, A[20:13], net28420, A[11:10], n316, A[8:3], n309, A[1], 
        n274}), .B({B[31:30], n236, n248, B[27], n216, B[25:23], n32, B[21:20], 
        n27, B[18:2], n306, n191}), .CI(1'b0), .DIFF({N122, N121, N120, N119, 
        N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91}) );
  ALU_DATA_W32_DW01_add_2 add_125 ( .A({net34616, n113, n181, A[28:26], n241, 
        A[24:13], net28420, net41315, A[10], n318, A[8:3], n311, A[1], n321}), 
        .B({B[31:30], n236, n248, B[27], n216, B[25], n5, B[23], n213, B[21:2], 
        n307, n324}), .CI(1'b0), .SUM({N90, N89, N88, N87, N86, N85, N84, N83, 
        N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, N66, N65, N64, N63, N62, N61, N60, N59}) );
  ALU_DATA_W32_DW01_cmp6_1 r80 ( .A({B[31:29], n93, B[27:22], n59, B[20:19], 
        n34, n33, B[16], n201, n215, n276, n238, n223, n245, n218, n273, n222, 
        n221, n261, n278, net28241, net34566, n68, n225}), .B({A[31:26], n241, 
        A[24:22], n257, A[20:18], n281, A[16], n104, n235, n314, net28422, 
        net34655, A[10], n317, n320, n312, n187, n303, n305, n182, n310, n275, 
        n322}), .TC(1'b0), .LE(N794), .GE(N795), .NE(N796) );
  CLKBUF_X1 U3 ( .A(n230), .Z(n1) );
  CLKBUF_X3 U4 ( .A(net34351), .Z(net34889) );
  INV_X1 U6 ( .A(n559), .ZN(n2) );
  NOR2_X1 U7 ( .A1(n3), .A2(n4), .ZN(n681) );
  AND2_X1 U8 ( .A1(N82), .A2(net27181), .ZN(n3) );
  NAND2_X1 U9 ( .A1(n139), .A2(n138), .ZN(n4) );
  BUF_X1 U10 ( .A(B[24]), .Z(n5) );
  BUF_X2 U12 ( .A(A[22]), .Z(n6) );
  AND3_X1 U13 ( .A1(n484), .A2(n674), .A3(n642), .ZN(n244) );
  CLKBUF_X1 U15 ( .A(A[10]), .Z(n315) );
  INV_X1 U16 ( .A(n278), .ZN(n7) );
  INV_X1 U17 ( .A(n7), .ZN(n8) );
  NAND2_X2 U18 ( .A1(n366), .A2(net35893), .ZN(n546) );
  OR4_X2 U19 ( .A1(n222), .A2(B[6]), .A3(B[8]), .A4(B[9]), .ZN(n824) );
  OAI22_X1 U20 ( .A1(net25237), .A2(n166), .B1(net27195), .B2(n165), .ZN(
        net35986) );
  INV_X1 U21 ( .A(net25138), .ZN(n165) );
  INV_X1 U22 ( .A(net25136), .ZN(n166) );
  NAND4_X1 U23 ( .A1(n179), .A2(n19), .A3(n10), .A4(net25114), .ZN(net35985)
         );
  NAND2_X1 U24 ( .A1(n177), .A2(n181), .ZN(n179) );
  OAI22_X1 U25 ( .A1(net27165), .A2(n164), .B1(net27195), .B2(n158), .ZN(n168)
         );
  OAI21_X1 U26 ( .B1(net25237), .B2(n161), .A(n173), .ZN(n167) );
  INV_X1 U27 ( .A(net25132), .ZN(n164) );
  INV_X1 U28 ( .A(net25114), .ZN(n74) );
  BUF_X1 U29 ( .A(B[3]), .Z(net28242) );
  INV_X1 U30 ( .A(net34232), .ZN(n156) );
  INV_X1 U31 ( .A(net25443), .ZN(n171) );
  NAND2_X1 U32 ( .A1(net27203), .A2(n178), .ZN(n155) );
  INV_X1 U33 ( .A(n161), .ZN(n178) );
  NAND2_X1 U34 ( .A1(n232), .A2(net25131), .ZN(n173) );
  NAND2_X1 U35 ( .A1(n149), .A2(n150), .ZN(n480) );
  NAND2_X1 U36 ( .A1(n174), .A2(A[29]), .ZN(n150) );
  AND3_X1 U37 ( .A1(n521), .A2(n627), .A3(n598), .ZN(n133) );
  AND3_X1 U38 ( .A1(n508), .A2(n643), .A3(n613), .ZN(n240) );
  BUF_X1 U39 ( .A(net20206), .Z(net27179) );
  BUF_X1 U40 ( .A(n517), .Z(n122) );
  INV_X1 U41 ( .A(net25113), .ZN(n80) );
  INV_X1 U42 ( .A(n133), .ZN(n593) );
  BUF_X1 U43 ( .A(A[0]), .Z(n321) );
  NAND2_X1 U44 ( .A1(net35871), .A2(n74), .ZN(net25366) );
  OAI221_X1 U45 ( .B1(n842), .B2(net35616), .C1(n841), .C2(net27408), .A(n513), 
        .ZN(net25130) );
  INV_X1 U46 ( .A(n55), .ZN(n417) );
  BUF_X1 U47 ( .A(net33654), .Z(net27181) );
  INV_X1 U48 ( .A(n79), .ZN(n81) );
  AOI211_X1 U49 ( .C1(net35985), .C2(net35893), .A(net35986), .B(n12), .ZN(n78) );
  BUF_X1 U50 ( .A(A[2]), .Z(n309) );
  INV_X1 U51 ( .A(n244), .ZN(n500) );
  BUF_X1 U52 ( .A(n84), .Z(net27191) );
  NAND2_X1 U53 ( .A1(n169), .A2(n171), .ZN(n153) );
  NOR2_X1 U54 ( .A1(net25114), .A2(n156), .ZN(n152) );
  NAND2_X1 U55 ( .A1(net27527), .A2(net25442), .ZN(n169) );
  NAND2_X1 U56 ( .A1(net25238), .A2(net35893), .ZN(n154) );
  AND2_X1 U57 ( .A1(net27165), .A2(net34616), .ZN(n9) );
  OR2_X1 U58 ( .A1(net34836), .A2(n160), .ZN(n10) );
  INV_X1 U59 ( .A(net34906), .ZN(n177) );
  AND3_X1 U60 ( .A1(n141), .A2(n142), .A3(n143), .ZN(n11) );
  AND2_X1 U61 ( .A1(net25137), .A2(n232), .ZN(n12) );
  INV_X1 U62 ( .A(net27195), .ZN(net27201) );
  OR2_X1 U63 ( .A1(n261), .A2(B[31]), .ZN(n13) );
  OR2_X1 U64 ( .A1(B[18]), .A2(B[16]), .ZN(n14) );
  AND2_X1 U65 ( .A1(n349), .A2(n350), .ZN(n15) );
  AND2_X1 U66 ( .A1(n77), .A2(n76), .ZN(n16) );
  INV_X1 U67 ( .A(net25130), .ZN(n161) );
  OR2_X1 U68 ( .A1(n180), .A2(net20044), .ZN(n19) );
  OR2_X1 U69 ( .A1(net25236), .A2(net25237), .ZN(n20) );
  INV_X1 U70 ( .A(n439), .ZN(n22) );
  INV_X1 U71 ( .A(n63), .ZN(net34906) );
  BUF_X1 U72 ( .A(net35631), .Z(net27151) );
  CLKBUF_X1 U73 ( .A(n42), .Z(n23) );
  AND2_X1 U74 ( .A1(n42), .A2(net35893), .ZN(n24) );
  INV_X1 U75 ( .A(net27165), .ZN(net35893) );
  AND2_X2 U76 ( .A1(n42), .A2(n232), .ZN(n299) );
  INV_X1 U77 ( .A(n23), .ZN(net25596) );
  CLKBUF_X1 U78 ( .A(n267), .Z(n25) );
  INV_X1 U79 ( .A(n553), .ZN(n26) );
  AND3_X1 U80 ( .A1(n675), .A2(n706), .A3(n506), .ZN(n108) );
  BUF_X1 U81 ( .A(A[16]), .Z(n226) );
  CLKBUF_X1 U82 ( .A(B[19]), .Z(n27) );
  CLKBUF_X1 U83 ( .A(n114), .Z(n28) );
  AND3_X1 U84 ( .A1(n691), .A2(n659), .A3(n520), .ZN(n114) );
  BUF_X1 U85 ( .A(n324), .Z(n29) );
  BUF_X1 U86 ( .A(B[1]), .Z(n308) );
  INV_X1 U87 ( .A(n256), .ZN(n577) );
  AND3_X1 U88 ( .A1(n483), .A2(n612), .A3(n588), .ZN(n256) );
  CLKBUF_X1 U89 ( .A(B[27]), .Z(n30) );
  INV_X1 U90 ( .A(n546), .ZN(n31) );
  BUF_X1 U91 ( .A(net20206), .Z(net27177) );
  AOI221_X1 U92 ( .B1(n736), .B2(net25231), .C1(n30), .C2(n735), .A(n761), 
        .ZN(n749) );
  INV_X1 U93 ( .A(net27159), .ZN(net35616) );
  CLKBUF_X1 U94 ( .A(B[22]), .Z(n32) );
  CLKBUF_X1 U95 ( .A(B[17]), .Z(n33) );
  CLKBUF_X1 U96 ( .A(B[18]), .Z(n34) );
  INV_X1 U97 ( .A(n191), .ZN(n35) );
  BUF_X1 U98 ( .A(n338), .Z(n36) );
  BUF_X1 U99 ( .A(B[3]), .Z(net28241) );
  INV_X1 U100 ( .A(net27141), .ZN(net27137) );
  CLKBUF_X1 U101 ( .A(net25169), .Z(n37) );
  OR2_X1 U102 ( .A1(net27143), .A2(n73), .ZN(n38) );
  NAND2_X1 U103 ( .A1(n38), .A2(net25583), .ZN(net25484) );
  CLKBUF_X1 U104 ( .A(n308), .Z(n68) );
  NAND2_X1 U105 ( .A1(N73), .A2(net27183), .ZN(n39) );
  NAND2_X1 U106 ( .A1(n92), .A2(n529), .ZN(n40) );
  NAND2_X1 U107 ( .A1(N105), .A2(net27191), .ZN(n41) );
  AND3_X1 U108 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n530) );
  BUF_X1 U109 ( .A(net33654), .Z(net27183) );
  INV_X1 U110 ( .A(n28), .ZN(n529) );
  AND2_X2 U111 ( .A1(n69), .A2(net33657), .ZN(n42) );
  INV_X1 U112 ( .A(n219), .ZN(net27141) );
  AND2_X1 U113 ( .A1(n478), .A2(n745), .ZN(n43) );
  AND2_X1 U114 ( .A1(n286), .A2(net25131), .ZN(n44) );
  AND2_X1 U115 ( .A1(n744), .A2(net25130), .ZN(n45) );
  NOR3_X1 U116 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n453) );
  CLKBUF_X3 U117 ( .A(A[13]), .Z(n314) );
  INV_X2 U118 ( .A(n232), .ZN(net18434) );
  NOR2_X2 U119 ( .A1(net20020), .A2(net20024), .ZN(n232) );
  AND2_X1 U120 ( .A1(n189), .A2(n458), .ZN(n46) );
  AND2_X1 U121 ( .A1(n479), .A2(n696), .ZN(n47) );
  AND2_X1 U122 ( .A1(net27209), .A2(n632), .ZN(n48) );
  NOR3_X1 U123 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n403) );
  OR4_X1 U124 ( .A1(B[27]), .A2(B[26]), .A3(B[29]), .A4(B[28]), .ZN(n823) );
  BUF_X1 U125 ( .A(A[17]), .Z(n281) );
  BUF_X1 U126 ( .A(B[7]), .Z(n222) );
  BUF_X1 U127 ( .A(B[0]), .Z(n324) );
  NOR2_X1 U128 ( .A1(n167), .A2(n168), .ZN(net35981) );
  INV_X1 U129 ( .A(net25238), .ZN(n158) );
  NAND2_X1 U130 ( .A1(n348), .A2(n15), .ZN(RES[0]) );
  CLKBUF_X1 U131 ( .A(A[21]), .Z(n49) );
  NAND2_X1 U132 ( .A1(N78), .A2(net27183), .ZN(n50) );
  NAND2_X1 U133 ( .A1(n296), .A2(net25132), .ZN(n51) );
  NAND2_X1 U134 ( .A1(N110), .A2(net27191), .ZN(n52) );
  AND3_X1 U135 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n617) );
  BUF_X2 U136 ( .A(net20206), .Z(n53) );
  BUF_X2 U137 ( .A(net20206), .Z(n54) );
  AND3_X2 U138 ( .A1(n482), .A2(n738), .A3(n705), .ZN(n55) );
  BUF_X1 U139 ( .A(B[10]), .Z(n56) );
  OR2_X1 U140 ( .A1(net18434), .A2(net25169), .ZN(n57) );
  NAND2_X1 U141 ( .A1(n57), .A2(n579), .ZN(n408) );
  BUF_X1 U142 ( .A(n408), .Z(n94) );
  AND2_X1 U143 ( .A1(n8), .A2(n284), .ZN(n58) );
  CLKBUF_X1 U144 ( .A(B[21]), .Z(n59) );
  NAND2_X1 U145 ( .A1(N76), .A2(net27183), .ZN(n60) );
  NAND2_X1 U146 ( .A1(n297), .A2(n776), .ZN(n61) );
  NAND2_X1 U147 ( .A1(N108), .A2(net27191), .ZN(n62) );
  AND3_X1 U148 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n589) );
  NOR2_X1 U149 ( .A1(n112), .A2(n29), .ZN(n63) );
  NAND2_X1 U150 ( .A1(N74), .A2(net27183), .ZN(n64) );
  NAND2_X1 U151 ( .A1(n92), .A2(n553), .ZN(n65) );
  NAND2_X1 U152 ( .A1(N106), .A2(net27191), .ZN(n66) );
  AND3_X1 U153 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n554) );
  INV_X1 U154 ( .A(n108), .ZN(n553) );
  BUF_X1 U155 ( .A(B[0]), .Z(n282) );
  NAND2_X1 U156 ( .A1(n307), .A2(n282), .ZN(net33834) );
  BUF_X2 U157 ( .A(A[21]), .Z(n257) );
  BUF_X2 U158 ( .A(B[2]), .Z(net34566) );
  BUF_X1 U159 ( .A(net27127), .Z(net35004) );
  BUF_X1 U160 ( .A(B[4]), .Z(n278) );
  CLKBUF_X1 U161 ( .A(net25464), .Z(n67) );
  AND2_X1 U162 ( .A1(n210), .A2(n284), .ZN(n69) );
  NAND2_X1 U163 ( .A1(net27205), .A2(net25130), .ZN(n70) );
  NAND2_X1 U164 ( .A1(n92), .A2(n449), .ZN(n71) );
  NAND2_X1 U165 ( .A1(n478), .A2(n679), .ZN(n72) );
  AND3_X1 U166 ( .A1(n70), .A2(n71), .A3(n72), .ZN(n393) );
  NAND3_X1 U167 ( .A1(net25116), .A2(n75), .A3(n16), .ZN(RES[31]) );
  NAND2_X1 U168 ( .A1(B[31]), .A2(net25121), .ZN(n76) );
  OAI21_X1 U169 ( .B1(net34616), .B2(net27081), .A(net27103), .ZN(net25121) );
  INV_X1 U170 ( .A(net27105), .ZN(net27103) );
  INV_X2 U171 ( .A(net27095), .ZN(net27081) );
  MUX2_X1 U172 ( .A(net27095), .B(net33647), .S(B[30]), .Z(net25146) );
  AOI21_X1 U173 ( .B1(net27095), .B2(net25502), .A(net27105), .ZN(net25499) );
  AOI21_X1 U174 ( .B1(net27095), .B2(net25527), .A(net27105), .ZN(net25523) );
  CLKBUF_X1 U175 ( .A(net39040), .Z(net34616) );
  INV_X1 U176 ( .A(n73), .ZN(net39040) );
  INV_X1 U177 ( .A(A[31]), .ZN(n73) );
  OAI21_X1 U178 ( .B1(n54), .B2(n73), .A(net25112), .ZN(net25577) );
  OAI21_X1 U179 ( .B1(net34835), .B2(n73), .A(net25112), .ZN(net25464) );
  NAND2_X1 U180 ( .A1(n80), .A2(n74), .ZN(n77) );
  NAND2_X1 U181 ( .A1(n81), .A2(net33829), .ZN(n75) );
  MUX2_X1 U182 ( .A(net35981), .B(n78), .S(n82), .Z(n79) );
  INV_X1 U183 ( .A(n58), .ZN(n82) );
  INV_X2 U184 ( .A(n82), .ZN(net38433) );
  NAND2_X1 U185 ( .A1(N122), .A2(net27189), .ZN(n85) );
  AND3_X1 U186 ( .A1(n85), .A2(net34297), .A3(net34298), .ZN(net25116) );
  BUF_X1 U187 ( .A(n84), .Z(net27189) );
  AND3_X1 U188 ( .A1(FUNC[0]), .A2(net33684), .A3(n83), .ZN(n84) );
  BUF_X1 U189 ( .A(n84), .Z(net27187) );
  INV_X1 U190 ( .A(FUNC[2]), .ZN(n83) );
  AND3_X1 U191 ( .A1(net33684), .A2(n83), .A3(net25629), .ZN(net33654) );
  AND3_X1 U192 ( .A1(net33169), .A2(n83), .A3(net25629), .ZN(net33647) );
  NAND3_X1 U193 ( .A1(FUNC[0]), .A2(net33169), .A3(n83), .ZN(n124) );
  NAND3_X1 U194 ( .A1(FUNC[2]), .A2(net33684), .A3(net25629), .ZN(n123) );
  AND2_X1 U195 ( .A1(net33190), .A2(net33684), .ZN(net33657) );
  BUF_X1 U196 ( .A(A[11]), .Z(net41315) );
  CLKBUF_X1 U197 ( .A(A[25]), .Z(n241) );
  BUF_X2 U198 ( .A(A[25]), .Z(n242) );
  NAND2_X1 U199 ( .A1(net27203), .A2(n288), .ZN(n86) );
  AND2_X1 U200 ( .A1(N97), .A2(net27187), .ZN(n87) );
  AND2_X1 U201 ( .A1(n98), .A2(n175), .ZN(n88) );
  AND2_X1 U202 ( .A1(n31), .A2(n176), .ZN(n89) );
  NOR3_X1 U203 ( .A1(n89), .A2(n88), .A3(n87), .ZN(n384) );
  CLKBUF_X1 U204 ( .A(A[20]), .Z(n90) );
  CLKBUF_X1 U205 ( .A(n8), .Z(n91) );
  AND2_X2 U206 ( .A1(net20105), .A2(n288), .ZN(n92) );
  INV_X1 U207 ( .A(net25237), .ZN(net20105) );
  OR2_X1 U208 ( .A1(n535), .A2(n411), .ZN(n581) );
  BUF_X1 U209 ( .A(A[9]), .Z(n316) );
  INV_X1 U210 ( .A(net27408), .ZN(n174) );
  BUF_X1 U211 ( .A(B[28]), .Z(n93) );
  BUF_X2 U212 ( .A(A[7]), .Z(n312) );
  INV_X1 U213 ( .A(n134), .ZN(n95) );
  BUF_X1 U214 ( .A(A[4]), .Z(n305) );
  AND2_X1 U215 ( .A1(net28242), .A2(net34566), .ZN(net35871) );
  BUF_X1 U216 ( .A(B[1]), .Z(n306) );
  BUF_X1 U217 ( .A(B[1]), .Z(n307) );
  AND2_X1 U218 ( .A1(n236), .A2(n787), .ZN(n96) );
  AND2_X1 U219 ( .A1(net33829), .A2(n786), .ZN(n97) );
  NOR3_X1 U220 ( .A1(n96), .A2(n97), .A3(n785), .ZN(n793) );
  BUF_X1 U221 ( .A(B[10]), .Z(n245) );
  INV_X1 U222 ( .A(n566), .ZN(n98) );
  CLKBUF_X1 U223 ( .A(n34), .Z(n99) );
  NOR2_X1 U224 ( .A1(n152), .A2(n153), .ZN(net25429) );
  AND2_X1 U225 ( .A1(n479), .A2(n728), .ZN(n100) );
  AND2_X1 U226 ( .A1(n286), .A2(n800), .ZN(n101) );
  AND2_X1 U227 ( .A1(n744), .A2(n801), .ZN(n102) );
  NOR3_X1 U228 ( .A1(n100), .A2(n101), .A3(n102), .ZN(n437) );
  AOI221_X1 U229 ( .B1(n788), .B2(n94), .C1(n292), .C2(n119), .A(n585), .ZN(
        n591) );
  CLKBUF_X1 U230 ( .A(n33), .Z(n103) );
  AND4_X2 U231 ( .A1(n826), .A2(n825), .A3(n828), .A4(n827), .ZN(n284) );
  CLKBUF_X1 U232 ( .A(B[11]), .Z(n223) );
  INV_X2 U233 ( .A(n180), .ZN(net27123) );
  CLKBUF_X3 U234 ( .A(net33834), .Z(n180) );
  BUF_X1 U235 ( .A(A[15]), .Z(n104) );
  NAND2_X1 U236 ( .A1(n293), .A2(n728), .ZN(n105) );
  NAND2_X1 U237 ( .A1(n296), .A2(n795), .ZN(n106) );
  NAND2_X1 U238 ( .A1(n743), .A2(n794), .ZN(n107) );
  AND3_X1 U239 ( .A1(n105), .A2(n106), .A3(n107), .ZN(n730) );
  BUF_X2 U240 ( .A(n784), .Z(n293) );
  BUF_X1 U241 ( .A(B[9]), .Z(n218) );
  BUF_X1 U242 ( .A(A[12]), .Z(net28420) );
  CLKBUF_X1 U243 ( .A(B[6]), .Z(n221) );
  AOI21_X1 U244 ( .B1(net39040), .B2(n68), .A(n480), .ZN(n338) );
  OR2_X1 U245 ( .A1(n338), .A2(net18434), .ZN(n109) );
  NAND2_X1 U246 ( .A1(n579), .A2(n109), .ZN(n409) );
  BUF_X1 U247 ( .A(n409), .Z(n119) );
  AND2_X1 U248 ( .A1(n479), .A2(n742), .ZN(n110) );
  AND2_X1 U249 ( .A1(net27525), .A2(n445), .ZN(n111) );
  NOR3_X1 U250 ( .A1(n110), .A2(n111), .A3(n444), .ZN(n455) );
  NOR3_X1 U251 ( .A1(n824), .A2(B[30]), .A3(n13), .ZN(n825) );
  BUF_X1 U252 ( .A(B[5]), .Z(n261) );
  INV_X1 U253 ( .A(n306), .ZN(n112) );
  BUF_X2 U254 ( .A(A[30]), .Z(n113) );
  INV_X1 U255 ( .A(n294), .ZN(n115) );
  INV_X1 U256 ( .A(net25503), .ZN(n116) );
  AND2_X1 U257 ( .A1(net27207), .A2(net25238), .ZN(n117) );
  AND2_X1 U258 ( .A1(n92), .A2(n606), .ZN(n118) );
  NOR3_X1 U259 ( .A1(n117), .A2(n118), .A3(n450), .ZN(n452) );
  BUF_X1 U260 ( .A(n24), .Z(net27207) );
  INV_X1 U261 ( .A(n240), .ZN(n606) );
  CLKBUF_X1 U262 ( .A(B[8]), .Z(n273) );
  AOI221_X4 U263 ( .B1(n303), .B2(net35005), .C1(n305), .C2(net27131), .A(n272), .ZN(n271) );
  BUF_X1 U264 ( .A(n552), .Z(n190) );
  CLKBUF_X1 U265 ( .A(n207), .Z(n120) );
  BUF_X1 U266 ( .A(n517), .Z(n125) );
  BUF_X1 U267 ( .A(n517), .Z(n126) );
  NAND2_X1 U268 ( .A1(n42), .A2(net27203), .ZN(n517) );
  AND2_X1 U269 ( .A1(n734), .A2(n733), .ZN(n128) );
  AND2_X1 U270 ( .A1(B[30]), .A2(n810), .ZN(n129) );
  AND2_X1 U271 ( .A1(net33829), .A2(n809), .ZN(n130) );
  NOR3_X1 U272 ( .A1(n129), .A2(n130), .A3(n808), .ZN(n814) );
  AND2_X1 U273 ( .A1(net33829), .A2(n766), .ZN(n131) );
  AND2_X1 U274 ( .A1(n765), .A2(A[28]), .ZN(n132) );
  NOR3_X1 U275 ( .A1(n131), .A2(n132), .A3(n764), .ZN(n770) );
  CLKBUF_X1 U276 ( .A(n425), .Z(n134) );
  OR2_X1 U277 ( .A1(net18434), .A2(net25143), .ZN(n135) );
  NAND2_X1 U278 ( .A1(n135), .A2(n11), .ZN(n266) );
  CLKBUF_X1 U279 ( .A(n723), .Z(n137) );
  INV_X2 U280 ( .A(n468), .ZN(n478) );
  NAND2_X1 U281 ( .A1(n287), .A2(net25132), .ZN(n138) );
  NAND2_X1 U282 ( .A1(N114), .A2(net27189), .ZN(n139) );
  OR2_X1 U283 ( .A1(net18434), .A2(net25150), .ZN(n140) );
  NAND2_X1 U284 ( .A1(n140), .A2(n11), .ZN(n267) );
  OR2_X1 U285 ( .A1(n594), .A2(net25237), .ZN(n141) );
  OR2_X1 U286 ( .A1(net27167), .A2(n133), .ZN(n142) );
  OR2_X1 U287 ( .A1(n114), .A2(net27195), .ZN(n143) );
  NAND2_X2 U288 ( .A1(net28242), .A2(net20020), .ZN(net25237) );
  NAND2_X2 U289 ( .A1(net34566), .A2(net20024), .ZN(net27195) );
  NAND2_X1 U290 ( .A1(N121), .A2(net27187), .ZN(n144) );
  NAND2_X1 U291 ( .A1(N89), .A2(net27181), .ZN(n145) );
  INV_X1 U292 ( .A(n812), .ZN(n147) );
  AND3_X1 U293 ( .A1(n145), .A2(n144), .A3(n147), .ZN(n813) );
  INV_X2 U294 ( .A(n180), .ZN(net27121) );
  NAND3_X1 U295 ( .A1(n20), .A2(n154), .A3(n155), .ZN(net25231) );
  INV_X1 U296 ( .A(net34351), .ZN(net35631) );
  INV_X1 U297 ( .A(net27151), .ZN(net34836) );
  BUF_X4 U298 ( .A(net18431), .Z(net27165) );
  CLKBUF_X1 U299 ( .A(net18431), .Z(net27167) );
  NAND2_X1 U300 ( .A1(n42), .A2(net35893), .ZN(net25503) );
  INV_X1 U301 ( .A(A[29]), .ZN(net20047) );
  INV_X1 U302 ( .A(net20047), .ZN(n181) );
  CLKBUF_X1 U303 ( .A(net34889), .Z(net35624) );
  INV_X1 U304 ( .A(A[30]), .ZN(n160) );
  OR2_X1 U305 ( .A1(n160), .A2(net34835), .ZN(n149) );
  CLKBUF_X1 U306 ( .A(A[3]), .Z(n182) );
  INV_X1 U307 ( .A(n839), .ZN(n185) );
  BUF_X1 U308 ( .A(A[9]), .Z(n318) );
  CLKBUF_X1 U309 ( .A(A[6]), .Z(n187) );
  BUF_X2 U310 ( .A(net27127), .Z(net35005) );
  BUF_X1 U311 ( .A(net27125), .Z(net35006) );
  INV_X1 U312 ( .A(net33834), .ZN(net27125) );
  INV_X1 U313 ( .A(n676), .ZN(n188) );
  BUF_X1 U314 ( .A(B[0]), .Z(n191) );
  INV_X1 U315 ( .A(n58), .ZN(net34986) );
  INV_X1 U316 ( .A(n548), .ZN(n189) );
  NAND2_X2 U317 ( .A1(n366), .A2(n232), .ZN(n548) );
  CLKBUF_X1 U318 ( .A(n309), .Z(n193) );
  CLKBUF_X1 U319 ( .A(n59), .Z(n194) );
  CLKBUF_X1 U320 ( .A(n27), .Z(n199) );
  INV_X1 U321 ( .A(n112), .ZN(n200) );
  BUF_X1 U322 ( .A(B[15]), .Z(n201) );
  INV_X1 U323 ( .A(n225), .ZN(n212) );
  CLKBUF_X1 U324 ( .A(B[22]), .Z(n213) );
  CLKBUF_X1 U325 ( .A(B[14]), .Z(n215) );
  CLKBUF_X1 U326 ( .A(B[26]), .Z(n216) );
  INV_X1 U327 ( .A(net27179), .ZN(net34869) );
  INV_X1 U328 ( .A(net27143), .ZN(net34866) );
  BUF_X1 U329 ( .A(A[2]), .Z(n311) );
  CLKBUF_X1 U330 ( .A(net41315), .Z(net34655) );
  INV_X2 U331 ( .A(net35631), .ZN(net34835) );
  INV_X1 U332 ( .A(n355), .ZN(n224) );
  OAI221_X4 U333 ( .B1(n846), .B2(net34836), .C1(n845), .C2(n329), .A(n512), 
        .ZN(net25131) );
  INV_X1 U334 ( .A(n35), .ZN(n225) );
  NOR3_X1 U335 ( .A1(n822), .A2(n33), .A3(n14), .ZN(n827) );
  AND2_X1 U336 ( .A1(N95), .A2(net27187), .ZN(n227) );
  AND2_X1 U337 ( .A1(n92), .A2(n457), .ZN(n228) );
  AND2_X1 U338 ( .A1(n196), .A2(n768), .ZN(n229) );
  NOR3_X1 U339 ( .A1(n229), .A2(n228), .A3(n227), .ZN(n368) );
  INV_X1 U340 ( .A(n546), .ZN(n230) );
  INV_X1 U341 ( .A(n614), .ZN(n231) );
  INV_X1 U342 ( .A(n599), .ZN(n233) );
  CLKBUF_X1 U343 ( .A(n222), .Z(n234) );
  CLKBUF_X1 U344 ( .A(A[14]), .Z(n235) );
  CLKBUF_X1 U345 ( .A(B[29]), .Z(n236) );
  CLKBUF_X1 U346 ( .A(n439), .Z(n237) );
  BUF_X1 U347 ( .A(B[12]), .Z(n238) );
  CLKBUF_X1 U348 ( .A(n201), .Z(n243) );
  INV_X1 U349 ( .A(n284), .ZN(n294) );
  OR4_X1 U350 ( .A1(B[20]), .A2(B[19]), .A3(B[21]), .A4(B[22]), .ZN(n822) );
  INV_X1 U351 ( .A(n761), .ZN(n246) );
  NAND2_X1 U352 ( .A1(n784), .A2(n9), .ZN(n734) );
  CLKBUF_X1 U353 ( .A(n93), .Z(n248) );
  CLKBUF_X1 U354 ( .A(n316), .Z(n317) );
  INV_X1 U355 ( .A(n599), .ZN(n249) );
  NAND2_X1 U356 ( .A1(N120), .A2(net27187), .ZN(n250) );
  NAND2_X1 U357 ( .A1(N88), .A2(net27181), .ZN(n251) );
  INV_X1 U358 ( .A(n791), .ZN(n252) );
  AND3_X1 U359 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n792) );
  CLKBUF_X1 U360 ( .A(n238), .Z(n255) );
  AOI221_X4 U361 ( .B1(n242), .B2(net27123), .C1(A[26]), .C2(net34866), .A(
        n302), .ZN(n295) );
  AOI221_X4 U362 ( .B1(n304), .B2(net27123), .C1(n323), .C2(n177), .A(n416), 
        .ZN(n415) );
  CLKBUF_X1 U363 ( .A(n221), .Z(n260) );
  CLKBUF_X1 U364 ( .A(n215), .Z(n262) );
  BUF_X1 U365 ( .A(A[0]), .Z(n274) );
  CLKBUF_X1 U366 ( .A(A[1]), .Z(n275) );
  CLKBUF_X1 U367 ( .A(B[13]), .Z(n276) );
  CLKBUF_X1 U368 ( .A(n273), .Z(n277) );
  CLKBUF_X1 U369 ( .A(n218), .Z(n280) );
  CLKBUF_X1 U370 ( .A(A[8]), .Z(n319) );
  CLKBUF_X1 U371 ( .A(A[20]), .Z(n283) );
  INV_X1 U372 ( .A(n516), .ZN(n286) );
  INV_X1 U373 ( .A(n516), .ZN(n287) );
  INV_X1 U374 ( .A(n516), .ZN(n743) );
  NAND2_X1 U375 ( .A1(n582), .A2(n581), .ZN(n288) );
  NAND2_X1 U376 ( .A1(N86), .A2(net27181), .ZN(n289) );
  NAND2_X1 U377 ( .A1(n299), .A2(net25132), .ZN(n290) );
  NAND2_X1 U378 ( .A1(N118), .A2(net27189), .ZN(n291) );
  AND3_X1 U379 ( .A1(n289), .A2(n290), .A3(n291), .ZN(n746) );
  INV_X1 U380 ( .A(net27201), .ZN(net27193) );
  BUF_X2 U381 ( .A(n784), .Z(n292) );
  NAND2_X1 U382 ( .A1(n282), .A2(n848), .ZN(net34351) );
  INV_X1 U383 ( .A(n122), .ZN(n296) );
  INV_X1 U384 ( .A(n122), .ZN(n297) );
  NAND2_X1 U385 ( .A1(N90), .A2(net27183), .ZN(net34297) );
  NAND2_X1 U386 ( .A1(net34616), .A2(n816), .ZN(net34298) );
  BUF_X2 U387 ( .A(n24), .Z(net27205) );
  BUF_X1 U388 ( .A(n24), .Z(net27209) );
  INV_X1 U389 ( .A(n546), .ZN(n768) );
  INV_X1 U390 ( .A(n122), .ZN(n744) );
  INV_X1 U391 ( .A(net27143), .ZN(net27131) );
  INV_X1 U392 ( .A(net27141), .ZN(net27133) );
  AND2_X2 U393 ( .A1(n736), .A2(net27175), .ZN(n298) );
  INV_X1 U394 ( .A(n582), .ZN(n784) );
  INV_X1 U395 ( .A(n566), .ZN(n552) );
  AND2_X1 U396 ( .A1(n478), .A2(net27175), .ZN(net34232) );
  INV_X1 U397 ( .A(n581), .ZN(n788) );
  AND2_X1 U398 ( .A1(n736), .A2(net27203), .ZN(n300) );
  INV_X1 U399 ( .A(n219), .ZN(net27143) );
  AOI22_X1 U400 ( .A1(n163), .A2(net27203), .B1(n162), .B2(net20105), .ZN(n211) );
  AOI22_X1 U401 ( .A1(n176), .A2(net27203), .B1(n175), .B2(net20105), .ZN(n269) );
  AOI22_X1 U402 ( .A1(n186), .A2(net27203), .B1(n136), .B2(net20105), .ZN(n412) );
  NOR2_X1 U403 ( .A1(n239), .A2(n294), .ZN(n208) );
  INV_X1 U404 ( .A(net27105), .ZN(net27101) );
  OAI221_X1 U405 ( .B1(net34835), .B2(n819), .C1(n839), .C2(net18425), .A(n413), .ZN(n136) );
  OAI221_X1 U406 ( .B1(n839), .B2(net35624), .C1(net27408), .C2(n840), .A(n545), .ZN(n151) );
  OAI221_X1 U407 ( .B1(net34835), .B2(n842), .C1(net34869), .C2(n843), .A(n414), .ZN(n186) );
  OAI221_X1 U408 ( .B1(n839), .B2(n180), .C1(net34906), .C2(n840), .A(n270), 
        .ZN(n176) );
  OAI221_X1 U409 ( .B1(n180), .B2(n819), .C1(n839), .C2(net27143), .A(n214), 
        .ZN(n163) );
  OAI221_X1 U410 ( .B1(n268), .B2(n837), .C1(n208), .C2(n206), .A(net34986), 
        .ZN(n258) );
  OAI221_X1 U411 ( .B1(n209), .B2(n836), .C1(n208), .C2(n206), .A(net34986), 
        .ZN(n197) );
  OAI221_X1 U412 ( .B1(n410), .B2(n838), .C1(n208), .C2(n206), .A(net34986), 
        .ZN(n401) );
  INV_X1 U413 ( .A(net27095), .ZN(net27083) );
  OAI221_X1 U414 ( .B1(net35616), .B2(n843), .C1(n329), .C2(n844), .A(n544), 
        .ZN(n196) );
  NOR2_X1 U415 ( .A1(n848), .A2(n29), .ZN(n219) );
  OAI221_X1 U416 ( .B1(n328), .B2(net27081), .C1(net27113), .C2(n842), .A(
        net27103), .ZN(n172) );
  OAI22_X1 U417 ( .A1(n329), .A2(net20044), .B1(net34836), .B2(n818), .ZN(n302) );
  OAI22_X1 U418 ( .A1(n832), .A2(net18434), .B1(n217), .B2(net27165), .ZN(n209) );
  OAI22_X1 U419 ( .A1(n329), .A2(n845), .B1(net34835), .B2(n844), .ZN(n220) );
  OAI22_X1 U420 ( .A1(n833), .A2(net18434), .B1(n271), .B2(net27165), .ZN(n268) );
  OAI22_X1 U421 ( .A1(net27408), .A2(n846), .B1(net34835), .B2(n845), .ZN(n272) );
  OAI22_X1 U422 ( .A1(n834), .A2(net18434), .B1(n415), .B2(net27165), .ZN(n410) );
  OAI22_X1 U423 ( .A1(net27408), .A2(n847), .B1(net35624), .B2(n846), .ZN(n416) );
  OAI22_X1 U424 ( .A1(n835), .A2(net18434), .B1(n541), .B2(net27165), .ZN(n540) );
  AOI211_X1 U425 ( .C1(n323), .C2(net35006), .A(n542), .B(n817), .ZN(n541) );
  OAI22_X1 U426 ( .A1(net34836), .A2(n847), .B1(net34906), .B2(n846), .ZN(n542) );
  AND2_X1 U427 ( .A1(net33657), .A2(n115), .ZN(net33829) );
  BUF_X1 U428 ( .A(net33654), .Z(net27185) );
  INV_X1 U429 ( .A(net27195), .ZN(net27203) );
  OAI21_X1 U430 ( .B1(net28241), .B2(n123), .A(net27101), .ZN(n203) );
  AOI22_X1 U431 ( .A1(n408), .A2(n206), .B1(n409), .B2(n208), .ZN(n407) );
  AOI22_X1 U432 ( .A1(n266), .A2(n206), .B1(n267), .B2(n208), .ZN(n265) );
  AOI22_X1 U433 ( .A1(n205), .A2(n206), .B1(n207), .B2(n208), .ZN(n204) );
  NOR2_X1 U434 ( .A1(n411), .A2(n294), .ZN(n206) );
  AOI221_X1 U435 ( .B1(A[26]), .B2(net27123), .C1(A[27]), .C2(n177), .A(n285), 
        .ZN(n279) );
  OAI22_X1 U436 ( .A1(net34869), .A2(net20047), .B1(net34835), .B2(net20044), 
        .ZN(n285) );
  AOI211_X1 U437 ( .C1(A[27]), .C2(net27123), .A(n253), .B(n254), .ZN(n247) );
  OAI22_X1 U438 ( .A1(net35616), .A2(net20047), .B1(net20044), .B2(net27143), 
        .ZN(n253) );
  AOI22_X1 U439 ( .A1(n257), .A2(net27127), .B1(A[20]), .B2(n63), .ZN(n521) );
  AOI22_X1 U440 ( .A1(n6), .A2(net35004), .B1(n257), .B2(net27133), .ZN(n508)
         );
  AOI22_X1 U441 ( .A1(n90), .A2(net35004), .B1(n231), .B2(net27133), .ZN(n483)
         );
  NAND2_X1 U442 ( .A1(n232), .A2(net39040), .ZN(n378) );
  NAND2_X1 U443 ( .A1(net28242), .A2(net34616), .ZN(n339) );
  AOI221_X1 U444 ( .B1(n276), .B2(n486), .C1(net34232), .C2(net25484), .A(n481), .ZN(n504) );
  AOI22_X1 U445 ( .A1(A[27]), .A2(net27121), .B1(A[26]), .B2(net27137), .ZN(
        n547) );
  AOI22_X1 U446 ( .A1(n188), .A2(net27123), .B1(n6), .B2(net27131), .ZN(n550)
         );
  AOI22_X1 U447 ( .A1(A[24]), .A2(net27125), .B1(net27133), .B2(A[23]), .ZN(
        n484) );
  AND2_X1 U448 ( .A1(n332), .A2(n333), .ZN(net33684) );
  AOI22_X1 U449 ( .A1(A[28]), .A2(net27125), .B1(A[27]), .B2(net27133), .ZN(
        n482) );
  AOI22_X1 U450 ( .A1(A[26]), .A2(net27127), .B1(n242), .B2(net27133), .ZN(
        n506) );
  AOI22_X1 U451 ( .A1(n242), .A2(net27125), .B1(A[24]), .B2(n63), .ZN(n520) );
  INV_X1 U452 ( .A(n124), .ZN(net27105) );
  AND2_X1 U453 ( .A1(net39040), .A2(n364), .ZN(n301) );
  AOI221_X1 U454 ( .B1(n262), .B2(n514), .C1(net34232), .C2(n67), .A(n511), 
        .ZN(n533) );
  AOI221_X1 U455 ( .B1(n327), .B2(net33647), .C1(net27095), .C2(n847), .A(
        net27105), .ZN(n405) );
  AOI221_X1 U456 ( .B1(n309), .B2(net33647), .C1(net27095), .C2(n846), .A(
        net27105), .ZN(n263) );
  AOI221_X1 U457 ( .B1(n323), .B2(net33647), .C1(net27095), .C2(n845), .A(
        net27105), .ZN(n202) );
  AOI221_X1 U458 ( .B1(n298), .B2(net25131), .C1(n199), .C2(n610), .A(n718), 
        .ZN(n620) );
  AOI221_X1 U459 ( .B1(n478), .B2(n727), .C1(n430), .C2(n315), .A(n429), .ZN(
        n438) );
  AND2_X1 U460 ( .A1(FUNC[0]), .A2(FUNC[2]), .ZN(net33190) );
  AND2_X1 U461 ( .A1(FUNC[1]), .A2(n332), .ZN(net33169) );
  CLKBUF_X1 U462 ( .A(n274), .Z(n322) );
  CLKBUF_X1 U463 ( .A(A[5]), .Z(n303) );
  AOI22_X1 U464 ( .A1(n281), .A2(net27123), .B1(n226), .B2(net27131), .ZN(n523) );
  OAI21_X1 U465 ( .B1(n234), .B2(n123), .A(n124), .ZN(n157) );
  CLKBUF_X1 U466 ( .A(A[4]), .Z(n304) );
  CLKBUF_X1 U467 ( .A(A[12]), .Z(net28421) );
  CLKBUF_X1 U468 ( .A(A[12]), .Z(net28422) );
  CLKBUF_X1 U469 ( .A(A[2]), .Z(n310) );
  CLKBUF_X1 U470 ( .A(n312), .Z(n313) );
  OAI21_X1 U471 ( .B1(n260), .B2(n123), .A(n124), .ZN(n170) );
  OAI21_X1 U472 ( .B1(net34566), .B2(net27081), .A(net27101), .ZN(n264) );
  OAI21_X1 U473 ( .B1(n261), .B2(n123), .A(n124), .ZN(n183) );
  OAI21_X1 U474 ( .B1(n91), .B2(n123), .A(n124), .ZN(n192) );
  OAI21_X1 U475 ( .B1(n277), .B2(n123), .A(n124), .ZN(n146) );
  OAI21_X1 U476 ( .B1(n280), .B2(n123), .A(net27101), .ZN(n121) );
  BUF_X1 U477 ( .A(A[8]), .Z(n320) );
  INV_X1 U478 ( .A(n845), .ZN(n323) );
  OAI21_X1 U479 ( .B1(n200), .B2(net27081), .A(net27101), .ZN(n406) );
  INV_X1 U480 ( .A(n308), .ZN(n848) );
  INV_X1 U481 ( .A(net25448), .ZN(net27527) );
  INV_X1 U482 ( .A(net25527), .ZN(net27525) );
  INV_X1 U483 ( .A(n235), .ZN(n325) );
  INV_X1 U484 ( .A(n325), .ZN(n326) );
  AOI22_X1 U485 ( .A1(net38433), .A2(n830), .B1(n193), .B2(n264), .ZN(n259) );
  AOI22_X1 U486 ( .A1(n249), .A2(net35005), .B1(n281), .B2(net27131), .ZN(n507) );
  AOI22_X1 U487 ( .A1(n231), .A2(net27121), .B1(n249), .B2(net27137), .ZN(n549) );
  OAI221_X1 U488 ( .B1(n320), .B2(n123), .C1(net27113), .C2(n840), .A(net27103), .ZN(n148) );
  INV_X1 U489 ( .A(n847), .ZN(n327) );
  INV_X1 U490 ( .A(n842), .ZN(n328) );
  OAI221_X1 U491 ( .B1(n303), .B2(net27081), .C1(net27113), .C2(n843), .A(n124), .ZN(n184) );
  AOI221_X1 U492 ( .B1(n328), .B2(net27121), .C1(n303), .C2(net34866), .A(n220), .ZN(n217) );
  AOI22_X1 U493 ( .A1(n303), .A2(net27123), .B1(n328), .B2(n177), .ZN(n497) );
  OAI221_X1 U494 ( .B1(n185), .B2(n123), .C1(n839), .C2(net27113), .A(net27103), .ZN(n127) );
  AOI22_X1 U495 ( .A1(n310), .A2(net35005), .B1(n323), .B2(net34866), .ZN(n487) );
  AOI22_X1 U496 ( .A1(net38433), .A2(n829), .B1(n323), .B2(n203), .ZN(n198) );
  OAI221_X1 U497 ( .B1(n305), .B2(net27081), .C1(net27113), .C2(n844), .A(n124), .ZN(n195) );
  AOI22_X1 U498 ( .A1(n323), .A2(net35006), .B1(n304), .B2(net27137), .ZN(n528) );
  AOI22_X1 U499 ( .A1(n305), .A2(net35005), .B1(n303), .B2(net34866), .ZN(n513) );
  AOI22_X1 U500 ( .A1(n226), .A2(net35006), .B1(net27527), .B2(net34866), .ZN(
        n485) );
  AOI22_X1 U501 ( .A1(net27527), .A2(net35006), .B1(n326), .B2(net27131), .ZN(
        n543) );
  AOI22_X1 U502 ( .A1(n314), .A2(net35005), .B1(n326), .B2(net34866), .ZN(n454) );
  AOI22_X1 U503 ( .A1(net28421), .A2(net27123), .B1(n314), .B2(net27137), .ZN(
        n465) );
  AOI22_X1 U504 ( .A1(n326), .A2(net27121), .B1(n314), .B2(n177), .ZN(n509) );
  AOI22_X1 U505 ( .A1(n314), .A2(net35006), .B1(net28422), .B2(net27137), .ZN(
        n522) );
  AOI22_X1 U506 ( .A1(net27525), .A2(net35005), .B1(net28422), .B2(n177), .ZN(
        n474) );
  AOI22_X1 U507 ( .A1(n315), .A2(net27123), .B1(net27525), .B2(net27137), .ZN(
        n488) );
  AOI22_X1 U508 ( .A1(net27525), .A2(net35006), .B1(n315), .B2(net27131), .ZN(
        n545) );
  AOI22_X1 U509 ( .A1(net28421), .A2(net27123), .B1(net27525), .B2(net27131), 
        .ZN(n413) );
  OAI221_X1 U510 ( .B1(n313), .B2(n123), .C1(net27113), .C2(n841), .A(net27103), .ZN(n159) );
  AOI22_X1 U511 ( .A1(n313), .A2(net35006), .B1(n319), .B2(net27137), .ZN(n527) );
  AOI22_X1 U512 ( .A1(n312), .A2(net27121), .B1(n328), .B2(net27137), .ZN(n544) );
  AOI22_X1 U513 ( .A1(n328), .A2(net27123), .B1(n313), .B2(net34866), .ZN(n489) );
  AOI22_X1 U514 ( .A1(n313), .A2(net27149), .B1(n328), .B2(n53), .ZN(n270) );
  AOI22_X1 U515 ( .A1(n319), .A2(net35005), .B1(n312), .B2(net34866), .ZN(n414) );
  AOI22_X1 U516 ( .A1(n320), .A2(net27159), .B1(n313), .B2(net27179), .ZN(n214) );
  AOI22_X1 U517 ( .A1(n831), .A2(net38433), .B1(n327), .B2(n406), .ZN(n402) );
  AOI22_X1 U518 ( .A1(n321), .A2(net27123), .B1(n327), .B2(net27137), .ZN(n512) );
  AOI22_X1 U519 ( .A1(n327), .A2(net27121), .B1(n193), .B2(net34866), .ZN(n496) );
  INV_X1 U520 ( .A(n275), .ZN(n847) );
  NAND2_X1 U521 ( .A1(n112), .A2(n35), .ZN(net27408) );
  NAND2_X1 U522 ( .A1(n112), .A2(n212), .ZN(n329) );
  INV_X2 U523 ( .A(n469), .ZN(n479) );
  INV_X1 U524 ( .A(net27165), .ZN(net27175) );
  INV_X1 U525 ( .A(net34889), .ZN(net27149) );
  INV_X1 U526 ( .A(net34889), .ZN(net27155) );
  INV_X1 U527 ( .A(net34889), .ZN(net27159) );
  INV_X1 U528 ( .A(net34889), .ZN(net27161) );
  INV_X1 U529 ( .A(net33834), .ZN(net27127) );
  INV_X1 U530 ( .A(net33647), .ZN(net27113) );
  INV_X1 U531 ( .A(n123), .ZN(net27095) );
  INV_X1 U532 ( .A(FUNC[3]), .ZN(n332) );
  NAND2_X1 U533 ( .A1(net33190), .A2(net33169), .ZN(n239) );
  INV_X1 U534 ( .A(FUNC[0]), .ZN(net25629) );
  NAND3_X1 U535 ( .A1(net33169), .A2(FUNC[2]), .A3(net25629), .ZN(n411) );
  INV_X1 U536 ( .A(n282), .ZN(n820) );
  NAND2_X1 U537 ( .A1(n848), .A2(n820), .ZN(net18425) );
  INV_X1 U538 ( .A(net34566), .ZN(net20020) );
  INV_X1 U539 ( .A(net28242), .ZN(net20024) );
  NAND2_X1 U540 ( .A1(net20020), .A2(net20024), .ZN(net18431) );
  NAND2_X1 U541 ( .A1(n8), .A2(n284), .ZN(n210) );
  INV_X1 U542 ( .A(FUNC[1]), .ZN(n333) );
  MUX2_X1 U543 ( .A(net27083), .B(net27113), .S(n225), .Z(n330) );
  NAND2_X1 U544 ( .A1(n330), .A2(net27103), .ZN(n331) );
  AOI22_X1 U545 ( .A1(n224), .A2(n331), .B1(N91), .B2(net27189), .ZN(n350) );
  INV_X1 U546 ( .A(net18425), .ZN(net20206) );
  NAND2_X1 U547 ( .A1(n54), .A2(n322), .ZN(n685) );
  INV_X1 U548 ( .A(n685), .ZN(n817) );
  NAND2_X1 U549 ( .A1(n210), .A2(n284), .ZN(n535) );
  AOI22_X1 U550 ( .A1(n817), .A2(net27207), .B1(N59), .B2(net27185), .ZN(n349)
         );
  NOR2_X1 U551 ( .A1(FUNC[2]), .A2(n332), .ZN(n347) );
  MUX2_X1 U552 ( .A(N794), .B(N796), .S(FUNC[1]), .Z(n335) );
  AND2_X1 U553 ( .A1(N795), .A2(n333), .ZN(n334) );
  MUX2_X1 U554 ( .A(n335), .B(n334), .S(FUNC[0]), .Z(n346) );
  INV_X1 U555 ( .A(n322), .ZN(n355) );
  AOI21_X1 U556 ( .B1(net27095), .B2(n355), .A(net27105), .ZN(n344) );
  AOI221_X1 U557 ( .B1(n196), .B2(net27203), .C1(n151), .C2(net20105), .A(n540), .ZN(n341) );
  NAND2_X1 U558 ( .A1(n242), .A2(net27159), .ZN(n722) );
  NAND2_X1 U559 ( .A1(A[24]), .A2(n53), .ZN(n690) );
  NAND3_X1 U560 ( .A1(n547), .A2(n722), .A3(n690), .ZN(n456) );
  INV_X1 U561 ( .A(A[28]), .ZN(net20044) );
  AOI22_X1 U562 ( .A1(n113), .A2(net27137), .B1(net39040), .B2(net35005), .ZN(
        n336) );
  OAI221_X1 U563 ( .B1(net20047), .B2(net34835), .C1(net20044), .C2(net27408), 
        .A(n336), .ZN(n767) );
  NAND2_X1 U564 ( .A1(n257), .A2(net27161), .ZN(n658) );
  NAND2_X1 U565 ( .A1(n283), .A2(n53), .ZN(n626) );
  NAND3_X1 U566 ( .A1(n550), .A2(n658), .A3(n626), .ZN(n458) );
  INV_X1 U567 ( .A(n458), .ZN(n567) );
  NAND2_X1 U568 ( .A1(n281), .A2(net27149), .ZN(n597) );
  NAND2_X1 U569 ( .A1(n226), .A2(n53), .ZN(n563) );
  NAND3_X1 U570 ( .A1(n549), .A2(n597), .A3(n563), .ZN(n572) );
  INV_X1 U571 ( .A(n572), .ZN(n397) );
  OAI22_X1 U572 ( .A1(n567), .A2(net27195), .B1(net27165), .B2(n397), .ZN(n337) );
  AOI221_X1 U573 ( .B1(net20105), .B2(n456), .C1(n767), .C2(n232), .A(n337), 
        .ZN(n340) );
  MUX2_X1 U574 ( .A(n341), .B(n340), .S(net38433), .Z(n343) );
  INV_X1 U575 ( .A(n411), .ZN(n363) );
  INV_X1 U576 ( .A(n239), .ZN(n364) );
  OAI21_X1 U577 ( .B1(n363), .B2(n364), .A(n115), .ZN(n342) );
  OAI22_X1 U578 ( .A1(n212), .A2(n344), .B1(n343), .B2(n342), .ZN(n345) );
  NAND2_X1 U579 ( .A1(n301), .A2(n294), .ZN(n441) );
  INV_X1 U580 ( .A(n441), .ZN(n419) );
  AOI211_X1 U581 ( .C1(n347), .C2(n346), .A(n419), .B(n345), .ZN(n348) );
  AOI22_X1 U582 ( .A1(N92), .A2(net27187), .B1(N60), .B2(net27185), .ZN(n353)
         );
  INV_X1 U583 ( .A(n327), .ZN(n354) );
  OAI22_X1 U584 ( .A1(net34869), .A2(n354), .B1(net34836), .B2(n355), .ZN(n777) );
  NAND2_X1 U585 ( .A1(n402), .A2(n401), .ZN(n351) );
  AOI211_X1 U586 ( .C1(net27205), .C2(n777), .A(n419), .B(n351), .ZN(n352) );
  OAI211_X1 U587 ( .C1(n405), .C2(n112), .A(n353), .B(n352), .ZN(RES[1]) );
  AOI22_X1 U588 ( .A1(N93), .A2(net27187), .B1(N61), .B2(net27185), .ZN(n358)
         );
  INV_X1 U589 ( .A(n193), .ZN(n846) );
  OAI222_X1 U590 ( .A1(n846), .A2(n329), .B1(net34906), .B2(n355), .C1(
        net35624), .C2(n354), .ZN(n800) );
  NAND2_X1 U591 ( .A1(n259), .A2(n258), .ZN(n356) );
  AOI211_X1 U592 ( .C1(net27205), .C2(n800), .A(n419), .B(n356), .ZN(n357) );
  OAI211_X1 U593 ( .C1(n263), .C2(net20020), .A(n358), .B(n357), .ZN(RES[2])
         );
  AOI22_X1 U594 ( .A1(N94), .A2(net27187), .B1(N62), .B2(net27185), .ZN(n361)
         );
  INV_X1 U595 ( .A(n182), .ZN(n845) );
  NAND2_X1 U596 ( .A1(n198), .A2(n197), .ZN(n359) );
  AOI211_X1 U597 ( .C1(net27205), .C2(net25131), .A(n419), .B(n359), .ZN(n360)
         );
  OAI211_X1 U598 ( .C1(n202), .C2(net20024), .A(n361), .B(n360), .ZN(RES[3])
         );
  NAND2_X1 U599 ( .A1(n363), .A2(n58), .ZN(n468) );
  INV_X1 U600 ( .A(n767), .ZN(n467) );
  INV_X1 U601 ( .A(n456), .ZN(n569) );
  OAI222_X1 U602 ( .A1(n467), .A2(net25237), .B1(n569), .B2(net27193), .C1(
        net27165), .C2(n567), .ZN(n631) );
  NOR2_X1 U603 ( .A1(net28242), .A2(net25596), .ZN(n362) );
  INV_X1 U604 ( .A(n304), .ZN(n844) );
  OAI221_X1 U605 ( .B1(n845), .B2(net34836), .C1(n844), .C2(net27408), .A(n496), .ZN(n565) );
  INV_X1 U606 ( .A(n565), .ZN(n686) );
  MUX2_X1 U607 ( .A(n686), .B(n685), .S(net34566), .Z(n755) );
  INV_X1 U608 ( .A(n755), .ZN(n622) );
  AOI221_X1 U609 ( .B1(n478), .B2(n631), .C1(n362), .C2(n622), .A(n419), .ZN(
        n370) );
  NAND2_X1 U610 ( .A1(n69), .A2(n364), .ZN(n582) );
  NAND2_X1 U611 ( .A1(n582), .A2(n581), .ZN(n366) );
  NAND2_X1 U612 ( .A1(net27203), .A2(n288), .ZN(n566) );
  NAND2_X1 U613 ( .A1(n364), .A2(n58), .ZN(n469) );
  INV_X1 U614 ( .A(n631), .ZN(n365) );
  NAND2_X1 U615 ( .A1(n365), .A2(n378), .ZN(n633) );
  INV_X1 U616 ( .A(n548), .ZN(n571) );
  AOI222_X1 U617 ( .A1(n151), .A2(n98), .B1(n479), .B2(n633), .C1(n189), .C2(
        n572), .ZN(n369) );
  NAND2_X1 U618 ( .A1(net20105), .A2(n288), .ZN(n568) );
  NAND2_X1 U619 ( .A1(n314), .A2(net27149), .ZN(n525) );
  NAND2_X1 U620 ( .A1(net28421), .A2(net27179), .ZN(n460) );
  NAND3_X1 U621 ( .A1(n543), .A2(n525), .A3(n460), .ZN(n457) );
  AOI222_X1 U622 ( .A1(n192), .A2(n304), .B1(N63), .B2(net27185), .C1(n195), 
        .C2(n91), .ZN(n367) );
  NAND4_X1 U623 ( .A1(n369), .A2(n370), .A3(n368), .A4(n367), .ZN(RES[4]) );
  NAND2_X1 U624 ( .A1(n6), .A2(net27155), .ZN(n674) );
  NAND2_X1 U625 ( .A1(n257), .A2(n54), .ZN(n642) );
  NAND2_X1 U626 ( .A1(A[26]), .A2(net27155), .ZN(n738) );
  NAND2_X1 U627 ( .A1(n242), .A2(n54), .ZN(n705) );
  OAI22_X1 U628 ( .A1(net27165), .A2(n244), .B1(n55), .B2(net27193), .ZN(n371)
         );
  INV_X1 U629 ( .A(n371), .ZN(n373) );
  OAI211_X1 U630 ( .C1(n36), .C2(net25237), .A(n373), .B(n378), .ZN(n647) );
  NAND2_X1 U631 ( .A1(n233), .A2(net27161), .ZN(n612) );
  NAND2_X1 U632 ( .A1(n281), .A2(n53), .ZN(n588) );
  INV_X1 U633 ( .A(n777), .ZN(n420) );
  OAI21_X1 U634 ( .B1(n420), .B2(n126), .A(n441), .ZN(n372) );
  AOI221_X1 U635 ( .B1(n479), .B2(n647), .C1(n571), .C2(n577), .A(n372), .ZN(
        n377) );
  INV_X1 U636 ( .A(n303), .ZN(n843) );
  OAI221_X1 U637 ( .B1(n844), .B2(net35624), .C1(n843), .C2(n329), .A(n487), 
        .ZN(n778) );
  NAND2_X1 U638 ( .A1(n326), .A2(net27159), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n314), .A2(n53), .ZN(n494) );
  NAND3_X1 U640 ( .A1(n485), .A2(n539), .A3(n494), .ZN(n498) );
  INV_X1 U641 ( .A(n480), .ZN(net25583) );
  INV_X1 U642 ( .A(net25484), .ZN(net25169) );
  OAI21_X1 U643 ( .B1(n37), .B2(net25237), .A(n373), .ZN(n648) );
  AOI222_X1 U644 ( .A1(net27205), .A2(n778), .B1(n92), .B2(n498), .C1(n478), 
        .C2(n648), .ZN(n376) );
  AOI222_X1 U645 ( .A1(N96), .A2(net27187), .B1(n136), .B2(n552), .C1(n230), 
        .C2(n186), .ZN(n375) );
  AOI222_X1 U646 ( .A1(n183), .A2(n303), .B1(N64), .B2(net27185), .C1(n261), 
        .C2(n184), .ZN(n374) );
  NAND4_X1 U647 ( .A1(n375), .A2(n376), .A3(n377), .A4(n374), .ZN(RES[5]) );
  NAND2_X1 U648 ( .A1(net27525), .A2(net27149), .ZN(n461) );
  NAND2_X1 U649 ( .A1(net27179), .A2(n315), .ZN(n432) );
  NAND3_X1 U650 ( .A1(n522), .A2(n461), .A3(n432), .ZN(n175) );
  NAND2_X1 U651 ( .A1(net27179), .A2(n113), .ZN(net25112) );
  INV_X1 U652 ( .A(net25577), .ZN(net25150) );
  NAND2_X1 U653 ( .A1(A[23]), .A2(net27161), .ZN(n691) );
  NAND2_X1 U654 ( .A1(n6), .A2(net27177), .ZN(n659) );
  INV_X1 U655 ( .A(A[27]), .ZN(n818) );
  NAND2_X1 U656 ( .A1(A[26]), .A2(net27177), .ZN(n723) );
  AOI22_X1 U657 ( .A1(A[28]), .A2(n63), .B1(A[29]), .B2(net27125), .ZN(n379)
         );
  OAI211_X1 U658 ( .C1(n818), .C2(net34889), .A(n379), .B(n723), .ZN(n425) );
  INV_X1 U659 ( .A(n425), .ZN(n594) );
  OAI22_X1 U660 ( .A1(net27165), .A2(n28), .B1(n95), .B2(net27193), .ZN(n380)
         );
  INV_X1 U661 ( .A(n380), .ZN(n382) );
  OAI211_X1 U662 ( .C1(net25150), .C2(net25237), .A(n378), .B(n382), .ZN(n664)
         );
  NAND2_X1 U663 ( .A1(n231), .A2(net27155), .ZN(n627) );
  NAND2_X1 U664 ( .A1(n233), .A2(net27177), .ZN(n598) );
  INV_X1 U665 ( .A(n800), .ZN(n716) );
  OAI21_X1 U666 ( .B1(n716), .B2(n125), .A(n441), .ZN(n381) );
  AOI221_X1 U667 ( .B1(n479), .B2(n664), .C1(n571), .C2(n593), .A(n381), .ZN(
        n386) );
  INV_X1 U668 ( .A(n187), .ZN(n842) );
  OAI221_X1 U669 ( .B1(n843), .B2(net34835), .C1(n842), .C2(net34869), .A(n528), .ZN(n801) );
  NAND2_X1 U670 ( .A1(net27527), .A2(net27159), .ZN(n564) );
  NAND2_X1 U671 ( .A1(n326), .A2(net27179), .ZN(n524) );
  NAND3_X1 U672 ( .A1(n523), .A2(n564), .A3(n524), .ZN(n433) );
  INV_X1 U673 ( .A(net25464), .ZN(net25143) );
  OAI21_X1 U674 ( .B1(net25143), .B2(net25237), .A(n382), .ZN(n663) );
  AOI222_X1 U675 ( .A1(net27205), .A2(n801), .B1(n92), .B2(n433), .C1(n478), 
        .C2(n663), .ZN(n385) );
  AOI222_X1 U676 ( .A1(n170), .A2(n328), .B1(N65), .B2(net27185), .C1(n260), 
        .C2(n172), .ZN(n383) );
  NAND4_X1 U677 ( .A1(n384), .A2(n383), .A3(n386), .A4(n385), .ZN(RES[6]) );
  NAND2_X1 U678 ( .A1(net28422), .A2(net27161), .ZN(n495) );
  NAND2_X1 U679 ( .A1(net27525), .A2(n54), .ZN(n448) );
  NAND3_X1 U680 ( .A1(n509), .A2(n495), .A3(n448), .ZN(n162) );
  NAND2_X1 U681 ( .A1(A[24]), .A2(net27149), .ZN(n706) );
  NAND2_X1 U682 ( .A1(A[23]), .A2(net27179), .ZN(n675) );
  NAND2_X1 U683 ( .A1(net27177), .A2(A[27]), .ZN(n739) );
  AOI22_X1 U684 ( .A1(A[29]), .A2(n63), .B1(A[30]), .B2(net27127), .ZN(n387)
         );
  OAI211_X1 U685 ( .C1(net20044), .C2(net34889), .A(n739), .B(n387), .ZN(n439)
         );
  INV_X1 U686 ( .A(n439), .ZN(n607) );
  OAI22_X1 U687 ( .A1(net27165), .A2(n26), .B1(n607), .B2(net27193), .ZN(n388)
         );
  INV_X1 U688 ( .A(n388), .ZN(n390) );
  NAND2_X1 U689 ( .A1(n390), .A2(n339), .ZN(n680) );
  NAND2_X1 U690 ( .A1(n90), .A2(net27159), .ZN(n643) );
  NAND2_X1 U691 ( .A1(n231), .A2(n53), .ZN(n613) );
  INV_X1 U692 ( .A(net25131), .ZN(net25236) );
  OAI21_X1 U693 ( .B1(net25236), .B2(n126), .A(n441), .ZN(n389) );
  AOI221_X1 U694 ( .B1(n479), .B2(n680), .C1(n571), .C2(n606), .A(n389), .ZN(
        n394) );
  INV_X1 U695 ( .A(n312), .ZN(n841) );
  NAND2_X1 U696 ( .A1(n226), .A2(net27151), .ZN(n587) );
  NAND2_X1 U697 ( .A1(net27527), .A2(n54), .ZN(n538) );
  NAND3_X1 U698 ( .A1(n507), .A2(n587), .A3(n538), .ZN(n449) );
  NAND2_X1 U699 ( .A1(net39040), .A2(n54), .ZN(net25114) );
  OAI21_X1 U700 ( .B1(net25237), .B2(net25114), .A(n390), .ZN(n679) );
  AOI222_X1 U701 ( .A1(N98), .A2(net27187), .B1(n98), .B2(n162), .C1(n230), 
        .C2(n163), .ZN(n392) );
  AOI222_X1 U702 ( .A1(n157), .A2(n312), .B1(N66), .B2(net27185), .C1(n234), 
        .C2(n159), .ZN(n391) );
  NAND4_X1 U703 ( .A1(n392), .A2(n393), .A3(n394), .A4(n391), .ZN(RES[7]) );
  NAND2_X1 U704 ( .A1(n42), .A2(net20105), .ZN(n516) );
  OAI22_X1 U705 ( .A1(n467), .A2(net27193), .B1(net27165), .B2(n569), .ZN(n695) );
  INV_X1 U706 ( .A(n695), .ZN(n396) );
  OAI21_X1 U707 ( .B1(n396), .B2(n468), .A(n441), .ZN(n395) );
  AOI221_X1 U708 ( .B1(n817), .B2(n287), .C1(n297), .C2(n565), .A(n395), .ZN(
        n404) );
  NAND2_X1 U709 ( .A1(n396), .A2(n339), .ZN(n696) );
  INV_X1 U710 ( .A(n319), .ZN(n840) );
  OAI221_X1 U711 ( .B1(n841), .B2(net35616), .C1(n840), .C2(n329), .A(n497), 
        .ZN(n632) );
  INV_X1 U712 ( .A(n457), .ZN(n835) );
  OAI22_X1 U713 ( .A1(n397), .A2(n568), .B1(n835), .B2(n86), .ZN(n398) );
  AOI221_X1 U714 ( .B1(n151), .B2(n768), .C1(N99), .C2(net27187), .A(n398), 
        .ZN(n400) );
  AOI222_X1 U715 ( .A1(n146), .A2(n319), .B1(N67), .B2(net27185), .C1(n277), 
        .C2(n148), .ZN(n399) );
  NAND4_X1 U716 ( .A1(n400), .A2(n403), .A3(n404), .A4(n399), .ZN(RES[8]) );
  NAND2_X1 U717 ( .A1(n417), .A2(net27175), .ZN(n418) );
  OAI211_X1 U718 ( .C1(n36), .C2(net27195), .A(n339), .B(n418), .ZN(n710) );
  OAI21_X1 U719 ( .B1(n37), .B2(net27195), .A(n418), .ZN(n703) );
  AOI221_X1 U720 ( .B1(n479), .B2(n710), .C1(n478), .C2(n703), .A(n419), .ZN(
        n424) );
  INV_X1 U721 ( .A(n778), .ZN(n491) );
  INV_X1 U722 ( .A(n318), .ZN(n839) );
  OAI221_X1 U723 ( .B1(n840), .B2(net34835), .C1(n839), .C2(net34869), .A(n489), .ZN(n649) );
  INV_X1 U724 ( .A(n649), .ZN(n780) );
  OAI222_X1 U725 ( .A1(n491), .A2(net27193), .B1(net27165), .B2(n780), .C1(
        n420), .C2(net25237), .ZN(n711) );
  AOI222_X1 U726 ( .A1(n98), .A2(n498), .B1(n23), .B2(n711), .C1(n92), .C2(
        n577), .ZN(n423) );
  AOI222_X1 U727 ( .A1(N100), .A2(net27187), .B1(n189), .B2(n500), .C1(n768), 
        .C2(n136), .ZN(n422) );
  AOI222_X1 U728 ( .A1(n121), .A2(n317), .B1(N68), .B2(net27185), .C1(n280), 
        .C2(n127), .ZN(n421) );
  NAND4_X1 U729 ( .A1(n422), .A2(n423), .A3(n424), .A4(n421), .ZN(RES[9]) );
  NAND2_X1 U730 ( .A1(n134), .A2(net27175), .ZN(n431) );
  OAI21_X1 U731 ( .B1(net25143), .B2(net27195), .A(n431), .ZN(n727) );
  MUX2_X1 U732 ( .A(net27081), .B(net27113), .S(n56), .Z(n426) );
  NAND2_X1 U733 ( .A1(n426), .A2(net27103), .ZN(n430) );
  INV_X1 U734 ( .A(n315), .ZN(n819) );
  AOI21_X1 U735 ( .B1(net27095), .B2(n819), .A(net27105), .ZN(n428) );
  INV_X1 U736 ( .A(n56), .ZN(n427) );
  OAI21_X1 U737 ( .B1(n428), .B2(n427), .A(n441), .ZN(n429) );
  OAI211_X1 U738 ( .C1(net25150), .C2(net27195), .A(n339), .B(n431), .ZN(n728)
         );
  OAI211_X1 U739 ( .C1(n839), .C2(net34836), .A(n527), .B(n432), .ZN(n665) );
  INV_X1 U740 ( .A(n433), .ZN(n833) );
  OAI22_X1 U741 ( .A1(n28), .A2(n548), .B1(n833), .B2(n86), .ZN(n434) );
  AOI221_X1 U742 ( .B1(net27207), .B2(n665), .C1(n92), .C2(n593), .A(n434), 
        .ZN(n436) );
  AOI222_X1 U743 ( .A1(N69), .A2(net27183), .B1(n31), .B2(n175), .C1(N101), 
        .C2(net27189), .ZN(n435) );
  NAND4_X1 U744 ( .A1(n436), .A2(n437), .A3(n438), .A4(n435), .ZN(RES[10]) );
  NAND2_X1 U745 ( .A1(n237), .A2(net27175), .ZN(n446) );
  INV_X1 U746 ( .A(n446), .ZN(n742) );
  MUX2_X1 U747 ( .A(net27083), .B(net27113), .S(n223), .Z(n440) );
  NAND2_X1 U748 ( .A1(n440), .A2(net27103), .ZN(n445) );
  INV_X1 U749 ( .A(net34655), .ZN(net25527) );
  INV_X1 U750 ( .A(n223), .ZN(n443) );
  NAND3_X1 U751 ( .A1(n479), .A2(net34616), .A3(net27165), .ZN(n442) );
  NAND2_X1 U752 ( .A1(n442), .A2(n441), .ZN(n470) );
  INV_X1 U753 ( .A(n470), .ZN(n505) );
  OAI21_X1 U754 ( .B1(net25523), .B2(n443), .A(n505), .ZN(n444) );
  OAI21_X1 U755 ( .B1(net27193), .B2(net25114), .A(n446), .ZN(n745) );
  AOI22_X1 U756 ( .A1(net27123), .A2(n320), .B1(net27137), .B2(n185), .ZN(n447) );
  OAI211_X1 U757 ( .C1(n819), .C2(net34836), .A(n448), .B(n447), .ZN(net25238)
         );
  INV_X1 U758 ( .A(n449), .ZN(n832) );
  OAI22_X1 U759 ( .A1(n26), .A2(n548), .B1(n832), .B2(n86), .ZN(n450) );
  AOI222_X1 U760 ( .A1(N70), .A2(net27183), .B1(n31), .B2(n162), .C1(N102), 
        .C2(net27191), .ZN(n451) );
  NAND4_X1 U761 ( .A1(n452), .A2(n453), .A3(n455), .A4(n451), .ZN(RES[11]) );
  AOI222_X1 U762 ( .A1(n1), .A2(n457), .B1(n571), .B2(n456), .C1(n98), .C2(
        n572), .ZN(n477) );
  AOI222_X1 U763 ( .A1(N71), .A2(net27183), .B1(n92), .B2(n458), .C1(N103), 
        .C2(net27191), .ZN(n476) );
  INV_X1 U764 ( .A(n632), .ZN(n757) );
  AOI22_X1 U765 ( .A1(net27123), .A2(n317), .B1(n315), .B2(net27137), .ZN(n459) );
  NAND3_X1 U766 ( .A1(n461), .A2(n460), .A3(n459), .ZN(n697) );
  INV_X1 U767 ( .A(n697), .ZN(n756) );
  MUX2_X1 U768 ( .A(net27095), .B(net33647), .S(n255), .Z(n462) );
  OAI21_X1 U769 ( .B1(net27105), .B2(n462), .A(net28421), .ZN(n463) );
  OAI221_X1 U770 ( .B1(n757), .B2(n125), .C1(n756), .C2(net25503), .A(n463), 
        .ZN(n473) );
  INV_X1 U771 ( .A(net28422), .ZN(net25502) );
  INV_X1 U772 ( .A(n255), .ZN(n466) );
  NAND3_X1 U773 ( .A1(n23), .A2(net28241), .A3(n622), .ZN(n464) );
  OAI21_X1 U774 ( .B1(net25499), .B2(n466), .A(n464), .ZN(n472) );
  AOI211_X1 U775 ( .C1(n469), .C2(n468), .A(net27165), .B(n467), .ZN(n471) );
  NOR4_X1 U776 ( .A1(n473), .A2(n472), .A3(n471), .A4(n470), .ZN(n475) );
  NAND3_X1 U777 ( .A1(n477), .A2(n476), .A3(n475), .ZN(RES[12]) );
  OAI21_X1 U778 ( .B1(n314), .B2(net27081), .A(net27103), .ZN(n486) );
  NAND2_X1 U779 ( .A1(n479), .A2(net27175), .ZN(n510) );
  OAI21_X1 U780 ( .B1(n36), .B2(n510), .A(n505), .ZN(n481) );
  MUX2_X1 U781 ( .A(net27083), .B(net27113), .S(n276), .Z(n490) );
  NAND2_X1 U782 ( .A1(n490), .A2(net27103), .ZN(n493) );
  OAI22_X1 U783 ( .A1(n780), .A2(n125), .B1(n491), .B2(n516), .ZN(n492) );
  AOI221_X1 U784 ( .B1(n314), .B2(n493), .C1(n299), .C2(n777), .A(n492), .ZN(
        n503) );
  NAND3_X1 U785 ( .A1(n488), .A2(n495), .A3(n494), .ZN(n776) );
  INV_X1 U786 ( .A(n498), .ZN(n834) );
  OAI22_X1 U787 ( .A1(n55), .A2(n548), .B1(n834), .B2(n546), .ZN(n499) );
  AOI221_X1 U788 ( .B1(net27207), .B2(n776), .C1(n190), .C2(n577), .A(n499), 
        .ZN(n502) );
  AOI222_X1 U789 ( .A1(N72), .A2(net27183), .B1(n92), .B2(n500), .C1(N104), 
        .C2(net27191), .ZN(n501) );
  NAND4_X1 U790 ( .A1(n502), .A2(n503), .A3(n504), .A4(n501), .ZN(RES[13]) );
  OAI21_X1 U791 ( .B1(n326), .B2(net27081), .A(net27103), .ZN(n514) );
  OAI21_X1 U792 ( .B1(net25150), .B2(n510), .A(n505), .ZN(n511) );
  MUX2_X1 U793 ( .A(net27083), .B(net27113), .S(n262), .Z(n515) );
  NAND2_X1 U794 ( .A1(n515), .A2(net27103), .ZN(n519) );
  INV_X1 U795 ( .A(n665), .ZN(n803) );
  INV_X1 U796 ( .A(n801), .ZN(n717) );
  OAI22_X1 U797 ( .A1(n803), .A2(n126), .B1(n717), .B2(n516), .ZN(n518) );
  AOI221_X1 U798 ( .B1(n326), .B2(n519), .C1(n299), .C2(n800), .A(n518), .ZN(
        n532) );
  NAND3_X1 U799 ( .A1(n474), .A2(n525), .A3(n524), .ZN(n799) );
  OAI22_X1 U800 ( .A1(n95), .A2(n548), .B1(n833), .B2(n546), .ZN(n526) );
  AOI221_X1 U801 ( .B1(net27207), .B2(n799), .C1(n190), .C2(n593), .A(n526), 
        .ZN(n531) );
  NAND4_X1 U802 ( .A1(n531), .A2(n532), .A3(n533), .A4(n530), .ZN(RES[14]) );
  MUX2_X1 U803 ( .A(net27083), .B(net27113), .S(n243), .Z(n534) );
  NAND2_X1 U804 ( .A1(n534), .A2(net27103), .ZN(net25442) );
  INV_X1 U805 ( .A(n104), .ZN(net25448) );
  AOI21_X1 U806 ( .B1(net27095), .B2(net25448), .A(net27105), .ZN(n537) );
  INV_X1 U807 ( .A(n243), .ZN(n536) );
  NAND2_X1 U808 ( .A1(n301), .A2(n535), .ZN(n733) );
  OAI21_X1 U809 ( .B1(n537), .B2(n536), .A(n733), .ZN(net25443) );
  AOI222_X1 U810 ( .A1(n296), .A2(net25238), .B1(n299), .B2(net25131), .C1(
        n743), .C2(net25130), .ZN(n556) );
  NAND3_X1 U811 ( .A1(n465), .A2(n539), .A3(n538), .ZN(net25132) );
  OAI22_X1 U812 ( .A1(n607), .A2(n548), .B1(n832), .B2(n546), .ZN(n551) );
  AOI221_X1 U813 ( .B1(n116), .B2(net25132), .C1(n190), .C2(n606), .A(n551), 
        .ZN(n555) );
  NAND4_X1 U814 ( .A1(n554), .A2(n556), .A3(net25429), .A4(n555), .ZN(RES[15])
         );
  NAND2_X1 U815 ( .A1(net33657), .A2(n58), .ZN(n621) );
  INV_X1 U816 ( .A(n621), .ZN(n736) );
  MUX2_X1 U817 ( .A(net27083), .B(net27113), .S(n2), .Z(n557) );
  NAND2_X1 U818 ( .A1(n557), .A2(net27103), .ZN(n562) );
  INV_X1 U819 ( .A(n226), .ZN(n558) );
  AOI21_X1 U820 ( .B1(net27095), .B2(n558), .A(net27105), .ZN(n560) );
  INV_X1 U821 ( .A(B[16]), .ZN(n559) );
  OAI21_X1 U822 ( .B1(n560), .B2(n559), .A(n733), .ZN(n561) );
  AOI221_X1 U823 ( .B1(n298), .B2(n817), .C1(n226), .C2(n562), .A(n561), .ZN(
        n576) );
  NAND3_X1 U824 ( .A1(n454), .A2(n564), .A3(n563), .ZN(n750) );
  AOI222_X1 U825 ( .A1(net27205), .A2(n750), .B1(n299), .B2(n565), .C1(n743), 
        .C2(n632), .ZN(n575) );
  OAI22_X1 U826 ( .A1(n569), .A2(n568), .B1(n567), .B2(n86), .ZN(n570) );
  AOI221_X1 U827 ( .B1(n297), .B2(n697), .C1(n571), .C2(n767), .A(n570), .ZN(
        n574) );
  AOI222_X1 U828 ( .A1(N75), .A2(net27183), .B1(n768), .B2(n572), .C1(N107), 
        .C2(net27191), .ZN(n573) );
  NAND4_X1 U829 ( .A1(n573), .A2(n576), .A3(n574), .A4(n575), .ZN(RES[16]) );
  OAI222_X1 U830 ( .A1(n55), .A2(net25237), .B1(net27167), .B2(n256), .C1(n244), .C2(net27195), .ZN(n578) );
  INV_X1 U831 ( .A(n578), .ZN(n579) );
  OAI21_X1 U832 ( .B1(n281), .B2(net27081), .A(net27103), .ZN(n580) );
  INV_X1 U833 ( .A(n733), .ZN(n718) );
  AOI221_X1 U834 ( .B1(n298), .B2(n777), .C1(n103), .C2(n580), .A(n718), .ZN(
        n592) );
  MUX2_X1 U835 ( .A(net27083), .B(net27113), .S(n103), .Z(n584) );
  INV_X1 U836 ( .A(n281), .ZN(n583) );
  AOI21_X1 U837 ( .B1(n584), .B2(net27101), .A(n583), .ZN(n585) );
  AOI22_X1 U838 ( .A1(n326), .A2(net27123), .B1(net27527), .B2(net27131), .ZN(
        n586) );
  NAND3_X1 U839 ( .A1(n588), .A2(n587), .A3(n586), .ZN(n771) );
  AOI222_X1 U840 ( .A1(n286), .A2(n649), .B1(net27209), .B2(n771), .C1(n299), 
        .C2(n778), .ZN(n590) );
  NAND4_X1 U841 ( .A1(n592), .A2(n591), .A3(n590), .A4(n589), .ZN(RES[17]) );
  OAI21_X1 U842 ( .B1(n249), .B2(net27081), .A(net27103), .ZN(n595) );
  AOI221_X1 U843 ( .B1(n298), .B2(n800), .C1(n99), .C2(n595), .A(n718), .ZN(
        n605) );
  AOI22_X1 U844 ( .A1(net27527), .A2(net27121), .B1(n226), .B2(net27137), .ZN(
        n596) );
  NAND3_X1 U845 ( .A1(n598), .A2(n597), .A3(n596), .ZN(n794) );
  MUX2_X1 U846 ( .A(net27083), .B(net27113), .S(n99), .Z(n600) );
  INV_X1 U847 ( .A(A[18]), .ZN(n599) );
  AOI21_X1 U848 ( .B1(n600), .B2(net27101), .A(n599), .ZN(n601) );
  AOI221_X1 U849 ( .B1(n292), .B2(n25), .C1(n116), .C2(n794), .A(n601), .ZN(
        n604) );
  AOI222_X1 U850 ( .A1(n287), .A2(n665), .B1(n788), .B2(n266), .C1(n299), .C2(
        n801), .ZN(n603) );
  AOI222_X1 U851 ( .A1(N77), .A2(net27183), .B1(n297), .B2(n799), .C1(N109), 
        .C2(net27191), .ZN(n602) );
  NAND4_X1 U852 ( .A1(n602), .A2(n604), .A3(n603), .A4(n605), .ZN(RES[18]) );
  OAI222_X1 U853 ( .A1(n22), .A2(net25237), .B1(net27167), .B2(n240), .C1(n108), .C2(net27195), .ZN(n608) );
  INV_X1 U854 ( .A(n608), .ZN(n609) );
  NAND2_X1 U855 ( .A1(n609), .A2(n378), .ZN(n207) );
  NAND2_X1 U856 ( .A1(n609), .A2(net25366), .ZN(n205) );
  OAI21_X1 U857 ( .B1(n231), .B2(net27081), .A(net27103), .ZN(n610) );
  AOI22_X1 U858 ( .A1(n226), .A2(net27121), .B1(n281), .B2(net27137), .ZN(n611) );
  NAND3_X1 U859 ( .A1(n613), .A2(n612), .A3(n611), .ZN(net25137) );
  MUX2_X1 U860 ( .A(net27083), .B(net27113), .S(n199), .Z(n615) );
  INV_X1 U861 ( .A(A[19]), .ZN(n614) );
  AOI21_X1 U862 ( .B1(n615), .B2(net27101), .A(n614), .ZN(n616) );
  AOI221_X1 U863 ( .B1(n293), .B2(n120), .C1(n116), .C2(net25137), .A(n616), 
        .ZN(n619) );
  AOI222_X1 U864 ( .A1(n286), .A2(net25238), .B1(n788), .B2(n205), .C1(n299), 
        .C2(net25130), .ZN(n618) );
  NAND4_X1 U865 ( .A1(n617), .A2(n619), .A3(n618), .A4(n620), .ZN(RES[19]) );
  OAI21_X1 U866 ( .B1(n283), .B2(net27081), .A(net27103), .ZN(n624) );
  NOR2_X1 U867 ( .A1(net28241), .A2(n621), .ZN(n623) );
  AOI221_X1 U868 ( .B1(B[20]), .B2(n624), .C1(n623), .C2(n622), .A(n718), .ZN(
        n637) );
  AOI22_X1 U869 ( .A1(n281), .A2(net27121), .B1(n249), .B2(net27131), .ZN(n625) );
  NAND3_X1 U870 ( .A1(n627), .A2(n626), .A3(n625), .ZN(n751) );
  MUX2_X1 U871 ( .A(net27083), .B(net27113), .S(B[20]), .Z(n629) );
  INV_X1 U872 ( .A(n283), .ZN(n628) );
  AOI21_X1 U873 ( .B1(n629), .B2(net27101), .A(n628), .ZN(n630) );
  AOI221_X1 U874 ( .B1(n116), .B2(n751), .C1(n788), .C2(n631), .A(n630), .ZN(
        n636) );
  AOI222_X1 U875 ( .A1(n287), .A2(n697), .B1(n293), .B2(n633), .C1(n299), .C2(
        n632), .ZN(n635) );
  AOI222_X1 U876 ( .A1(N79), .A2(net27181), .B1(n296), .B2(n750), .C1(N111), 
        .C2(net27191), .ZN(n634) );
  NAND4_X1 U877 ( .A1(n636), .A2(n637), .A3(n635), .A4(n634), .ZN(RES[20]) );
  INV_X1 U878 ( .A(n257), .ZN(n644) );
  AOI21_X1 U879 ( .B1(net27095), .B2(n644), .A(net27105), .ZN(n639) );
  INV_X1 U880 ( .A(n194), .ZN(n638) );
  OAI21_X1 U881 ( .B1(n639), .B2(n638), .A(n733), .ZN(n640) );
  AOI221_X1 U882 ( .B1(n300), .B2(n777), .C1(n298), .C2(n778), .A(n640), .ZN(
        n653) );
  AOI22_X1 U883 ( .A1(n249), .A2(net35005), .B1(n231), .B2(net27131), .ZN(n641) );
  NAND3_X1 U884 ( .A1(n643), .A2(n642), .A3(n641), .ZN(n772) );
  MUX2_X1 U885 ( .A(net27083), .B(net27113), .S(n194), .Z(n645) );
  AOI21_X1 U886 ( .B1(n645), .B2(net27101), .A(n644), .ZN(n646) );
  AOI221_X1 U887 ( .B1(n293), .B2(n647), .C1(net27205), .C2(n772), .A(n646), 
        .ZN(n652) );
  AOI222_X1 U888 ( .A1(n299), .A2(n649), .B1(n788), .B2(n648), .C1(n744), .C2(
        n771), .ZN(n651) );
  AOI222_X1 U889 ( .A1(N80), .A2(net27181), .B1(n287), .B2(n776), .C1(N112), 
        .C2(net27189), .ZN(n650) );
  NAND4_X1 U890 ( .A1(n651), .A2(n652), .A3(n650), .A4(n653), .ZN(RES[21]) );
  INV_X1 U891 ( .A(n6), .ZN(n660) );
  AOI21_X1 U892 ( .B1(net27095), .B2(n660), .A(net27105), .ZN(n655) );
  INV_X1 U893 ( .A(n32), .ZN(n654) );
  OAI21_X1 U894 ( .B1(n655), .B2(n654), .A(n733), .ZN(n656) );
  AOI221_X1 U895 ( .B1(n300), .B2(n800), .C1(n298), .C2(n801), .A(n656), .ZN(
        n669) );
  AOI22_X1 U896 ( .A1(n231), .A2(net27121), .B1(n283), .B2(net27137), .ZN(n657) );
  NAND3_X1 U897 ( .A1(n659), .A2(n658), .A3(n657), .ZN(n795) );
  MUX2_X1 U898 ( .A(net27083), .B(net27113), .S(n213), .Z(n661) );
  AOI21_X1 U899 ( .B1(n661), .B2(net27101), .A(n660), .ZN(n662) );
  AOI221_X1 U900 ( .B1(n297), .B2(n794), .C1(n116), .C2(n795), .A(n662), .ZN(
        n668) );
  AOI222_X1 U901 ( .A1(n299), .A2(n665), .B1(n292), .B2(n664), .C1(n788), .C2(
        n663), .ZN(n667) );
  AOI222_X1 U902 ( .A1(N81), .A2(net27181), .B1(n286), .B2(n799), .C1(N113), 
        .C2(net27189), .ZN(n666) );
  NAND4_X1 U903 ( .A1(n666), .A2(n668), .A3(n667), .A4(n669), .ZN(RES[22]) );
  INV_X1 U904 ( .A(A[23]), .ZN(n676) );
  AOI21_X1 U905 ( .B1(net27095), .B2(n676), .A(net27105), .ZN(n671) );
  INV_X1 U906 ( .A(B[23]), .ZN(n670) );
  OAI21_X1 U907 ( .B1(n671), .B2(n670), .A(n733), .ZN(n672) );
  AOI221_X1 U908 ( .B1(n300), .B2(net25131), .C1(n298), .C2(net25130), .A(n672), .ZN(n684) );
  AOI22_X1 U909 ( .A1(n283), .A2(net27121), .B1(n257), .B2(net27137), .ZN(n673) );
  NAND3_X1 U910 ( .A1(n675), .A2(n674), .A3(n673), .ZN(net25136) );
  MUX2_X1 U911 ( .A(net27083), .B(net27113), .S(B[23]), .Z(n677) );
  AOI21_X1 U912 ( .B1(n677), .B2(net27101), .A(n676), .ZN(n678) );
  AOI221_X1 U913 ( .B1(n297), .B2(net25137), .C1(net27205), .C2(net25136), .A(
        n678), .ZN(n683) );
  AOI222_X1 U914 ( .A1(n299), .A2(net25238), .B1(n293), .B2(n680), .C1(n788), 
        .C2(n679), .ZN(n682) );
  NAND4_X1 U915 ( .A1(n681), .A2(n683), .A3(n682), .A4(n684), .ZN(RES[23]) );
  OAI222_X1 U916 ( .A1(n686), .A2(net27193), .B1(net27165), .B2(n757), .C1(
        net25237), .C2(n685), .ZN(n688) );
  OAI21_X1 U917 ( .B1(A[24]), .B2(net27081), .A(net27101), .ZN(n687) );
  AOI221_X1 U918 ( .B1(n736), .B2(n688), .C1(n5), .C2(n687), .A(n718), .ZN(
        n701) );
  AOI22_X1 U919 ( .A1(n257), .A2(net27121), .B1(n6), .B2(net27131), .ZN(n689)
         );
  NAND3_X1 U920 ( .A1(n691), .A2(n690), .A3(n689), .ZN(n752) );
  MUX2_X1 U921 ( .A(net27083), .B(net27113), .S(n5), .Z(n693) );
  INV_X1 U922 ( .A(A[24]), .ZN(n692) );
  AOI21_X1 U923 ( .B1(n693), .B2(net27101), .A(n692), .ZN(n694) );
  AOI221_X1 U924 ( .B1(net27209), .B2(n752), .C1(n788), .C2(n695), .A(n694), 
        .ZN(n700) );
  AOI222_X1 U925 ( .A1(n299), .A2(n697), .B1(n744), .B2(n751), .C1(n293), .C2(
        n696), .ZN(n699) );
  AOI222_X1 U926 ( .A1(N83), .A2(net27181), .B1(n286), .B2(n750), .C1(N115), 
        .C2(net27189), .ZN(n698) );
  NAND4_X1 U927 ( .A1(n698), .A2(n700), .A3(n699), .A4(n701), .ZN(RES[24]) );
  OAI21_X1 U928 ( .B1(n242), .B2(net27081), .A(net27103), .ZN(n702) );
  AOI221_X1 U929 ( .B1(n788), .B2(n703), .C1(B[25]), .C2(n702), .A(n718), .ZN(
        n715) );
  AOI22_X1 U930 ( .A1(n6), .A2(net35006), .B1(n188), .B2(net27137), .ZN(n704)
         );
  NAND3_X1 U931 ( .A1(n706), .A2(n705), .A3(n704), .ZN(n773) );
  MUX2_X1 U932 ( .A(net27083), .B(net27113), .S(B[25]), .Z(n708) );
  INV_X1 U933 ( .A(n242), .ZN(n707) );
  AOI21_X1 U934 ( .B1(n708), .B2(net27101), .A(n707), .ZN(n709) );
  AOI221_X1 U935 ( .B1(n296), .B2(n772), .C1(net27205), .C2(n773), .A(n709), 
        .ZN(n714) );
  AOI222_X1 U936 ( .A1(n736), .A2(n711), .B1(n292), .B2(n710), .C1(n743), .C2(
        n771), .ZN(n713) );
  AOI222_X1 U937 ( .A1(N84), .A2(net27181), .B1(n299), .B2(n776), .C1(N116), 
        .C2(net27189), .ZN(n712) );
  NAND4_X1 U938 ( .A1(n712), .A2(n714), .A3(n713), .A4(n715), .ZN(RES[25]) );
  OAI222_X1 U939 ( .A1(n717), .A2(net27193), .B1(net27165), .B2(n803), .C1(
        n716), .C2(net25237), .ZN(n720) );
  OAI21_X1 U940 ( .B1(A[26]), .B2(net27081), .A(net27101), .ZN(n719) );
  AOI221_X1 U941 ( .B1(n736), .B2(n720), .C1(n216), .C2(n719), .A(n718), .ZN(
        n732) );
  AOI22_X1 U942 ( .A1(n188), .A2(net27121), .B1(A[24]), .B2(net27131), .ZN(
        n721) );
  NAND3_X1 U943 ( .A1(n137), .A2(n722), .A3(n721), .ZN(n796) );
  MUX2_X1 U944 ( .A(net27083), .B(net27113), .S(n216), .Z(n725) );
  INV_X1 U945 ( .A(A[26]), .ZN(n724) );
  AOI21_X1 U946 ( .B1(n725), .B2(net27101), .A(n724), .ZN(n726) );
  AOI221_X1 U947 ( .B1(n116), .B2(n796), .C1(n788), .C2(n727), .A(n726), .ZN(
        n731) );
  AOI222_X1 U948 ( .A1(N85), .A2(net27181), .B1(n299), .B2(n799), .C1(N117), 
        .C2(net27189), .ZN(n729) );
  NAND4_X1 U949 ( .A1(n729), .A2(n732), .A3(n730), .A4(n731), .ZN(RES[26]) );
  OAI21_X1 U950 ( .B1(A[27]), .B2(net27081), .A(net27101), .ZN(n735) );
  NAND2_X1 U951 ( .A1(n734), .A2(n733), .ZN(n761) );
  AOI22_X1 U952 ( .A1(A[24]), .A2(net27121), .B1(n242), .B2(net27131), .ZN(
        n737) );
  NAND3_X1 U953 ( .A1(n739), .A2(n738), .A3(n737), .ZN(net25138) );
  MUX2_X1 U954 ( .A(net27083), .B(net27113), .S(n30), .Z(n740) );
  AOI21_X1 U955 ( .B1(n740), .B2(net27101), .A(n818), .ZN(n741) );
  AOI221_X1 U956 ( .B1(n116), .B2(net25138), .C1(n742), .C2(n292), .A(n741), 
        .ZN(n748) );
  AOI222_X1 U957 ( .A1(n788), .A2(n745), .B1(n296), .B2(net25136), .C1(n743), 
        .C2(net25137), .ZN(n747) );
  NAND4_X1 U958 ( .A1(n746), .A2(n748), .A3(n747), .A4(n749), .ZN(RES[27]) );
  INV_X1 U959 ( .A(n750), .ZN(n754) );
  AOI22_X1 U960 ( .A1(net27201), .A2(n752), .B1(net20105), .B2(n751), .ZN(n753) );
  OAI221_X1 U961 ( .B1(net18434), .B2(n754), .C1(n295), .C2(net27165), .A(n753), .ZN(n759) );
  OAI222_X1 U962 ( .A1(n757), .A2(net27193), .B1(net27165), .B2(n756), .C1(
        net20024), .C2(n755), .ZN(n758) );
  MUX2_X1 U963 ( .A(n759), .B(n758), .S(net38433), .Z(n766) );
  MUX2_X1 U964 ( .A(net27083), .B(net27113), .S(n248), .Z(n760) );
  NAND2_X1 U965 ( .A1(n760), .A2(net27103), .ZN(n765) );
  AOI21_X1 U966 ( .B1(net27095), .B2(net20044), .A(net27105), .ZN(n763) );
  INV_X1 U967 ( .A(n248), .ZN(n762) );
  OAI21_X1 U968 ( .B1(n763), .B2(n762), .A(n128), .ZN(n764) );
  AOI222_X1 U969 ( .A1(N87), .A2(net27181), .B1(n31), .B2(n767), .C1(N119), 
        .C2(net27189), .ZN(n769) );
  NAND2_X1 U970 ( .A1(n770), .A2(n769), .ZN(RES[28]) );
  OAI21_X1 U971 ( .B1(n181), .B2(net27081), .A(net27103), .ZN(n787) );
  INV_X1 U972 ( .A(n771), .ZN(n775) );
  AOI22_X1 U973 ( .A1(net27201), .A2(n773), .B1(net20105), .B2(n772), .ZN(n774) );
  OAI221_X1 U974 ( .B1(net18434), .B2(n775), .C1(n279), .C2(net27165), .A(n774), .ZN(n783) );
  INV_X1 U975 ( .A(n776), .ZN(n781) );
  AOI22_X1 U976 ( .A1(net20105), .A2(n778), .B1(n777), .B2(n232), .ZN(n779) );
  OAI221_X1 U977 ( .B1(net27165), .B2(n781), .C1(n780), .C2(net27195), .A(n779), .ZN(n782) );
  MUX2_X1 U978 ( .A(n783), .B(n782), .S(net38433), .Z(n786) );
  NAND2_X1 U979 ( .A1(n292), .A2(net27175), .ZN(n807) );
  OAI21_X1 U980 ( .B1(n36), .B2(n807), .A(n246), .ZN(n785) );
  NAND2_X1 U981 ( .A1(n788), .A2(net27175), .ZN(net25113) );
  MUX2_X1 U982 ( .A(net27095), .B(net33647), .S(n236), .Z(n789) );
  OAI21_X1 U983 ( .B1(net27105), .B2(n789), .A(n181), .ZN(n790) );
  OAI21_X1 U984 ( .B1(n37), .B2(net25113), .A(n790), .ZN(n791) );
  NAND2_X1 U985 ( .A1(n792), .A2(n793), .ZN(RES[29]) );
  OAI21_X1 U986 ( .B1(n113), .B2(net27081), .A(net27101), .ZN(n810) );
  INV_X1 U987 ( .A(n794), .ZN(n798) );
  AOI22_X1 U988 ( .A1(net27203), .A2(n796), .B1(net20105), .B2(n795), .ZN(n797) );
  OAI221_X1 U989 ( .B1(net18434), .B2(n798), .C1(n247), .C2(net27165), .A(n797), .ZN(n806) );
  INV_X1 U990 ( .A(n799), .ZN(n804) );
  AOI22_X1 U991 ( .A1(net20105), .A2(n801), .B1(n800), .B2(n232), .ZN(n802) );
  OAI221_X1 U992 ( .B1(net27165), .B2(n804), .C1(n803), .C2(net27195), .A(n802), .ZN(n805) );
  MUX2_X1 U993 ( .A(n806), .B(n805), .S(net38433), .Z(n809) );
  OAI21_X1 U994 ( .B1(net25150), .B2(n807), .A(n128), .ZN(n808) );
  OAI21_X1 U995 ( .B1(net27105), .B2(net25146), .A(n113), .ZN(n811) );
  OAI21_X1 U996 ( .B1(net25143), .B2(net25113), .A(n811), .ZN(n812) );
  NAND2_X1 U997 ( .A1(n813), .A2(n814), .ZN(RES[30]) );
  MUX2_X1 U998 ( .A(net27081), .B(net27113), .S(B[31]), .Z(n815) );
  NAND3_X1 U999 ( .A1(n239), .A2(net27103), .A3(n815), .ZN(n816) );
  INV_X1 U1000 ( .A(n412), .ZN(n838) );
  INV_X1 U1001 ( .A(n407), .ZN(n831) );
  INV_X1 U1002 ( .A(n269), .ZN(n837) );
  INV_X1 U1003 ( .A(n265), .ZN(n830) );
  INV_X1 U1004 ( .A(net25112), .ZN(n254) );
  INV_X1 U1005 ( .A(n211), .ZN(n836) );
  INV_X1 U1006 ( .A(n204), .ZN(n829) );
  OR3_X1 U1007 ( .A1(B[15]), .A2(B[14]), .A3(B[13]), .ZN(n821) );
  NOR4_X1 U1008 ( .A1(n821), .A2(n56), .A3(n238), .A4(n223), .ZN(n828) );
  NOR4_X1 U1009 ( .A1(n823), .A2(B[23]), .A3(B[25]), .A4(B[24]), .ZN(n826) );
endmodule


module REG_PIPO_6_00_00_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [5:0] DIN;
  output [5:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21;

  DFFR_X1 \reg_mem_reg[5]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[5]) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n14), .ZN(n20) );
  INV_X1 U3 ( .A(n21), .ZN(n13) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n20), .B1(n14), .B2(DOUT[0]), .ZN(n21) );
  INV_X1 U5 ( .A(n19), .ZN(n12) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n20), .B1(n14), .B2(DOUT[1]), .ZN(n19) );
  INV_X1 U7 ( .A(n18), .ZN(n11) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n20), .B1(n14), .B2(DOUT[2]), .ZN(n18) );
  INV_X1 U9 ( .A(n17), .ZN(n10) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n20), .B1(n14), .B2(DOUT[3]), .ZN(n17) );
  INV_X1 U11 ( .A(n16), .ZN(n9) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n20), .B1(n14), .B2(DOUT[4]), .ZN(n16) );
  INV_X1 U13 ( .A(n15), .ZN(n3) );
  AOI22_X1 U14 ( .A1(DIN[5]), .A2(n20), .B1(n14), .B2(DOUT[5]), .ZN(n15) );
  INV_X1 U15 ( .A(EN), .ZN(n14) );
endmodule


module REG_PIPO_32_00000000_00000000_6 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n3) );
  BUF_X1 U4 ( .A(n169), .Z(n2) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U29 ( .A(DIN[21]), .ZN(n19) );
  OAI22_X1 U30 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U31 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U32 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U33 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U34 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U35 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U36 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U37 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U38 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U39 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U40 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U41 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U42 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U43 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U44 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U45 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U46 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U47 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U48 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U49 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U50 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U51 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U52 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U53 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U54 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U55 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U56 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U57 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U58 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U59 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U60 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U61 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U62 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U63 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U64 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U65 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U66 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U67 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U68 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U69 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U70 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U71 ( .A(DIN[20]), .ZN(n20) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_32_00000000_00000000_5 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n98, net25088, net34508, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175;

  DFFR_X1 \reg_mem_reg[30]  ( .D(n113), .CK(CLK), .RN(n17), .Q(DOUT[30]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n114), .CK(CLK), .RN(n17), .Q(DOUT[29]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n115), .CK(CLK), .RN(n17), .Q(DOUT[28]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n116), .CK(CLK), .RN(n17), .Q(DOUT[27]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n117), .CK(CLK), .RN(n17), .Q(DOUT[26]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n118), .CK(CLK), .RN(n17), .Q(DOUT[25]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n119), .CK(CLK), .RN(n17), .Q(DOUT[24]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n120), .CK(CLK), .RN(n17), .Q(DOUT[23]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n121), .CK(CLK), .RN(n17), .Q(DOUT[22]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n122), .CK(CLK), .RN(n16), .Q(DOUT[21]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n123), .CK(CLK), .RN(n16), .Q(DOUT[20]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n124), .CK(CLK), .RN(n16), .Q(DOUT[19]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n125), .CK(CLK), .RN(n16), .Q(DOUT[18]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n126), .CK(CLK), .RN(n16), .Q(DOUT[17]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n127), .CK(CLK), .RN(n16), .Q(DOUT[16]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n128), .CK(CLK), .RN(n16), .Q(DOUT[15]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n129), .CK(CLK), .RN(n16), .Q(DOUT[14]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n130), .CK(CLK), .RN(n16), .Q(DOUT[13]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n131), .CK(CLK), .RN(n16), .Q(DOUT[12]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n132), .CK(CLK), .RN(n16), .Q(DOUT[11]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n133), .CK(CLK), .RN(n15), .Q(DOUT[10]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n134), .CK(CLK), .RN(n15), .Q(DOUT[9]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n135), .CK(CLK), .RN(n15), .Q(DOUT[8]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n136), .CK(CLK), .RN(n15), .Q(DOUT[7]), .QN(
        n168) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n137), .CK(CLK), .RN(n15), .Q(DOUT[6]), .QN(
        n169) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n138), .CK(CLK), .RN(n15), .Q(DOUT[5]), .QN(
        n170) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n139), .CK(CLK), .RN(n15), .Q(DOUT[4]), .QN(
        n171) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n140), .CK(CLK), .RN(n15), .Q(DOUT[3]), .QN(
        n172) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n141), .CK(CLK), .RN(n15), .Q(DOUT[2]), .QN(
        n173) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n142), .CK(CLK), .RN(n15), .Q(DOUT[1]), .QN(
        n174) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n143), .CK(CLK), .RN(n15), .Q(DOUT[0]), .QN(
        n175) );
  DFFR_X1 \reg_mem_reg[31]  ( .D(n98), .CK(CLK), .RN(n17), .Q(DOUT[31]), .QN(
        n144) );
  OR2_X1 U2 ( .A1(n145), .A2(EN), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n2), .A2(n103), .ZN(n113) );
  OR2_X1 U4 ( .A1(n151), .A2(EN), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n33), .A2(n3), .ZN(n119) );
  OR2_X1 U6 ( .A1(n161), .A2(EN), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n23), .A2(n4), .ZN(n129) );
  OR2_X1 U8 ( .A1(n155), .A2(EN), .ZN(n5) );
  NAND2_X1 U9 ( .A1(n29), .A2(n5), .ZN(n123) );
  OR2_X1 U10 ( .A1(n157), .A2(EN), .ZN(n6) );
  NAND2_X1 U11 ( .A1(n6), .A2(n27), .ZN(n125) );
  OR2_X1 U12 ( .A1(n153), .A2(EN), .ZN(n7) );
  NAND2_X1 U13 ( .A1(n31), .A2(n7), .ZN(n121) );
  NAND2_X1 U14 ( .A1(DIN[31]), .A2(net25088), .ZN(n8) );
  NAND2_X1 U15 ( .A1(n8), .A2(net34508), .ZN(n98) );
  INV_X1 U16 ( .A(n1), .ZN(net25088) );
  OR2_X1 U17 ( .A1(INIT), .A2(n9), .ZN(n1) );
  INV_X1 U18 ( .A(EN), .ZN(n9) );
  OR2_X1 U19 ( .A1(n175), .A2(EN), .ZN(n10) );
  NAND2_X1 U20 ( .A1(n18), .A2(n10), .ZN(n143) );
  OR2_X1 U21 ( .A1(n160), .A2(EN), .ZN(n11) );
  NAND2_X1 U22 ( .A1(n24), .A2(n11), .ZN(n128) );
  OR2_X1 U23 ( .A1(n146), .A2(EN), .ZN(n12) );
  NAND2_X1 U24 ( .A1(n102), .A2(n12), .ZN(n114) );
  OR2_X1 U25 ( .A1(n152), .A2(EN), .ZN(n13) );
  NAND2_X1 U26 ( .A1(n32), .A2(n13), .ZN(n120) );
  OR2_X1 U27 ( .A1(n148), .A2(EN), .ZN(n14) );
  NAND2_X1 U28 ( .A1(n100), .A2(n14), .ZN(n116) );
  OR2_X1 U29 ( .A1(n144), .A2(EN), .ZN(net34508) );
  BUF_X1 U30 ( .A(RST_AN), .Z(n15) );
  BUF_X1 U31 ( .A(RST_AN), .Z(n16) );
  BUF_X1 U32 ( .A(RST_AN), .Z(n17) );
  INV_X1 U33 ( .A(DIN[1]), .ZN(n112) );
  OAI22_X1 U34 ( .A1(n169), .A2(EN), .B1(n107), .B2(n1), .ZN(n137) );
  INV_X1 U35 ( .A(DIN[6]), .ZN(n107) );
  OAI22_X1 U36 ( .A1(n170), .A2(EN), .B1(n108), .B2(n1), .ZN(n138) );
  INV_X1 U37 ( .A(DIN[5]), .ZN(n108) );
  OAI22_X1 U38 ( .A1(n168), .A2(EN), .B1(n106), .B2(n1), .ZN(n136) );
  INV_X1 U39 ( .A(DIN[7]), .ZN(n106) );
  OAI22_X1 U40 ( .A1(n166), .A2(EN), .B1(n104), .B2(n1), .ZN(n134) );
  INV_X1 U41 ( .A(DIN[9]), .ZN(n104) );
  OAI22_X1 U42 ( .A1(n173), .A2(EN), .B1(n111), .B2(n1), .ZN(n141) );
  INV_X1 U43 ( .A(DIN[2]), .ZN(n111) );
  OAI22_X1 U44 ( .A1(n167), .A2(EN), .B1(n1), .B2(n105), .ZN(n135) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n105) );
  OAI22_X1 U46 ( .A1(n172), .A2(EN), .B1(n110), .B2(n1), .ZN(n140) );
  INV_X1 U47 ( .A(DIN[3]), .ZN(n110) );
  OAI22_X1 U48 ( .A1(n171), .A2(EN), .B1(n109), .B2(n1), .ZN(n139) );
  INV_X1 U49 ( .A(DIN[4]), .ZN(n109) );
  OAI22_X1 U50 ( .A1(n174), .A2(EN), .B1(n112), .B2(n1), .ZN(n142) );
  NAND2_X1 U51 ( .A1(DIN[0]), .A2(net25088), .ZN(n18) );
  NAND2_X1 U52 ( .A1(DIN[10]), .A2(net25088), .ZN(n19) );
  OAI21_X1 U53 ( .B1(n165), .B2(EN), .A(n19), .ZN(n133) );
  NAND2_X1 U54 ( .A1(DIN[11]), .A2(net25088), .ZN(n20) );
  OAI21_X1 U55 ( .B1(n164), .B2(EN), .A(n20), .ZN(n132) );
  NAND2_X1 U56 ( .A1(DIN[12]), .A2(net25088), .ZN(n21) );
  OAI21_X1 U57 ( .B1(n163), .B2(EN), .A(n21), .ZN(n131) );
  NAND2_X1 U58 ( .A1(DIN[13]), .A2(net25088), .ZN(n22) );
  OAI21_X1 U59 ( .B1(n162), .B2(EN), .A(n22), .ZN(n130) );
  NAND2_X1 U60 ( .A1(DIN[14]), .A2(net25088), .ZN(n23) );
  NAND2_X1 U61 ( .A1(DIN[15]), .A2(net25088), .ZN(n24) );
  NAND2_X1 U62 ( .A1(DIN[16]), .A2(net25088), .ZN(n25) );
  OAI21_X1 U63 ( .B1(n159), .B2(EN), .A(n25), .ZN(n127) );
  NAND2_X1 U64 ( .A1(DIN[17]), .A2(net25088), .ZN(n26) );
  OAI21_X1 U65 ( .B1(n158), .B2(EN), .A(n26), .ZN(n126) );
  NAND2_X1 U66 ( .A1(DIN[18]), .A2(net25088), .ZN(n27) );
  NAND2_X1 U67 ( .A1(DIN[19]), .A2(net25088), .ZN(n28) );
  OAI21_X1 U68 ( .B1(n156), .B2(EN), .A(n28), .ZN(n124) );
  NAND2_X1 U69 ( .A1(DIN[20]), .A2(net25088), .ZN(n29) );
  NAND2_X1 U70 ( .A1(DIN[21]), .A2(net25088), .ZN(n30) );
  OAI21_X1 U71 ( .B1(n154), .B2(EN), .A(n30), .ZN(n122) );
  NAND2_X1 U72 ( .A1(DIN[22]), .A2(net25088), .ZN(n31) );
  NAND2_X1 U73 ( .A1(DIN[23]), .A2(net25088), .ZN(n32) );
  NAND2_X1 U74 ( .A1(DIN[24]), .A2(net25088), .ZN(n33) );
  NAND2_X1 U75 ( .A1(DIN[25]), .A2(net25088), .ZN(n34) );
  OAI21_X1 U76 ( .B1(n150), .B2(EN), .A(n34), .ZN(n118) );
  NAND2_X1 U77 ( .A1(DIN[26]), .A2(net25088), .ZN(n99) );
  OAI21_X1 U78 ( .B1(n149), .B2(EN), .A(n99), .ZN(n117) );
  NAND2_X1 U79 ( .A1(DIN[27]), .A2(net25088), .ZN(n100) );
  NAND2_X1 U80 ( .A1(DIN[28]), .A2(net25088), .ZN(n101) );
  OAI21_X1 U81 ( .B1(n147), .B2(EN), .A(n101), .ZN(n115) );
  NAND2_X1 U82 ( .A1(DIN[29]), .A2(net25088), .ZN(n102) );
  NAND2_X1 U83 ( .A1(DIN[30]), .A2(net25088), .ZN(n103) );
endmodule


module REG_PIPO_32_00000000_00000000_4 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U9 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U10 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U11 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U12 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U13 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U14 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U15 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U16 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U17 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U18 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U19 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U21 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U22 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U23 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U25 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U26 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U27 ( .A(DIN[31]), .ZN(n9) );
  OAI22_X1 U28 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U29 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U30 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U31 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U32 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U33 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U34 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U35 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U36 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U37 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U38 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U39 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U40 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U41 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U42 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U43 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U45 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U46 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U47 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U48 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U49 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U50 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U51 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U53 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U54 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U55 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U56 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U57 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U58 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U59 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U60 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U61 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U62 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U63 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U64 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U65 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U66 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U67 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U68 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U69 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U70 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U71 ( .A(DIN[21]), .ZN(n19) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_5_00_00_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n3), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n8), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n9), .CK(CLK), .RN(RST_AN), .Q(DOUT[2]) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n10), .CK(CLK), .RN(RST_AN), .Q(DOUT[1]) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  NOR2_X1 U2 ( .A1(INIT), .A2(n12), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(n11) );
  AOI22_X1 U4 ( .A1(DIN[0]), .A2(n17), .B1(n12), .B2(DOUT[0]), .ZN(n18) );
  INV_X1 U5 ( .A(n16), .ZN(n10) );
  AOI22_X1 U6 ( .A1(DIN[1]), .A2(n17), .B1(n12), .B2(DOUT[1]), .ZN(n16) );
  INV_X1 U7 ( .A(n15), .ZN(n9) );
  AOI22_X1 U8 ( .A1(DIN[2]), .A2(n17), .B1(n12), .B2(DOUT[2]), .ZN(n15) );
  INV_X1 U9 ( .A(n14), .ZN(n8) );
  AOI22_X1 U10 ( .A1(DIN[3]), .A2(n17), .B1(n12), .B2(DOUT[3]), .ZN(n14) );
  INV_X1 U11 ( .A(n13), .ZN(n3) );
  AOI22_X1 U12 ( .A1(DIN[4]), .A2(n17), .B1(n12), .B2(DOUT[4]), .ZN(n13) );
  INV_X1 U13 ( .A(EN), .ZN(n12) );
endmodule


module REG_PIPO_1_0_0 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [0:0] DIN;
  output [0:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n1, n3, n4, n2;

  DFFR_X1 \reg_mem_reg[0]  ( .D(n4), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]), .QN(
        n3) );
  NAND3_X1 U3 ( .A1(DIN[0]), .A2(n2), .A3(EN), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n3), .B2(EN), .A(n1), .ZN(n4) );
  INV_X1 U4 ( .A(INIT), .ZN(n2) );
endmodule


module REG_PIPO_32_00000000_00000000_3 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n168), .A2(EN), .B1(n2), .B2(n103), .ZN(n136) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n103) );
  OAI22_X1 U10 ( .A1(n167), .A2(EN), .B1(n2), .B2(n102), .ZN(n135) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n102) );
  OAI22_X1 U12 ( .A1(n166), .A2(EN), .B1(n2), .B2(n101), .ZN(n134) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n101) );
  OAI22_X1 U14 ( .A1(n165), .A2(EN), .B1(n2), .B2(n100), .ZN(n133) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n100) );
  OAI22_X1 U16 ( .A1(n164), .A2(EN), .B1(n2), .B2(n99), .ZN(n132) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n99) );
  OAI22_X1 U18 ( .A1(n163), .A2(EN), .B1(n2), .B2(n34), .ZN(n131) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n34) );
  OAI22_X1 U20 ( .A1(n162), .A2(EN), .B1(n2), .B2(n33), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n33) );
  OAI22_X1 U22 ( .A1(n161), .A2(EN), .B1(n2), .B2(n32), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n160), .A2(EN), .B1(n2), .B2(n31), .ZN(n128) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n159), .A2(EN), .B1(n2), .B2(n30), .ZN(n127) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n158), .A2(EN), .B1(n2), .B2(n29), .ZN(n126) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n29) );
  OAI22_X1 U30 ( .A1(n157), .A2(EN), .B1(n3), .B2(n28), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n28) );
  OAI22_X1 U32 ( .A1(n156), .A2(EN), .B1(n3), .B2(n27), .ZN(n124) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n27) );
  OAI22_X1 U34 ( .A1(n155), .A2(EN), .B1(n3), .B2(n26), .ZN(n123) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n154), .A2(EN), .B1(n3), .B2(n25), .ZN(n122) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n25) );
  OAI22_X1 U38 ( .A1(n153), .A2(EN), .B1(n3), .B2(n24), .ZN(n121) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n24) );
  OAI22_X1 U40 ( .A1(n152), .A2(EN), .B1(n3), .B2(n23), .ZN(n120) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n151), .A2(EN), .B1(n3), .B2(n22), .ZN(n119) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n22) );
  OAI22_X1 U44 ( .A1(n150), .A2(EN), .B1(n3), .B2(n21), .ZN(n118) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n21) );
  OAI22_X1 U46 ( .A1(n149), .A2(EN), .B1(n3), .B2(n20), .ZN(n117) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n20) );
  OAI22_X1 U48 ( .A1(n148), .A2(EN), .B1(n3), .B2(n19), .ZN(n116) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n19) );
  OAI22_X1 U50 ( .A1(n147), .A2(EN), .B1(n3), .B2(n18), .ZN(n115) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n18) );
  OAI22_X1 U52 ( .A1(n146), .A2(EN), .B1(n4), .B2(n17), .ZN(n114) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n17) );
  OAI22_X1 U54 ( .A1(n145), .A2(EN), .B1(n4), .B2(n16), .ZN(n113) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n16) );
  OAI22_X1 U56 ( .A1(n144), .A2(EN), .B1(n4), .B2(n15), .ZN(n112) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n15) );
  OAI22_X1 U58 ( .A1(n143), .A2(EN), .B1(n4), .B2(n14), .ZN(n111) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n14) );
  OAI22_X1 U60 ( .A1(n142), .A2(EN), .B1(n4), .B2(n13), .ZN(n110) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n13) );
  OAI22_X1 U62 ( .A1(n141), .A2(EN), .B1(n4), .B2(n12), .ZN(n109) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n12) );
  OAI22_X1 U64 ( .A1(n140), .A2(EN), .B1(n4), .B2(n11), .ZN(n108) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n11) );
  OAI22_X1 U66 ( .A1(n139), .A2(EN), .B1(n4), .B2(n10), .ZN(n107) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n10) );
  OAI22_X1 U68 ( .A1(n138), .A2(EN), .B1(n4), .B2(n9), .ZN(n106) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n9) );
  OAI22_X1 U70 ( .A1(n137), .A2(EN), .B1(n4), .B2(n8), .ZN(n105) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n8) );
  NAND2_X1 U72 ( .A1(n104), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_2 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n168), .A2(EN), .B1(n2), .B2(n103), .ZN(n136) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n103) );
  OAI22_X1 U10 ( .A1(n167), .A2(EN), .B1(n2), .B2(n102), .ZN(n135) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n102) );
  OAI22_X1 U12 ( .A1(n166), .A2(EN), .B1(n2), .B2(n101), .ZN(n134) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n101) );
  OAI22_X1 U14 ( .A1(n165), .A2(EN), .B1(n2), .B2(n100), .ZN(n133) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n100) );
  OAI22_X1 U16 ( .A1(n164), .A2(EN), .B1(n2), .B2(n99), .ZN(n132) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n99) );
  OAI22_X1 U18 ( .A1(n163), .A2(EN), .B1(n2), .B2(n34), .ZN(n131) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n34) );
  OAI22_X1 U20 ( .A1(n162), .A2(EN), .B1(n2), .B2(n33), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n33) );
  OAI22_X1 U22 ( .A1(n161), .A2(EN), .B1(n2), .B2(n32), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n160), .A2(EN), .B1(n2), .B2(n31), .ZN(n128) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n159), .A2(EN), .B1(n2), .B2(n30), .ZN(n127) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n158), .A2(EN), .B1(n2), .B2(n29), .ZN(n126) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n29) );
  OAI22_X1 U30 ( .A1(n157), .A2(EN), .B1(n3), .B2(n28), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n28) );
  OAI22_X1 U32 ( .A1(n156), .A2(EN), .B1(n3), .B2(n27), .ZN(n124) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n27) );
  OAI22_X1 U34 ( .A1(n155), .A2(EN), .B1(n3), .B2(n26), .ZN(n123) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n154), .A2(EN), .B1(n3), .B2(n25), .ZN(n122) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n25) );
  OAI22_X1 U38 ( .A1(n153), .A2(EN), .B1(n3), .B2(n24), .ZN(n121) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n24) );
  OAI22_X1 U40 ( .A1(n152), .A2(EN), .B1(n3), .B2(n23), .ZN(n120) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n151), .A2(EN), .B1(n3), .B2(n22), .ZN(n119) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n22) );
  OAI22_X1 U44 ( .A1(n150), .A2(EN), .B1(n3), .B2(n21), .ZN(n118) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n21) );
  OAI22_X1 U46 ( .A1(n149), .A2(EN), .B1(n3), .B2(n20), .ZN(n117) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n20) );
  OAI22_X1 U48 ( .A1(n148), .A2(EN), .B1(n3), .B2(n19), .ZN(n116) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n19) );
  OAI22_X1 U50 ( .A1(n147), .A2(EN), .B1(n3), .B2(n18), .ZN(n115) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n18) );
  OAI22_X1 U52 ( .A1(n146), .A2(EN), .B1(n4), .B2(n17), .ZN(n114) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n17) );
  OAI22_X1 U54 ( .A1(n145), .A2(EN), .B1(n4), .B2(n16), .ZN(n113) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n16) );
  OAI22_X1 U56 ( .A1(n144), .A2(EN), .B1(n4), .B2(n15), .ZN(n112) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n15) );
  OAI22_X1 U58 ( .A1(n143), .A2(EN), .B1(n4), .B2(n14), .ZN(n111) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n14) );
  OAI22_X1 U60 ( .A1(n142), .A2(EN), .B1(n4), .B2(n13), .ZN(n110) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n13) );
  OAI22_X1 U62 ( .A1(n141), .A2(EN), .B1(n4), .B2(n12), .ZN(n109) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n12) );
  OAI22_X1 U64 ( .A1(n140), .A2(EN), .B1(n4), .B2(n11), .ZN(n108) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n11) );
  OAI22_X1 U66 ( .A1(n139), .A2(EN), .B1(n4), .B2(n10), .ZN(n107) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n10) );
  OAI22_X1 U68 ( .A1(n138), .A2(EN), .B1(n4), .B2(n9), .ZN(n106) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n9) );
  OAI22_X1 U70 ( .A1(n137), .A2(EN), .B1(n4), .B2(n8), .ZN(n105) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n8) );
  NAND2_X1 U72 ( .A1(n104), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n104) );
endmodule


module REG_PIPO_32_00000000_00000000_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [31:0] DIN;
  output [31:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169;

  DFFR_X1 \reg_mem_reg[31]  ( .D(n105), .CK(CLK), .RN(n7), .Q(DOUT[31]), .QN(
        n137) );
  DFFR_X1 \reg_mem_reg[30]  ( .D(n106), .CK(CLK), .RN(n7), .Q(DOUT[30]), .QN(
        n138) );
  DFFR_X1 \reg_mem_reg[29]  ( .D(n107), .CK(CLK), .RN(n7), .Q(DOUT[29]), .QN(
        n139) );
  DFFR_X1 \reg_mem_reg[28]  ( .D(n108), .CK(CLK), .RN(n7), .Q(DOUT[28]), .QN(
        n140) );
  DFFR_X1 \reg_mem_reg[27]  ( .D(n109), .CK(CLK), .RN(n7), .Q(DOUT[27]), .QN(
        n141) );
  DFFR_X1 \reg_mem_reg[26]  ( .D(n110), .CK(CLK), .RN(n7), .Q(DOUT[26]), .QN(
        n142) );
  DFFR_X1 \reg_mem_reg[25]  ( .D(n111), .CK(CLK), .RN(n7), .Q(DOUT[25]), .QN(
        n143) );
  DFFR_X1 \reg_mem_reg[24]  ( .D(n112), .CK(CLK), .RN(n7), .Q(DOUT[24]), .QN(
        n144) );
  DFFR_X1 \reg_mem_reg[23]  ( .D(n113), .CK(CLK), .RN(n7), .Q(DOUT[23]), .QN(
        n145) );
  DFFR_X1 \reg_mem_reg[22]  ( .D(n114), .CK(CLK), .RN(n7), .Q(DOUT[22]), .QN(
        n146) );
  DFFR_X1 \reg_mem_reg[21]  ( .D(n115), .CK(CLK), .RN(n6), .Q(DOUT[21]), .QN(
        n147) );
  DFFR_X1 \reg_mem_reg[20]  ( .D(n116), .CK(CLK), .RN(n6), .Q(DOUT[20]), .QN(
        n148) );
  DFFR_X1 \reg_mem_reg[19]  ( .D(n117), .CK(CLK), .RN(n6), .Q(DOUT[19]), .QN(
        n149) );
  DFFR_X1 \reg_mem_reg[18]  ( .D(n118), .CK(CLK), .RN(n6), .Q(DOUT[18]), .QN(
        n150) );
  DFFR_X1 \reg_mem_reg[17]  ( .D(n119), .CK(CLK), .RN(n6), .Q(DOUT[17]), .QN(
        n151) );
  DFFR_X1 \reg_mem_reg[16]  ( .D(n120), .CK(CLK), .RN(n6), .Q(DOUT[16]), .QN(
        n152) );
  DFFR_X1 \reg_mem_reg[15]  ( .D(n121), .CK(CLK), .RN(n6), .Q(DOUT[15]), .QN(
        n153) );
  DFFR_X1 \reg_mem_reg[14]  ( .D(n122), .CK(CLK), .RN(n6), .Q(DOUT[14]), .QN(
        n154) );
  DFFR_X1 \reg_mem_reg[13]  ( .D(n123), .CK(CLK), .RN(n6), .Q(DOUT[13]), .QN(
        n155) );
  DFFR_X1 \reg_mem_reg[12]  ( .D(n124), .CK(CLK), .RN(n6), .Q(DOUT[12]), .QN(
        n156) );
  DFFR_X1 \reg_mem_reg[11]  ( .D(n125), .CK(CLK), .RN(n6), .Q(DOUT[11]), .QN(
        n157) );
  DFFR_X1 \reg_mem_reg[10]  ( .D(n126), .CK(CLK), .RN(n5), .Q(DOUT[10]), .QN(
        n158) );
  DFFR_X1 \reg_mem_reg[9]  ( .D(n127), .CK(CLK), .RN(n5), .Q(DOUT[9]), .QN(
        n159) );
  DFFR_X1 \reg_mem_reg[8]  ( .D(n128), .CK(CLK), .RN(n5), .Q(DOUT[8]), .QN(
        n160) );
  DFFR_X1 \reg_mem_reg[7]  ( .D(n129), .CK(CLK), .RN(n5), .Q(DOUT[7]), .QN(
        n161) );
  DFFR_X1 \reg_mem_reg[6]  ( .D(n130), .CK(CLK), .RN(n5), .Q(DOUT[6]), .QN(
        n162) );
  DFFR_X1 \reg_mem_reg[5]  ( .D(n131), .CK(CLK), .RN(n5), .Q(DOUT[5]), .QN(
        n163) );
  DFFR_X1 \reg_mem_reg[4]  ( .D(n132), .CK(CLK), .RN(n5), .Q(DOUT[4]), .QN(
        n164) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n133), .CK(CLK), .RN(n5), .Q(DOUT[3]), .QN(
        n165) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n134), .CK(CLK), .RN(n5), .Q(DOUT[2]), .QN(
        n166) );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n135), .CK(CLK), .RN(n5), .Q(DOUT[1]), .QN(
        n167) );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n136), .CK(CLK), .RN(n5), .Q(DOUT[0]), .QN(
        n168) );
  BUF_X1 U2 ( .A(n169), .Z(n4) );
  BUF_X1 U3 ( .A(n169), .Z(n2) );
  BUF_X1 U4 ( .A(n169), .Z(n3) );
  BUF_X1 U5 ( .A(RST_AN), .Z(n5) );
  BUF_X1 U6 ( .A(RST_AN), .Z(n6) );
  BUF_X1 U7 ( .A(RST_AN), .Z(n7) );
  OAI22_X1 U8 ( .A1(n168), .A2(EN), .B1(n2), .B2(n104), .ZN(n136) );
  INV_X1 U9 ( .A(DIN[0]), .ZN(n104) );
  OAI22_X1 U10 ( .A1(n167), .A2(EN), .B1(n2), .B2(n103), .ZN(n135) );
  INV_X1 U11 ( .A(DIN[1]), .ZN(n103) );
  OAI22_X1 U12 ( .A1(n166), .A2(EN), .B1(n2), .B2(n102), .ZN(n134) );
  INV_X1 U13 ( .A(DIN[2]), .ZN(n102) );
  OAI22_X1 U14 ( .A1(n165), .A2(EN), .B1(n2), .B2(n101), .ZN(n133) );
  INV_X1 U15 ( .A(DIN[3]), .ZN(n101) );
  OAI22_X1 U16 ( .A1(n164), .A2(EN), .B1(n2), .B2(n100), .ZN(n132) );
  INV_X1 U17 ( .A(DIN[4]), .ZN(n100) );
  OAI22_X1 U18 ( .A1(n163), .A2(EN), .B1(n2), .B2(n99), .ZN(n131) );
  INV_X1 U19 ( .A(DIN[5]), .ZN(n99) );
  OAI22_X1 U20 ( .A1(n162), .A2(EN), .B1(n2), .B2(n34), .ZN(n130) );
  INV_X1 U21 ( .A(DIN[6]), .ZN(n34) );
  OAI22_X1 U22 ( .A1(n161), .A2(EN), .B1(n2), .B2(n33), .ZN(n129) );
  INV_X1 U23 ( .A(DIN[7]), .ZN(n33) );
  OAI22_X1 U24 ( .A1(n160), .A2(EN), .B1(n2), .B2(n32), .ZN(n128) );
  INV_X1 U25 ( .A(DIN[8]), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n159), .A2(EN), .B1(n2), .B2(n31), .ZN(n127) );
  INV_X1 U27 ( .A(DIN[9]), .ZN(n31) );
  OAI22_X1 U28 ( .A1(n158), .A2(EN), .B1(n2), .B2(n30), .ZN(n126) );
  INV_X1 U29 ( .A(DIN[10]), .ZN(n30) );
  OAI22_X1 U30 ( .A1(n157), .A2(EN), .B1(n3), .B2(n29), .ZN(n125) );
  INV_X1 U31 ( .A(DIN[11]), .ZN(n29) );
  OAI22_X1 U32 ( .A1(n156), .A2(EN), .B1(n3), .B2(n28), .ZN(n124) );
  INV_X1 U33 ( .A(DIN[12]), .ZN(n28) );
  OAI22_X1 U34 ( .A1(n155), .A2(EN), .B1(n3), .B2(n27), .ZN(n123) );
  INV_X1 U35 ( .A(DIN[13]), .ZN(n27) );
  OAI22_X1 U36 ( .A1(n154), .A2(EN), .B1(n3), .B2(n26), .ZN(n122) );
  INV_X1 U37 ( .A(DIN[14]), .ZN(n26) );
  OAI22_X1 U38 ( .A1(n153), .A2(EN), .B1(n3), .B2(n25), .ZN(n121) );
  INV_X1 U39 ( .A(DIN[15]), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n152), .A2(EN), .B1(n3), .B2(n24), .ZN(n120) );
  INV_X1 U41 ( .A(DIN[16]), .ZN(n24) );
  OAI22_X1 U42 ( .A1(n151), .A2(EN), .B1(n3), .B2(n23), .ZN(n119) );
  INV_X1 U43 ( .A(DIN[17]), .ZN(n23) );
  OAI22_X1 U44 ( .A1(n150), .A2(EN), .B1(n3), .B2(n22), .ZN(n118) );
  INV_X1 U45 ( .A(DIN[18]), .ZN(n22) );
  OAI22_X1 U46 ( .A1(n149), .A2(EN), .B1(n3), .B2(n21), .ZN(n117) );
  INV_X1 U47 ( .A(DIN[19]), .ZN(n21) );
  OAI22_X1 U48 ( .A1(n148), .A2(EN), .B1(n3), .B2(n20), .ZN(n116) );
  INV_X1 U49 ( .A(DIN[20]), .ZN(n20) );
  OAI22_X1 U50 ( .A1(n147), .A2(EN), .B1(n3), .B2(n19), .ZN(n115) );
  INV_X1 U51 ( .A(DIN[21]), .ZN(n19) );
  OAI22_X1 U52 ( .A1(n146), .A2(EN), .B1(n4), .B2(n18), .ZN(n114) );
  INV_X1 U53 ( .A(DIN[22]), .ZN(n18) );
  OAI22_X1 U54 ( .A1(n145), .A2(EN), .B1(n4), .B2(n17), .ZN(n113) );
  INV_X1 U55 ( .A(DIN[23]), .ZN(n17) );
  OAI22_X1 U56 ( .A1(n144), .A2(EN), .B1(n4), .B2(n16), .ZN(n112) );
  INV_X1 U57 ( .A(DIN[24]), .ZN(n16) );
  OAI22_X1 U58 ( .A1(n143), .A2(EN), .B1(n4), .B2(n15), .ZN(n111) );
  INV_X1 U59 ( .A(DIN[25]), .ZN(n15) );
  OAI22_X1 U60 ( .A1(n142), .A2(EN), .B1(n4), .B2(n14), .ZN(n110) );
  INV_X1 U61 ( .A(DIN[26]), .ZN(n14) );
  OAI22_X1 U62 ( .A1(n141), .A2(EN), .B1(n4), .B2(n13), .ZN(n109) );
  INV_X1 U63 ( .A(DIN[27]), .ZN(n13) );
  OAI22_X1 U64 ( .A1(n140), .A2(EN), .B1(n4), .B2(n12), .ZN(n108) );
  INV_X1 U65 ( .A(DIN[28]), .ZN(n12) );
  OAI22_X1 U66 ( .A1(n139), .A2(EN), .B1(n4), .B2(n11), .ZN(n107) );
  INV_X1 U67 ( .A(DIN[29]), .ZN(n11) );
  OAI22_X1 U68 ( .A1(n138), .A2(EN), .B1(n4), .B2(n10), .ZN(n106) );
  INV_X1 U69 ( .A(DIN[30]), .ZN(n10) );
  OAI22_X1 U70 ( .A1(n137), .A2(EN), .B1(n4), .B2(n9), .ZN(n105) );
  INV_X1 U71 ( .A(DIN[31]), .ZN(n9) );
  NAND2_X1 U72 ( .A1(n8), .A2(EN), .ZN(n169) );
  INV_X1 U73 ( .A(INIT), .ZN(n8) );
endmodule


module REG_PIPO_5_00_00_1 ( CLK, RST_AN, EN, INIT, DIN, DOUT );
  input [4:0] DIN;
  output [4:0] DOUT;
  input CLK, RST_AN, EN, INIT;
  wire   n23, n24, n3, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22;

  DFFR_X1 \reg_mem_reg[4]  ( .D(n11), .CK(CLK), .RN(RST_AN), .Q(DOUT[4]) );
  DFFR_X1 \reg_mem_reg[3]  ( .D(n12), .CK(CLK), .RN(RST_AN), .Q(DOUT[3]) );
  DFFR_X1 \reg_mem_reg[2]  ( .D(n13), .CK(CLK), .RN(RST_AN), .Q(n23), .QN(n9)
         );
  DFFR_X1 \reg_mem_reg[1]  ( .D(n14), .CK(CLK), .RN(RST_AN), .Q(n24), .QN(n3)
         );
  DFFR_X1 \reg_mem_reg[0]  ( .D(n15), .CK(CLK), .RN(RST_AN), .Q(DOUT[0]) );
  INV_X1 U2 ( .A(n3), .ZN(DOUT[1]) );
  INV_X1 U3 ( .A(n9), .ZN(DOUT[2]) );
  INV_X1 U4 ( .A(n22), .ZN(n15) );
  AOI22_X1 U5 ( .A1(DIN[0]), .A2(n21), .B1(n16), .B2(DOUT[0]), .ZN(n22) );
  INV_X1 U6 ( .A(n20), .ZN(n14) );
  AOI22_X1 U7 ( .A1(DIN[1]), .A2(n21), .B1(n16), .B2(n24), .ZN(n20) );
  INV_X1 U8 ( .A(n19), .ZN(n13) );
  AOI22_X1 U9 ( .A1(DIN[2]), .A2(n21), .B1(n16), .B2(n23), .ZN(n19) );
  INV_X1 U10 ( .A(n18), .ZN(n12) );
  AOI22_X1 U11 ( .A1(DIN[3]), .A2(n21), .B1(n16), .B2(DOUT[3]), .ZN(n18) );
  INV_X1 U12 ( .A(n17), .ZN(n11) );
  AOI22_X1 U13 ( .A1(DIN[4]), .A2(n21), .B1(n16), .B2(DOUT[4]), .ZN(n17) );
  INV_X1 U14 ( .A(EN), .ZN(n16) );
  NOR2_X1 U15 ( .A1(INIT), .A2(n16), .ZN(n21) );
endmodule


module DATAPATH_DW01_add_2 ( A, B, CI, SUM, CO );
  input [30:0] A;
  input [30:0] B;
  output [30:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U2 ( .A(A[11]), .B(n1), .Z(SUM[11]) );
  NOR2_X1 U3 ( .A1(n6), .A2(n47), .ZN(n1) );
  XOR2_X1 U4 ( .A(n28), .B(A[20]), .Z(SUM[20]) );
  XOR2_X1 U5 ( .A(n24), .B(A[24]), .Z(SUM[24]) );
  XNOR2_X1 U6 ( .A(n2), .B(A[27]), .ZN(SUM[27]) );
  NAND2_X1 U7 ( .A1(A[26]), .A2(n12), .ZN(n2) );
  XNOR2_X1 U8 ( .A(n3), .B(A[23]), .ZN(SUM[23]) );
  NAND2_X1 U9 ( .A1(A[22]), .A2(n9), .ZN(n3) );
  XOR2_X1 U10 ( .A(n7), .B(A[16]), .Z(SUM[16]) );
  XOR2_X1 U11 ( .A(A[19]), .B(n4), .Z(SUM[19]) );
  NOR2_X1 U12 ( .A1(n31), .A2(n33), .ZN(n4) );
  XNOR2_X1 U13 ( .A(n5), .B(A[30]), .ZN(SUM[30]) );
  NAND2_X1 U14 ( .A1(n10), .A2(A[29]), .ZN(n5) );
  XOR2_X1 U15 ( .A(n6), .B(n47), .Z(SUM[10]) );
  XOR2_X1 U16 ( .A(n13), .B(n51), .Z(SUM[9]) );
  NOR2_X1 U17 ( .A1(n49), .A2(n41), .ZN(n14) );
  NOR2_X1 U18 ( .A1(n46), .A2(n40), .ZN(n45) );
  OR2_X1 U19 ( .A1(n51), .A2(n13), .ZN(n6) );
  INV_X1 U20 ( .A(n25), .ZN(n27) );
  INV_X1 U21 ( .A(n29), .ZN(n32) );
  INV_X1 U22 ( .A(n20), .ZN(n23) );
  NOR2_X1 U23 ( .A1(n36), .A2(n8), .ZN(n7) );
  OR2_X1 U24 ( .A1(n34), .A2(n35), .ZN(n8) );
  XOR2_X1 U25 ( .A(A[13]), .B(n44), .Z(SUM[13]) );
  XOR2_X1 U26 ( .A(A[5]), .B(n17), .Z(SUM[5]) );
  XOR2_X1 U27 ( .A(A[8]), .B(n14), .Z(SUM[8]) );
  AND2_X1 U28 ( .A1(n17), .A2(A[5]), .ZN(n16) );
  AND2_X1 U29 ( .A1(n44), .A2(A[13]), .ZN(n43) );
  NOR2_X1 U30 ( .A1(n20), .A2(n21), .ZN(n19) );
  XNOR2_X1 U31 ( .A(n15), .B(A[7]), .ZN(SUM[7]) );
  NAND2_X1 U32 ( .A1(n16), .A2(A[6]), .ZN(n15) );
  XNOR2_X1 U33 ( .A(n42), .B(A[15]), .ZN(SUM[15]) );
  NAND2_X1 U34 ( .A1(n43), .A2(A[14]), .ZN(n42) );
  XNOR2_X1 U35 ( .A(A[3]), .B(SUM[2]), .ZN(SUM[3]) );
  XOR2_X1 U36 ( .A(A[14]), .B(n43), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(A[6]), .B(n16), .Z(SUM[6]) );
  XOR2_X1 U38 ( .A(A[12]), .B(n45), .Z(SUM[12]) );
  XOR2_X1 U39 ( .A(A[4]), .B(n38), .Z(SUM[4]) );
  NAND4_X1 U40 ( .A1(A[4]), .A2(A[5]), .A3(A[6]), .A4(A[7]), .ZN(n41) );
  NAND4_X1 U41 ( .A1(A[11]), .A2(A[10]), .A3(A[9]), .A4(A[8]), .ZN(n40) );
  NOR2_X1 U42 ( .A1(n25), .A2(n26), .ZN(n24) );
  NOR2_X1 U43 ( .A1(n29), .A2(n30), .ZN(n28) );
  NOR2_X1 U44 ( .A1(n48), .A2(n49), .ZN(n17) );
  AND2_X1 U45 ( .A1(A[12]), .A2(n45), .ZN(n44) );
  XOR2_X1 U46 ( .A(A[21]), .B(n27), .Z(SUM[21]) );
  XOR2_X1 U47 ( .A(A[17]), .B(n32), .Z(SUM[17]) );
  XOR2_X1 U48 ( .A(A[18]), .B(n11), .Z(SUM[18]) );
  XOR2_X1 U49 ( .A(n9), .B(A[22]), .Z(SUM[22]) );
  XOR2_X1 U50 ( .A(n23), .B(A[25]), .Z(SUM[25]) );
  XOR2_X1 U51 ( .A(n19), .B(A[28]), .Z(SUM[28]) );
  XNOR2_X1 U52 ( .A(n12), .B(n22), .ZN(SUM[26]) );
  XOR2_X1 U53 ( .A(n10), .B(A[29]), .Z(SUM[29]) );
  NOR2_X1 U54 ( .A1(SUM[2]), .A2(n50), .ZN(n38) );
  NAND2_X1 U55 ( .A1(n28), .A2(A[20]), .ZN(n25) );
  NAND2_X1 U56 ( .A1(n24), .A2(A[24]), .ZN(n20) );
  NAND2_X1 U57 ( .A1(n7), .A2(A[16]), .ZN(n29) );
  NAND2_X1 U58 ( .A1(n14), .A2(A[8]), .ZN(n13) );
  AND2_X1 U59 ( .A1(A[21]), .A2(n27), .ZN(n9) );
  AND2_X1 U60 ( .A1(n19), .A2(A[28]), .ZN(n10) );
  AND2_X1 U61 ( .A1(A[17]), .A2(n32), .ZN(n11) );
  NAND2_X1 U62 ( .A1(A[12]), .A2(A[13]), .ZN(n35) );
  AND2_X1 U63 ( .A1(A[25]), .A2(n23), .ZN(n12) );
  NAND2_X1 U64 ( .A1(A[14]), .A2(A[15]), .ZN(n34) );
  INV_X1 U65 ( .A(A[2]), .ZN(SUM[2]) );
  INV_X1 U66 ( .A(A[4]), .ZN(n48) );
  INV_X1 U67 ( .A(A[18]), .ZN(n33) );
  INV_X1 U68 ( .A(A[26]), .ZN(n22) );
  INV_X1 U69 ( .A(A[9]), .ZN(n51) );
  INV_X1 U70 ( .A(A[3]), .ZN(n50) );
  NAND3_X1 U71 ( .A1(A[26]), .A2(A[27]), .A3(A[25]), .ZN(n21) );
  NAND3_X1 U72 ( .A1(A[22]), .A2(A[23]), .A3(A[21]), .ZN(n26) );
  NAND3_X1 U73 ( .A1(A[18]), .A2(A[19]), .A3(A[17]), .ZN(n30) );
  INV_X1 U74 ( .A(n11), .ZN(n31) );
  NAND3_X1 U75 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n36) );
  INV_X1 U76 ( .A(n40), .ZN(n39) );
  INV_X1 U77 ( .A(n41), .ZN(n37) );
  INV_X1 U78 ( .A(n14), .ZN(n46) );
  INV_X1 U79 ( .A(A[10]), .ZN(n47) );
  INV_X1 U80 ( .A(n38), .ZN(n49) );
endmodule


module DATAPATH ( CLK, RST_AN, .CTRL_WORD({\CTRL_WORD[J_TYPE_IMM_SEL] , 
        \CTRL_WORD[R_TYPE_SEL] , \CTRL_WORD[IMM_SEL] , 
        \CTRL_WORD[PC_PLS_4_SEL] , \CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] , \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] , 
        \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] , 
        \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] , 
        \CTRL_WORD[RF_WEN] }), INSTR_CU, .HZRD_SIG({\HZRD_SIG[STALL_FD] , 
        \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , 
        \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] }), .DP_SIG({
        \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] , 
        \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] , 
        \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] , 
        \DP_SIG[INSTR_OPCODE_M][0] }), IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] INSTR_CU;
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN, \CTRL_WORD[J_TYPE_IMM_SEL] , \CTRL_WORD[R_TYPE_SEL] ,
         \CTRL_WORD[IMM_SEL] , \CTRL_WORD[PC_PLS_4_SEL] ,
         \CTRL_WORD[ALU_FUNC][3] , \CTRL_WORD[ALU_FUNC][2] ,
         \CTRL_WORD[ALU_FUNC][1] , \CTRL_WORD[ALU_FUNC][0] ,
         \CTRL_WORD[JUMP_EN] , \CTRL_WORD[BRANCH_EN] ,
         \CTRL_WORD[COMP_0_INVERT] , \CTRL_WORD[DMEM_WEN] ,
         \CTRL_WORD[RF_WB_DMEM_DOUT_SEL] , \CTRL_WORD[JAL_EN] ,
         \CTRL_WORD[RF_WEN] , \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] ,
         \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] ,
         \HZRD_SIG[FLUSH_MWB] ;
  output \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  wire   \npc_f[31] , n144, n145, n146, n147, n148, n149, n150, n151, n153,
         n154, n155, n156, n157, n158, n160, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n184, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n277, n278, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n302, net17712, net17717, net17718, net26009,
         net26007, net26021, net26019, net26025, net26023, net26033, net26031,
         net26029, net34307, net34306, net34464, net34633, net34948, net34947,
         net34991, net34990, net36835, net36877, net38403, net38918, net44768,
         n162, n1, n2, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n152,
         n159, n161, n183, n185, n186;
  wire   [30:0] pc_pls_4_f;
  wire   [31:0] pc_pls_4_d;
  wire   [31:0] instr_d;
  wire   [4:0] rf_waddr_d;
  wire   [31:0] rf_dout1_d;
  wire   [31:0] rf_dout2_d;
  wire   [4:0] rf_waddr_wb;
  wire   [31:16] imm_d;
  wire   [5:0] instr_opcode_e;
  wire   [31:0] pc_pls_4_e;
  wire   [31:0] rf_dout1_e;
  wire   [31:0] rf_dout2_e;
  wire   [31:0] imm_e;
  wire   [4:0] rs2_e;
  wire   [4:0] rs3_e;
  wire   [31:0] alu_a_e;
  wire   [31:0] alu_out_e;
  wire   [31:0] pc_pls_4_m;
  wire   [4:0] rf_waddr_m;
  wire   [31:0] pc_pls_4_wb;
  wire   [31:0] alu_out_wb;
  wire   [31:0] dmem_dout_wb;
  assign INSTR_CU[31] = IMEM_DOUT[31];
  assign INSTR_CU[30] = IMEM_DOUT[30];
  assign INSTR_CU[29] = IMEM_DOUT[29];
  assign INSTR_CU[28] = IMEM_DOUT[28];
  assign INSTR_CU[27] = IMEM_DOUT[27];
  assign INSTR_CU[26] = IMEM_DOUT[26];
  assign INSTR_CU[25] = IMEM_DOUT[25];
  assign INSTR_CU[24] = IMEM_DOUT[24];
  assign INSTR_CU[23] = IMEM_DOUT[23];
  assign INSTR_CU[22] = IMEM_DOUT[22];
  assign INSTR_CU[21] = IMEM_DOUT[21];
  assign INSTR_CU[20] = IMEM_DOUT[20];
  assign INSTR_CU[19] = IMEM_DOUT[19];
  assign INSTR_CU[18] = IMEM_DOUT[18];
  assign INSTR_CU[17] = IMEM_DOUT[17];
  assign INSTR_CU[16] = IMEM_DOUT[16];
  assign INSTR_CU[15] = IMEM_DOUT[15];
  assign INSTR_CU[14] = IMEM_DOUT[14];
  assign INSTR_CU[13] = IMEM_DOUT[13];
  assign INSTR_CU[12] = IMEM_DOUT[12];
  assign INSTR_CU[11] = IMEM_DOUT[11];
  assign INSTR_CU[10] = IMEM_DOUT[10];
  assign INSTR_CU[9] = IMEM_DOUT[9];
  assign INSTR_CU[8] = IMEM_DOUT[8];
  assign INSTR_CU[7] = IMEM_DOUT[7];
  assign INSTR_CU[6] = IMEM_DOUT[6];
  assign INSTR_CU[5] = IMEM_DOUT[5];
  assign INSTR_CU[4] = IMEM_DOUT[4];
  assign INSTR_CU[3] = IMEM_DOUT[3];
  assign INSTR_CU[2] = IMEM_DOUT[2];
  assign INSTR_CU[1] = IMEM_DOUT[1];
  assign INSTR_CU[0] = IMEM_DOUT[0];

  REG_PIPO_32_fffffffc_fffffffc U_PC_REG ( .CLK(CLK), .RST_AN(n40), .EN(1'b1), 
        .INIT(1'b0), .DIN({\npc_f[31] , n43, n44, n45, n46, n47, n48, n49, n50, 
        n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
        n65, n66, n67, n68, n69, n70, n71, n72, n119}), .DOUT(IMEM_ADDR) );
  REG_PIPO_32_00000000_00000000_0 U_PC_PLS_4_REG_FD ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN({1'b0, pc_pls_4_f}), 
        .DOUT(pc_pls_4_d) );
  REG_PIPO_32_00000000_00000000_11 U_INSTR_REG_FD ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_FD] ), .DIN(IMEM_DOUT), .DOUT(instr_d) );
  RF_ADDR_W5_DATA_W32 U_RF ( .CLK(CLK), .RST_AN(n39), .ENABLE(1'b1), .RD1(1'b1), .RD2(1'b1), .WR(\CTRL_WORD[RF_WEN] ), .ADD_WR(rf_waddr_d), .ADD_RD1(
        instr_d[25:21]), .ADD_RD2(instr_d[20:16]), .DATAIN({n120, n17, n1, 
        net17712, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
        n131, n132, n133, n134, n135, n136, n137, n138, n139, n8, n140, n141, 
        n142, n143, n152, n159, n161, n183}), .OUT1(rf_dout1_d), .OUT2(
        rf_dout2_d) );
  REG_PIPO_6_00_00_0 U_INSTR_OPCODE_REG_DE ( .CLK(CLK), .RST_AN(n39), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[31:26]), .DOUT(instr_opcode_e) );
  REG_PIPO_32_00000000_00000000_10 U_PC_PLS_4_REG_DE ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(pc_pls_4_d), .DOUT(
        pc_pls_4_e) );
  REG_PIPO_32_00000000_00000000_9 U_RF_DOUT1_REG_DE ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout1_d), .DOUT(
        rf_dout1_e) );
  REG_PIPO_32_00000000_00000000_8 U_RF_DOUT2_REG_DE ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN(rf_dout2_d), .DOUT(
        rf_dout2_e) );
  REG_PIPO_32_00000000_00000000_7 U_IMM_REG_DE ( .CLK(CLK), .RST_AN(n40), .EN(
        1'b1), .INIT(\HZRD_SIG[FLUSH_DE] ), .DIN({imm_d[31], imm_d[31], 
        imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[31], imm_d[24:16], 
        instr_d[15:0]}), .DOUT(imm_e) );
  REG_PIPO_5_00_00_0 U_RS2_REG_DE ( .CLK(CLK), .RST_AN(n39), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[20:16]), .DOUT(rs2_e) );
  REG_PIPO_5_00_00_3 U_RS3_REG_DE ( .CLK(CLK), .RST_AN(n39), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_DE] ), .DIN(instr_d[15:11]), .DOUT(rs3_e) );
  ALU_DATA_W32 U_ALU ( .FUNC({\CTRL_WORD[ALU_FUNC][3] , 
        \CTRL_WORD[ALU_FUNC][2] , \CTRL_WORD[ALU_FUNC][1] , 
        \CTRL_WORD[ALU_FUNC][0] }), .A(alu_a_e), .B({n89, n90, n91, n92, n93, 
        n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
        n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
        net17718, net17717}), .RES(alu_out_e) );
  REG_PIPO_6_00_00_1 U_INSTR_OPCODE_REG_EM ( .CLK(CLK), .RST_AN(n39), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(instr_opcode_e), .DOUT({
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }) );
  REG_PIPO_32_00000000_00000000_6 U_PC_PLS_4_REG_EM ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(pc_pls_4_e), .DOUT(
        pc_pls_4_m) );
  REG_PIPO_32_00000000_00000000_5 U_ALU_OUT_REG_EM ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(alu_out_e), .DOUT(
        DMEM_RWADDR) );
  REG_PIPO_32_00000000_00000000_4 U_DMEM_DOUT_REG_EM ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN(rf_dout2_e), .DOUT(
        DMEM_DIN) );
  REG_PIPO_5_00_00_2 U_RF_WADDR_REG_EM ( .CLK(CLK), .RST_AN(n39), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_EM] ), .DIN({n73, n74, n75, n76, n77}), .DOUT(
        rf_waddr_m) );
  REG_PIPO_1_0_0 U_IS_0_REG_EM ( .CLK(CLK), .RST_AN(n40), .EN(1'b1), .INIT(
        \HZRD_SIG[FLUSH_EM] ), .DIN(n302), .DOUT(\DP_SIG[CMPR_0_IS_0_M] ) );
  REG_PIPO_32_00000000_00000000_3 U_PC_PLS_4_REG_MWB ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(pc_pls_4_m), .DOUT(
        pc_pls_4_wb) );
  REG_PIPO_32_00000000_00000000_2 U_ALU_OUT_REG_MWB ( .CLK(CLK), .RST_AN(n40), 
        .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_RWADDR), .DOUT(
        alu_out_wb) );
  REG_PIPO_32_00000000_00000000_1 U_DMEM_DOUT_REG_MWB ( .CLK(CLK), .RST_AN(n40), .EN(1'b1), .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(DMEM_DOUT), .DOUT(dmem_dout_wb) );
  REG_PIPO_5_00_00_1 U_RF_WADDR_REG_MWB ( .CLK(CLK), .RST_AN(n39), .EN(1'b1), 
        .INIT(\HZRD_SIG[FLUSH_MWB] ), .DIN(rf_waddr_m), .DOUT(rf_waddr_wb) );
  DATAPATH_DW01_add_2 add_242 ( .A(IMEM_ADDR[30:0]), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(pc_pls_4_f) );
  BUF_X1 U5 ( .A(n151), .Z(net34948) );
  OR3_X2 U7 ( .A1(n14), .A2(n13), .A3(n15), .ZN(n1) );
  BUF_X2 U8 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n24) );
  CLKBUF_X2 U9 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n22) );
  BUF_X2 U10 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net34464) );
  MUX2_X1 U11 ( .A(rf_dout2_e[25]), .B(imm_e[25]), .S(net34633), .Z(n95) );
  BUF_X1 U12 ( .A(n37), .Z(n31) );
  OAI21_X2 U13 ( .B1(n25), .B2(n86), .A(n286), .ZN(alu_a_e[23]) );
  CLKBUF_X3 U14 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(net26019) );
  BUF_X1 U15 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(net26021) );
  BUF_X1 U16 ( .A(n23), .Z(n38) );
  BUF_X1 U17 ( .A(n151), .Z(net26029) );
  OR3_X2 U18 ( .A1(n19), .A2(n18), .A3(n20), .ZN(n17) );
  CLKBUF_X3 U19 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net34306) );
  OAI21_X2 U20 ( .B1(n25), .B2(n82), .A(n282), .ZN(alu_a_e[27]) );
  AOI222_X1 U21 ( .A1(dmem_dout_wb[28]), .A2(net26021), .B1(net38918), .B2(
        alu_out_wb[28]), .C1(net26031), .C2(pc_pls_4_wb[28]), .ZN(n162) );
  INV_X1 U22 ( .A(n162), .ZN(net17712) );
  NOR2_X2 U23 ( .A1(n7), .A2(n6), .ZN(net38918) );
  BUF_X2 U24 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(n6) );
  NOR2_X1 U25 ( .A1(n6), .A2(n2), .ZN(n151) );
  NOR2_X1 U26 ( .A1(n6), .A2(n2), .ZN(net36835) );
  NOR2_X1 U27 ( .A1(n7), .A2(n6), .ZN(n150) );
  INV_X1 U28 ( .A(n2), .ZN(n7) );
  INV_X1 U29 ( .A(\CTRL_WORD[JAL_EN] ), .ZN(n2) );
  BUF_X1 U30 ( .A(n150), .Z(net44768) );
  CLKBUF_X1 U31 ( .A(\CTRL_WORD[RF_WB_DMEM_DOUT_SEL] ), .Z(net38403) );
  BUF_X1 U32 ( .A(net26007), .Z(net36877) );
  OR3_X2 U33 ( .A1(n10), .A2(n9), .A3(n11), .ZN(n8) );
  BUF_X2 U34 ( .A(n37), .Z(n30) );
  AND2_X1 U35 ( .A1(dmem_dout_wb[8]), .A2(net26021), .ZN(n9) );
  AND2_X1 U36 ( .A1(net44768), .A2(alu_out_wb[8]), .ZN(n10) );
  AND2_X1 U37 ( .A1(pc_pls_4_wb[8]), .A2(net26031), .ZN(n11) );
  MUX2_X1 U38 ( .A(rf_dout2_e[1]), .B(imm_e[1]), .S(n12), .Z(net17718) );
  BUF_X1 U39 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(n12) );
  MUX2_X1 U40 ( .A(rf_dout2_e[0]), .B(imm_e[0]), .S(n12), .Z(net17717) );
  AND2_X1 U41 ( .A1(dmem_dout_wb[29]), .A2(net38403), .ZN(n13) );
  AND2_X1 U42 ( .A1(net34991), .A2(alu_out_wb[29]), .ZN(n14) );
  AND2_X1 U43 ( .A1(pc_pls_4_wb[29]), .A2(net36835), .ZN(n15) );
  OR2_X1 U44 ( .A1(n33), .A2(n87), .ZN(n16) );
  NAND2_X2 U45 ( .A1(n16), .A2(n287), .ZN(alu_a_e[22]) );
  BUF_X1 U46 ( .A(n151), .Z(net34947) );
  BUF_X1 U47 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n21) );
  MUX2_X1 U48 ( .A(pc_pls_4_e[19]), .B(rf_dout1_e[19]), .S(n32), .Z(
        alu_a_e[19]) );
  BUF_X2 U49 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net26009) );
  OAI21_X2 U50 ( .B1(n33), .B2(n83), .A(n283), .ZN(alu_a_e[26]) );
  AND2_X1 U51 ( .A1(dmem_dout_wb[30]), .A2(net26019), .ZN(n18) );
  AND2_X1 U52 ( .A1(net34990), .A2(alu_out_wb[30]), .ZN(n19) );
  AND2_X1 U53 ( .A1(pc_pls_4_wb[30]), .A2(net36835), .ZN(n20) );
  BUF_X1 U54 ( .A(n150), .Z(net34991) );
  BUF_X1 U55 ( .A(n150), .Z(net26023) );
  BUF_X1 U56 ( .A(n151), .Z(net26033) );
  CLKBUF_X2 U57 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net26007) );
  CLKBUF_X1 U58 ( .A(n37), .Z(n29) );
  OR2_X2 U59 ( .A1(rf_waddr_wb[0]), .A2(\CTRL_WORD[JAL_EN] ), .ZN(
        rf_waddr_d[0]) );
  OAI21_X1 U60 ( .B1(n30), .B2(n79), .A(n278), .ZN(alu_a_e[30]) );
  OAI21_X2 U61 ( .B1(n25), .B2(n81), .A(n281), .ZN(alu_a_e[28]) );
  BUF_X2 U62 ( .A(n23), .Z(n37) );
  BUF_X1 U63 ( .A(n150), .Z(net34990) );
  BUF_X1 U64 ( .A(\CTRL_WORD[PC_PLS_4_SEL] ), .Z(n23) );
  MUX2_X1 U65 ( .A(rf_dout1_e[18]), .B(pc_pls_4_e[18]), .S(n38), .Z(
        alu_a_e[18]) );
  MUX2_X1 U66 ( .A(rf_dout1_e[16]), .B(pc_pls_4_e[16]), .S(n37), .Z(
        alu_a_e[16]) );
  INV_X1 U67 ( .A(n32), .ZN(n25) );
  INV_X1 U68 ( .A(n32), .ZN(n33) );
  OAI21_X2 U69 ( .B1(n25), .B2(n85), .A(n285), .ZN(alu_a_e[24]) );
  CLKBUF_X1 U70 ( .A(net26007), .Z(net34633) );
  INV_X1 U71 ( .A(n149), .ZN(n139) );
  MUX2_X1 U72 ( .A(rf_dout2_e[10]), .B(imm_e[10]), .S(net34306), .Z(n110) );
  OAI21_X1 U73 ( .B1(n33), .B2(n80), .A(n280), .ZN(alu_a_e[29]) );
  CLKBUF_X1 U74 ( .A(\CTRL_WORD[IMM_SEL] ), .Z(net34307) );
  MUX2_X1 U75 ( .A(rf_dout2_e[11]), .B(imm_e[11]), .S(net34306), .Z(n109) );
  OAI21_X1 U76 ( .B1(n33), .B2(n88), .A(n288), .ZN(alu_a_e[21]) );
  MUX2_X1 U77 ( .A(rf_dout2_e[2]), .B(imm_e[2]), .S(net34464), .Z(n118) );
  OAI21_X1 U78 ( .B1(n33), .B2(n78), .A(n277), .ZN(alu_a_e[31]) );
  MUX2_X1 U79 ( .A(rf_dout2_e[4]), .B(imm_e[4]), .S(net26007), .Z(n116) );
  OAI21_X1 U80 ( .B1(n33), .B2(n84), .A(n284), .ZN(alu_a_e[25]) );
  NAND2_X1 U81 ( .A1(rf_dout1_e[20]), .A2(n26), .ZN(n27) );
  NAND2_X1 U82 ( .A1(pc_pls_4_e[20]), .A2(n25), .ZN(n28) );
  NAND2_X2 U83 ( .A1(n27), .A2(n28), .ZN(alu_a_e[20]) );
  INV_X1 U84 ( .A(n29), .ZN(n26) );
  OR2_X2 U85 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[2]), .ZN(
        rf_waddr_d[2]) );
  BUF_X1 U86 ( .A(n42), .Z(n34) );
  BUF_X1 U87 ( .A(n42), .Z(n35) );
  BUF_X1 U88 ( .A(n42), .Z(n36) );
  BUF_X1 U89 ( .A(n150), .Z(net26025) );
  BUF_X1 U90 ( .A(n151), .Z(net26031) );
  INV_X1 U91 ( .A(rf_dout1_e[31]), .ZN(n78) );
  NAND2_X1 U92 ( .A1(pc_pls_4_e[31]), .A2(n30), .ZN(n277) );
  INV_X1 U93 ( .A(rf_dout1_e[26]), .ZN(n83) );
  NAND2_X1 U94 ( .A1(pc_pls_4_e[26]), .A2(n31), .ZN(n283) );
  INV_X1 U95 ( .A(rf_dout1_e[25]), .ZN(n84) );
  NAND2_X1 U96 ( .A1(pc_pls_4_e[25]), .A2(n31), .ZN(n284) );
  INV_X1 U97 ( .A(rf_dout1_e[27]), .ZN(n82) );
  NAND2_X1 U98 ( .A1(pc_pls_4_e[27]), .A2(n31), .ZN(n282) );
  INV_X1 U99 ( .A(rf_dout1_e[24]), .ZN(n85) );
  NAND2_X1 U100 ( .A1(pc_pls_4_e[24]), .A2(n30), .ZN(n285) );
  INV_X1 U101 ( .A(rf_dout1_e[23]), .ZN(n86) );
  NAND2_X1 U102 ( .A1(pc_pls_4_e[23]), .A2(n30), .ZN(n286) );
  INV_X1 U103 ( .A(rf_dout1_e[21]), .ZN(n88) );
  NAND2_X1 U104 ( .A1(pc_pls_4_e[21]), .A2(n29), .ZN(n288) );
  INV_X1 U105 ( .A(rf_dout1_e[22]), .ZN(n87) );
  NAND2_X1 U106 ( .A1(pc_pls_4_e[22]), .A2(n29), .ZN(n287) );
  INV_X1 U107 ( .A(rf_dout1_e[29]), .ZN(n80) );
  NAND2_X1 U108 ( .A1(pc_pls_4_e[29]), .A2(n31), .ZN(n280) );
  INV_X1 U109 ( .A(rf_dout1_e[28]), .ZN(n81) );
  NAND2_X1 U110 ( .A1(pc_pls_4_e[28]), .A2(n31), .ZN(n281) );
  AOI222_X1 U111 ( .A1(dmem_dout_wb[9]), .A2(net26021), .B1(net38918), .B2(
        alu_out_wb[9]), .C1(pc_pls_4_wb[9]), .C2(net36835), .ZN(n149) );
  NOR4_X1 U112 ( .A1(rf_dout1_e[23]), .A2(rf_dout1_e[22]), .A3(rf_dout1_e[21]), 
        .A4(rf_dout1_e[20]), .ZN(n222) );
  NOR4_X1 U113 ( .A1(rf_dout1_e[5]), .A2(rf_dout1_e[4]), .A3(rf_dout1_e[3]), 
        .A4(rf_dout1_e[31]), .ZN(n225) );
  AOI222_X1 U114 ( .A1(dmem_dout_wb[6]), .A2(net26019), .B1(net38918), .B2(
        alu_out_wb[6]), .C1(pc_pls_4_wb[6]), .C2(net36835), .ZN(n154) );
  AOI222_X1 U115 ( .A1(dmem_dout_wb[7]), .A2(net26021), .B1(net26023), .B2(
        alu_out_wb[7]), .C1(pc_pls_4_wb[7]), .C2(net26033), .ZN(n153) );
  AOI222_X1 U116 ( .A1(dmem_dout_wb[3]), .A2(net26019), .B1(net34990), .B2(
        alu_out_wb[3]), .C1(pc_pls_4_wb[3]), .C2(net34947), .ZN(n157) );
  AOI222_X1 U117 ( .A1(dmem_dout_wb[4]), .A2(net38403), .B1(net34991), .B2(
        alu_out_wb[4]), .C1(pc_pls_4_wb[4]), .C2(net34947), .ZN(n156) );
  AOI222_X1 U118 ( .A1(dmem_dout_wb[5]), .A2(net26021), .B1(net26023), .B2(
        alu_out_wb[5]), .C1(pc_pls_4_wb[5]), .C2(net34948), .ZN(n155) );
  AOI222_X1 U119 ( .A1(dmem_dout_wb[31]), .A2(net26019), .B1(net34990), .B2(
        alu_out_wb[31]), .C1(pc_pls_4_wb[31]), .C2(net34948), .ZN(n158) );
  NAND2_X1 U120 ( .A1(n227), .A2(n228), .ZN(imm_d[31]) );
  NAND2_X1 U121 ( .A1(instr_d[25]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n228) );
  INV_X1 U122 ( .A(\CTRL_WORD[R_TYPE_SEL] ), .ZN(n186) );
  NAND2_X1 U123 ( .A1(n227), .A2(n231), .ZN(imm_d[22]) );
  NAND2_X1 U124 ( .A1(instr_d[22]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n231) );
  NAND2_X1 U125 ( .A1(n227), .A2(n230), .ZN(imm_d[23]) );
  NAND2_X1 U126 ( .A1(instr_d[23]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n230) );
  NAND2_X1 U127 ( .A1(n227), .A2(n229), .ZN(imm_d[24]) );
  NAND2_X1 U128 ( .A1(instr_d[24]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n229) );
  NAND2_X1 U129 ( .A1(n227), .A2(n237), .ZN(imm_d[16]) );
  NAND2_X1 U130 ( .A1(instr_d[16]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n237) );
  NAND2_X1 U131 ( .A1(n227), .A2(n236), .ZN(imm_d[17]) );
  NAND2_X1 U132 ( .A1(instr_d[17]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n236) );
  NAND2_X1 U133 ( .A1(n227), .A2(n235), .ZN(imm_d[18]) );
  NAND2_X1 U134 ( .A1(instr_d[18]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n235) );
  NAND2_X1 U135 ( .A1(n227), .A2(n234), .ZN(imm_d[19]) );
  NAND2_X1 U136 ( .A1(instr_d[19]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n234) );
  NAND2_X1 U137 ( .A1(n227), .A2(n233), .ZN(imm_d[20]) );
  NAND2_X1 U138 ( .A1(instr_d[20]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n233) );
  NAND2_X1 U139 ( .A1(n227), .A2(n232), .ZN(imm_d[21]) );
  NAND2_X1 U140 ( .A1(instr_d[21]), .A2(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n232) );
  OR2_X1 U141 ( .A1(\CTRL_WORD[JAL_EN] ), .A2(rf_waddr_wb[1]), .ZN(
        rf_waddr_d[1]) );
  NAND4_X1 U142 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(n218) );
  NOR4_X1 U143 ( .A1(rf_dout1_e[12]), .A2(rf_dout1_e[11]), .A3(rf_dout1_e[10]), 
        .A4(rf_dout1_e[0]), .ZN(n219) );
  NOR4_X1 U144 ( .A1(rf_dout1_e[16]), .A2(rf_dout1_e[15]), .A3(rf_dout1_e[14]), 
        .A4(rf_dout1_e[13]), .ZN(n220) );
  NOR4_X1 U145 ( .A1(rf_dout1_e[1]), .A2(rf_dout1_e[19]), .A3(rf_dout1_e[18]), 
        .A4(rf_dout1_e[17]), .ZN(n221) );
  NAND4_X1 U146 ( .A1(n223), .A2(n224), .A3(n225), .A4(n226), .ZN(n217) );
  NOR4_X1 U147 ( .A1(rf_dout1_e[27]), .A2(rf_dout1_e[26]), .A3(rf_dout1_e[25]), 
        .A4(rf_dout1_e[24]), .ZN(n223) );
  NOR4_X1 U148 ( .A1(rf_dout1_e[30]), .A2(rf_dout1_e[2]), .A3(rf_dout1_e[29]), 
        .A4(rf_dout1_e[28]), .ZN(n224) );
  NOR4_X1 U149 ( .A1(rf_dout1_e[9]), .A2(rf_dout1_e[8]), .A3(rf_dout1_e[7]), 
        .A4(rf_dout1_e[6]), .ZN(n226) );
  NAND2_X1 U150 ( .A1(instr_d[15]), .A2(n185), .ZN(n227) );
  INV_X1 U151 ( .A(\CTRL_WORD[J_TYPE_IMM_SEL] ), .ZN(n185) );
  AOI222_X1 U152 ( .A1(dmem_dout_wb[0]), .A2(net26021), .B1(net38918), .B2(
        alu_out_wb[0]), .C1(pc_pls_4_wb[0]), .C2(net26029), .ZN(n182) );
  AOI222_X1 U153 ( .A1(dmem_dout_wb[1]), .A2(net26021), .B1(net38918), .B2(
        alu_out_wb[1]), .C1(pc_pls_4_wb[1]), .C2(net36835), .ZN(n171) );
  AOI222_X1 U154 ( .A1(dmem_dout_wb[2]), .A2(net26021), .B1(net26023), .B2(
        alu_out_wb[2]), .C1(pc_pls_4_wb[2]), .C2(net26031), .ZN(n160) );
  AOI222_X1 U155 ( .A1(dmem_dout_wb[12]), .A2(net26019), .B1(net26023), .B2(
        alu_out_wb[12]), .C1(pc_pls_4_wb[12]), .C2(net26033), .ZN(n179) );
  AOI222_X1 U156 ( .A1(dmem_dout_wb[13]), .A2(net26019), .B1(net38918), .B2(
        alu_out_wb[13]), .C1(pc_pls_4_wb[13]), .C2(net36835), .ZN(n178) );
  AOI222_X1 U157 ( .A1(dmem_dout_wb[14]), .A2(net26019), .B1(net38918), .B2(
        alu_out_wb[14]), .C1(net34948), .C2(pc_pls_4_wb[14]), .ZN(n177) );
  AOI222_X1 U158 ( .A1(dmem_dout_wb[15]), .A2(net38403), .B1(net26025), .B2(
        alu_out_wb[15]), .C1(pc_pls_4_wb[15]), .C2(net34947), .ZN(n176) );
  AOI222_X1 U159 ( .A1(dmem_dout_wb[16]), .A2(net38403), .B1(net44768), .B2(
        alu_out_wb[16]), .C1(pc_pls_4_wb[16]), .C2(net36835), .ZN(n175) );
  AOI222_X1 U160 ( .A1(dmem_dout_wb[17]), .A2(net38403), .B1(net34991), .B2(
        alu_out_wb[17]), .C1(pc_pls_4_wb[17]), .C2(net34947), .ZN(n174) );
  AOI222_X1 U161 ( .A1(dmem_dout_wb[18]), .A2(net26019), .B1(net38918), .B2(
        alu_out_wb[18]), .C1(pc_pls_4_wb[18]), .C2(net26029), .ZN(n173) );
  AOI222_X1 U162 ( .A1(dmem_dout_wb[19]), .A2(net26019), .B1(net34991), .B2(
        alu_out_wb[19]), .C1(pc_pls_4_wb[19]), .C2(net26033), .ZN(n172) );
  AOI222_X1 U163 ( .A1(dmem_dout_wb[20]), .A2(net26021), .B1(net44768), .B2(
        alu_out_wb[20]), .C1(pc_pls_4_wb[20]), .C2(net34947), .ZN(n170) );
  AOI222_X1 U164 ( .A1(dmem_dout_wb[21]), .A2(net26019), .B1(net38918), .B2(
        alu_out_wb[21]), .C1(pc_pls_4_wb[21]), .C2(net34948), .ZN(n169) );
  AOI222_X1 U165 ( .A1(dmem_dout_wb[22]), .A2(net38403), .B1(net26025), .B2(
        alu_out_wb[22]), .C1(pc_pls_4_wb[22]), .C2(net36835), .ZN(n168) );
  AOI222_X1 U166 ( .A1(dmem_dout_wb[23]), .A2(net26019), .B1(net38918), .B2(
        alu_out_wb[23]), .C1(pc_pls_4_wb[23]), .C2(net26031), .ZN(n167) );
  AOI222_X1 U167 ( .A1(dmem_dout_wb[24]), .A2(net26021), .B1(net38918), .B2(
        alu_out_wb[24]), .C1(pc_pls_4_wb[24]), .C2(net26029), .ZN(n166) );
  AOI222_X1 U168 ( .A1(dmem_dout_wb[25]), .A2(net26021), .B1(net26025), .B2(
        alu_out_wb[25]), .C1(pc_pls_4_wb[25]), .C2(net26031), .ZN(n165) );
  AOI222_X1 U169 ( .A1(dmem_dout_wb[26]), .A2(net26019), .B1(net44768), .B2(
        alu_out_wb[26]), .C1(pc_pls_4_wb[26]), .C2(net26031), .ZN(n164) );
  AOI222_X1 U170 ( .A1(dmem_dout_wb[27]), .A2(net26019), .B1(net34990), .B2(
        alu_out_wb[27]), .C1(pc_pls_4_wb[27]), .C2(net26033), .ZN(n163) );
  AOI222_X1 U171 ( .A1(dmem_dout_wb[10]), .A2(net38403), .B1(net38918), .B2(
        alu_out_wb[10]), .C1(pc_pls_4_wb[10]), .C2(net36835), .ZN(n181) );
  AOI222_X1 U172 ( .A1(dmem_dout_wb[11]), .A2(net26021), .B1(net26025), .B2(
        alu_out_wb[11]), .C1(pc_pls_4_wb[11]), .C2(net26033), .ZN(n180) );
  NOR2_X1 U173 ( .A1(n217), .A2(n218), .ZN(n302) );
  INV_X1 U174 ( .A(rf_dout1_e[30]), .ZN(n79) );
  NAND2_X1 U175 ( .A1(pc_pls_4_e[30]), .A2(n30), .ZN(n278) );
  AND2_X1 U176 ( .A1(DMEM_RWADDR[31]), .A2(n184), .ZN(\npc_f[31] ) );
  INV_X1 U177 ( .A(n148), .ZN(n77) );
  AOI22_X1 U178 ( .A1(rs2_e[0]), .A2(n186), .B1(rs3_e[0]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n148) );
  INV_X1 U179 ( .A(n147), .ZN(n76) );
  AOI22_X1 U180 ( .A1(rs2_e[1]), .A2(n186), .B1(rs3_e[1]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n147) );
  INV_X1 U181 ( .A(n146), .ZN(n75) );
  AOI22_X1 U182 ( .A1(rs2_e[2]), .A2(n186), .B1(rs3_e[2]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n146) );
  INV_X1 U183 ( .A(n145), .ZN(n74) );
  AOI22_X1 U184 ( .A1(rs2_e[3]), .A2(n186), .B1(rs3_e[3]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n145) );
  INV_X1 U185 ( .A(n144), .ZN(n73) );
  AOI22_X1 U186 ( .A1(rs2_e[4]), .A2(n186), .B1(rs3_e[4]), .B2(
        \CTRL_WORD[R_TYPE_SEL] ), .ZN(n144) );
  BUF_X2 U187 ( .A(RST_AN), .Z(n39) );
  BUF_X2 U188 ( .A(RST_AN), .Z(n40) );
  INV_X1 U189 ( .A(n158), .ZN(n120) );
  INV_X1 U190 ( .A(n155), .ZN(n142) );
  INV_X1 U191 ( .A(n156), .ZN(n143) );
  INV_X1 U192 ( .A(n157), .ZN(n152) );
  INV_X1 U193 ( .A(n153), .ZN(n140) );
  INV_X1 U194 ( .A(n154), .ZN(n141) );
  INV_X1 U195 ( .A(n180), .ZN(n137) );
  INV_X1 U196 ( .A(n181), .ZN(n138) );
  INV_X1 U197 ( .A(n163), .ZN(n121) );
  INV_X1 U198 ( .A(n164), .ZN(n122) );
  INV_X1 U199 ( .A(n165), .ZN(n123) );
  INV_X1 U200 ( .A(n166), .ZN(n124) );
  INV_X1 U201 ( .A(n167), .ZN(n125) );
  INV_X1 U202 ( .A(n168), .ZN(n126) );
  INV_X1 U203 ( .A(n169), .ZN(n127) );
  INV_X1 U204 ( .A(n170), .ZN(n128) );
  INV_X1 U205 ( .A(n172), .ZN(n129) );
  INV_X1 U206 ( .A(n173), .ZN(n130) );
  INV_X1 U207 ( .A(n174), .ZN(n131) );
  INV_X1 U208 ( .A(n175), .ZN(n132) );
  INV_X1 U209 ( .A(n176), .ZN(n133) );
  INV_X1 U210 ( .A(n177), .ZN(n134) );
  INV_X1 U211 ( .A(n178), .ZN(n135) );
  INV_X1 U212 ( .A(n179), .ZN(n136) );
  INV_X1 U213 ( .A(n160), .ZN(n159) );
  INV_X1 U214 ( .A(n171), .ZN(n161) );
  INV_X1 U215 ( .A(n182), .ZN(n183) );
  MUX2_X1 U216 ( .A(rf_dout1_e[12]), .B(pc_pls_4_e[12]), .S(n22), .Z(
        alu_a_e[12]) );
  MUX2_X1 U217 ( .A(rf_dout1_e[7]), .B(pc_pls_4_e[7]), .S(n24), .Z(alu_a_e[7])
         );
  INV_X1 U218 ( .A(n23), .ZN(n32) );
  MUX2_X1 U219 ( .A(rf_dout1_e[14]), .B(pc_pls_4_e[14]), .S(n38), .Z(
        alu_a_e[14]) );
  OR2_X1 U220 ( .A1(rf_waddr_wb[3]), .A2(\CTRL_WORD[JAL_EN] ), .ZN(
        rf_waddr_d[3]) );
  OR2_X1 U221 ( .A1(rf_waddr_wb[4]), .A2(\CTRL_WORD[JAL_EN] ), .ZN(
        rf_waddr_d[4]) );
  MUX2_X1 U222 ( .A(rf_dout2_e[3]), .B(imm_e[3]), .S(net26007), .Z(n117) );
  MUX2_X1 U223 ( .A(rf_dout2_e[5]), .B(imm_e[5]), .S(net26009), .Z(n115) );
  MUX2_X1 U224 ( .A(rf_dout2_e[6]), .B(imm_e[6]), .S(net26009), .Z(n114) );
  MUX2_X1 U225 ( .A(rf_dout2_e[7]), .B(imm_e[7]), .S(net26009), .Z(n113) );
  MUX2_X1 U226 ( .A(rf_dout2_e[8]), .B(imm_e[8]), .S(net26009), .Z(n112) );
  MUX2_X1 U227 ( .A(rf_dout2_e[9]), .B(imm_e[9]), .S(net34464), .Z(n111) );
  MUX2_X1 U228 ( .A(rf_dout2_e[12]), .B(imm_e[12]), .S(net34306), .Z(n108) );
  MUX2_X1 U229 ( .A(rf_dout2_e[13]), .B(imm_e[13]), .S(net26009), .Z(n107) );
  MUX2_X1 U230 ( .A(rf_dout2_e[14]), .B(imm_e[14]), .S(net34464), .Z(n106) );
  MUX2_X1 U231 ( .A(rf_dout2_e[15]), .B(imm_e[15]), .S(net34464), .Z(n105) );
  MUX2_X1 U232 ( .A(rf_dout2_e[16]), .B(imm_e[16]), .S(net26007), .Z(n104) );
  MUX2_X1 U233 ( .A(rf_dout2_e[17]), .B(imm_e[17]), .S(net34307), .Z(n103) );
  MUX2_X1 U234 ( .A(rf_dout2_e[18]), .B(imm_e[18]), .S(net36877), .Z(n102) );
  MUX2_X1 U235 ( .A(rf_dout2_e[19]), .B(imm_e[19]), .S(net34307), .Z(n101) );
  MUX2_X1 U236 ( .A(rf_dout2_e[20]), .B(imm_e[20]), .S(net34306), .Z(n100) );
  MUX2_X1 U237 ( .A(rf_dout2_e[21]), .B(imm_e[21]), .S(net34464), .Z(n99) );
  MUX2_X1 U238 ( .A(rf_dout2_e[22]), .B(imm_e[22]), .S(net26007), .Z(n98) );
  MUX2_X1 U239 ( .A(rf_dout2_e[23]), .B(imm_e[23]), .S(net36877), .Z(n97) );
  MUX2_X1 U240 ( .A(rf_dout2_e[24]), .B(imm_e[24]), .S(net34633), .Z(n96) );
  MUX2_X1 U241 ( .A(rf_dout2_e[26]), .B(imm_e[26]), .S(net34464), .Z(n94) );
  MUX2_X1 U242 ( .A(rf_dout2_e[27]), .B(imm_e[27]), .S(net34306), .Z(n93) );
  MUX2_X1 U243 ( .A(rf_dout2_e[28]), .B(imm_e[28]), .S(net34307), .Z(n92) );
  MUX2_X1 U244 ( .A(rf_dout2_e[29]), .B(imm_e[29]), .S(net34307), .Z(n91) );
  MUX2_X1 U245 ( .A(rf_dout2_e[30]), .B(imm_e[30]), .S(net34633), .Z(n90) );
  MUX2_X1 U246 ( .A(rf_dout2_e[31]), .B(imm_e[31]), .S(net34306), .Z(n89) );
  MUX2_X1 U247 ( .A(rf_dout1_e[0]), .B(pc_pls_4_e[0]), .S(n21), .Z(alu_a_e[0])
         );
  MUX2_X1 U248 ( .A(rf_dout1_e[1]), .B(pc_pls_4_e[1]), .S(n21), .Z(alu_a_e[1])
         );
  MUX2_X1 U249 ( .A(rf_dout1_e[2]), .B(pc_pls_4_e[2]), .S(n24), .Z(alu_a_e[2])
         );
  MUX2_X1 U250 ( .A(rf_dout1_e[3]), .B(pc_pls_4_e[3]), .S(n24), .Z(alu_a_e[3])
         );
  MUX2_X1 U251 ( .A(rf_dout1_e[4]), .B(pc_pls_4_e[4]), .S(n21), .Z(alu_a_e[4])
         );
  MUX2_X1 U252 ( .A(rf_dout1_e[5]), .B(pc_pls_4_e[5]), .S(n24), .Z(alu_a_e[5])
         );
  MUX2_X1 U253 ( .A(rf_dout1_e[6]), .B(pc_pls_4_e[6]), .S(n24), .Z(alu_a_e[6])
         );
  MUX2_X1 U254 ( .A(rf_dout1_e[8]), .B(pc_pls_4_e[8]), .S(n24), .Z(alu_a_e[8])
         );
  MUX2_X1 U255 ( .A(rf_dout1_e[9]), .B(pc_pls_4_e[9]), .S(n22), .Z(alu_a_e[9])
         );
  MUX2_X1 U256 ( .A(rf_dout1_e[10]), .B(pc_pls_4_e[10]), .S(n22), .Z(
        alu_a_e[10]) );
  MUX2_X1 U257 ( .A(rf_dout1_e[11]), .B(pc_pls_4_e[11]), .S(n22), .Z(
        alu_a_e[11]) );
  MUX2_X1 U258 ( .A(rf_dout1_e[13]), .B(pc_pls_4_e[13]), .S(n21), .Z(
        alu_a_e[13]) );
  MUX2_X1 U259 ( .A(rf_dout1_e[15]), .B(pc_pls_4_e[15]), .S(n22), .Z(
        alu_a_e[15]) );
  MUX2_X1 U260 ( .A(rf_dout1_e[17]), .B(pc_pls_4_e[17]), .S(n37), .Z(
        alu_a_e[17]) );
  XOR2_X1 U261 ( .A(\DP_SIG[CMPR_0_IS_0_M] ), .B(\CTRL_WORD[COMP_0_INVERT] ), 
        .Z(n41) );
  MUX2_X1 U262 ( .A(\CTRL_WORD[JUMP_EN] ), .B(n41), .S(\CTRL_WORD[BRANCH_EN] ), 
        .Z(n184) );
  INV_X1 U263 ( .A(n184), .ZN(n42) );
  MUX2_X1 U264 ( .A(DMEM_RWADDR[0]), .B(pc_pls_4_f[0]), .S(n34), .Z(n119) );
  MUX2_X1 U265 ( .A(DMEM_RWADDR[1]), .B(pc_pls_4_f[1]), .S(n34), .Z(n72) );
  MUX2_X1 U266 ( .A(DMEM_RWADDR[2]), .B(pc_pls_4_f[2]), .S(n34), .Z(n71) );
  MUX2_X1 U267 ( .A(DMEM_RWADDR[3]), .B(pc_pls_4_f[3]), .S(n34), .Z(n70) );
  MUX2_X1 U268 ( .A(DMEM_RWADDR[4]), .B(pc_pls_4_f[4]), .S(n34), .Z(n69) );
  MUX2_X1 U269 ( .A(DMEM_RWADDR[5]), .B(pc_pls_4_f[5]), .S(n34), .Z(n68) );
  MUX2_X1 U270 ( .A(DMEM_RWADDR[6]), .B(pc_pls_4_f[6]), .S(n34), .Z(n67) );
  MUX2_X1 U271 ( .A(DMEM_RWADDR[7]), .B(pc_pls_4_f[7]), .S(n34), .Z(n66) );
  MUX2_X1 U272 ( .A(DMEM_RWADDR[8]), .B(pc_pls_4_f[8]), .S(n34), .Z(n65) );
  MUX2_X1 U273 ( .A(DMEM_RWADDR[9]), .B(pc_pls_4_f[9]), .S(n34), .Z(n64) );
  MUX2_X1 U274 ( .A(DMEM_RWADDR[10]), .B(pc_pls_4_f[10]), .S(n34), .Z(n63) );
  MUX2_X1 U275 ( .A(DMEM_RWADDR[11]), .B(pc_pls_4_f[11]), .S(n35), .Z(n62) );
  MUX2_X1 U276 ( .A(DMEM_RWADDR[12]), .B(pc_pls_4_f[12]), .S(n35), .Z(n61) );
  MUX2_X1 U277 ( .A(DMEM_RWADDR[13]), .B(pc_pls_4_f[13]), .S(n35), .Z(n60) );
  MUX2_X1 U278 ( .A(DMEM_RWADDR[14]), .B(pc_pls_4_f[14]), .S(n35), .Z(n59) );
  MUX2_X1 U279 ( .A(DMEM_RWADDR[15]), .B(pc_pls_4_f[15]), .S(n35), .Z(n58) );
  MUX2_X1 U280 ( .A(DMEM_RWADDR[16]), .B(pc_pls_4_f[16]), .S(n35), .Z(n57) );
  MUX2_X1 U281 ( .A(DMEM_RWADDR[17]), .B(pc_pls_4_f[17]), .S(n35), .Z(n56) );
  MUX2_X1 U282 ( .A(DMEM_RWADDR[18]), .B(pc_pls_4_f[18]), .S(n35), .Z(n55) );
  MUX2_X1 U283 ( .A(DMEM_RWADDR[19]), .B(pc_pls_4_f[19]), .S(n35), .Z(n54) );
  MUX2_X1 U284 ( .A(DMEM_RWADDR[20]), .B(pc_pls_4_f[20]), .S(n35), .Z(n53) );
  MUX2_X1 U285 ( .A(DMEM_RWADDR[21]), .B(pc_pls_4_f[21]), .S(n35), .Z(n52) );
  MUX2_X1 U286 ( .A(DMEM_RWADDR[22]), .B(pc_pls_4_f[22]), .S(n36), .Z(n51) );
  MUX2_X1 U287 ( .A(DMEM_RWADDR[23]), .B(pc_pls_4_f[23]), .S(n36), .Z(n50) );
  MUX2_X1 U288 ( .A(DMEM_RWADDR[24]), .B(pc_pls_4_f[24]), .S(n36), .Z(n49) );
  MUX2_X1 U289 ( .A(DMEM_RWADDR[25]), .B(pc_pls_4_f[25]), .S(n36), .Z(n48) );
  MUX2_X1 U290 ( .A(DMEM_RWADDR[26]), .B(pc_pls_4_f[26]), .S(n36), .Z(n47) );
  MUX2_X1 U291 ( .A(DMEM_RWADDR[27]), .B(pc_pls_4_f[27]), .S(n36), .Z(n46) );
  MUX2_X1 U292 ( .A(DMEM_RWADDR[28]), .B(pc_pls_4_f[28]), .S(n36), .Z(n45) );
  MUX2_X1 U293 ( .A(DMEM_RWADDR[29]), .B(pc_pls_4_f[29]), .S(n36), .Z(n44) );
  MUX2_X1 U294 ( .A(DMEM_RWADDR[30]), .B(pc_pls_4_f[30]), .S(n36), .Z(n43) );
endmodule


module HU ( CLK, RST_AN, .DP_SIG({\DP_SIG[CMPR_0_IS_0_M] , 
        \DP_SIG[INSTR_OPCODE_M][5] , \DP_SIG[INSTR_OPCODE_M][4] , 
        \DP_SIG[INSTR_OPCODE_M][3] , \DP_SIG[INSTR_OPCODE_M][2] , 
        \DP_SIG[INSTR_OPCODE_M][1] , \DP_SIG[INSTR_OPCODE_M][0] }), 
    .HZRD_SIG({\HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , 
        \HZRD_SIG[STALL_DE] , \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , 
        \HZRD_SIG[FLUSH_MWB] }) );
  input CLK, RST_AN, \DP_SIG[CMPR_0_IS_0_M] , \DP_SIG[INSTR_OPCODE_M][5] ,
         \DP_SIG[INSTR_OPCODE_M][4] , \DP_SIG[INSTR_OPCODE_M][3] ,
         \DP_SIG[INSTR_OPCODE_M][2] , \DP_SIG[INSTR_OPCODE_M][1] ,
         \DP_SIG[INSTR_OPCODE_M][0] ;
  output \HZRD_SIG[STALL_FD] , \HZRD_SIG[FLUSH_FD] , \HZRD_SIG[STALL_DE] ,
         \HZRD_SIG[FLUSH_DE] , \HZRD_SIG[FLUSH_EM] , \HZRD_SIG[FLUSH_MWB] ;
  wire   n2, n3, n4, n1, \HZRD_SIG[FLUSH_FD] , n6;
  assign \HZRD_SIG[FLUSH_MWB]  = 1'b0;
  assign \HZRD_SIG[STALL_DE]  = 1'b0;
  assign \HZRD_SIG[STALL_FD]  = 1'b0;
  assign \HZRD_SIG[FLUSH_DE]  = \HZRD_SIG[FLUSH_FD] ;
  assign \HZRD_SIG[FLUSH_EM]  = \HZRD_SIG[FLUSH_FD] ;

  OR4_X1 U3 ( .A1(\DP_SIG[INSTR_OPCODE_M][3] ), .A2(n2), .A3(
        \DP_SIG[INSTR_OPCODE_M][5] ), .A4(\DP_SIG[INSTR_OPCODE_M][4] ), .ZN(n1) );
  INV_X2 U4 ( .A(n1), .ZN(\HZRD_SIG[FLUSH_FD] ) );
  AOI22_X1 U5 ( .A1(n3), .A2(\DP_SIG[INSTR_OPCODE_M][2] ), .B1(
        \DP_SIG[INSTR_OPCODE_M][1] ), .B2(n6), .ZN(n2) );
  INV_X1 U6 ( .A(\DP_SIG[INSTR_OPCODE_M][2] ), .ZN(n6) );
  NOR2_X1 U7 ( .A1(\DP_SIG[INSTR_OPCODE_M][1] ), .A2(n4), .ZN(n3) );
  XNOR2_X1 U8 ( .A(\DP_SIG[INSTR_OPCODE_M][0] ), .B(\DP_SIG[CMPR_0_IS_0_M] ), 
        .ZN(n4) );
endmodule


module CPU ( CLK, RST_AN, IMEM_ADDR, IMEM_DOUT, DMEM_RWADDR, DMEM_WEN, 
        DMEM_DIN, DMEM_DOUT );
  output [31:0] IMEM_ADDR;
  input [31:0] IMEM_DOUT;
  output [31:0] DMEM_RWADDR;
  output [31:0] DMEM_DIN;
  input [31:0] DMEM_DOUT;
  input CLK, RST_AN;
  output DMEM_WEN;
  wire   \hzrd_sig[FLUSH_FD] , \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] ,
         \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] ,
         \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] ,
         \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] ,
         \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] ,
         \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] ,
         \ctrl_word[COMP_0_INVERT] , \ctrl_word[RF_WB_DMEM_DOUT_SEL] ,
         \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] , \dp_sig[CMPR_0_IS_0_M] ,
         \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] ,
         \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] ,
         \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] ;
  wire   [31:0] instr_cu;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  CU U_CU ( .CLK(CLK), .RST_AN(RST_AN), .INSTR(instr_cu), .HZRD_SIG({1'b0, 
        \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        1'b0}), .CTRL_WORD({\ctrl_word[J_TYPE_IMM_SEL] , 
        \ctrl_word[R_TYPE_SEL] , \ctrl_word[IMM_SEL] , 
        \ctrl_word[PC_PLS_4_SEL] , \ctrl_word[ALU_FUNC][3] , 
        \ctrl_word[ALU_FUNC][2] , \ctrl_word[ALU_FUNC][1] , 
        \ctrl_word[ALU_FUNC][0] , \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }) );
  DATAPATH U_DATAPATH ( .CLK(CLK), .RST_AN(RST_AN), .CTRL_WORD({
        \ctrl_word[J_TYPE_IMM_SEL] , \ctrl_word[R_TYPE_SEL] , 
        \ctrl_word[IMM_SEL] , \ctrl_word[PC_PLS_4_SEL] , 
        \ctrl_word[ALU_FUNC][3] , \ctrl_word[ALU_FUNC][2] , 
        \ctrl_word[ALU_FUNC][1] , \ctrl_word[ALU_FUNC][0] , 
        \ctrl_word[JUMP_EN] , \ctrl_word[BRANCH_EN] , 
        \ctrl_word[COMP_0_INVERT] , DMEM_WEN, \ctrl_word[RF_WB_DMEM_DOUT_SEL] , 
        \ctrl_word[JAL_EN] , \ctrl_word[RF_WEN] }), .INSTR_CU(instr_cu), 
        .HZRD_SIG({1'b0, \hzrd_sig[FLUSH_FD] , 1'b0, \hzrd_sig[FLUSH_DE] , 
        \hzrd_sig[FLUSH_EM] , 1'b0}), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), 
        .IMEM_ADDR(IMEM_ADDR), .IMEM_DOUT(IMEM_DOUT), .DMEM_RWADDR(DMEM_RWADDR), .DMEM_DIN(DMEM_DIN), .DMEM_DOUT(DMEM_DOUT) );
  HU U_HU ( .CLK(CLK), .RST_AN(RST_AN), .DP_SIG({\dp_sig[CMPR_0_IS_0_M] , 
        \dp_sig[INSTR_OPCODE_M][5] , \dp_sig[INSTR_OPCODE_M][4] , 
        \dp_sig[INSTR_OPCODE_M][3] , \dp_sig[INSTR_OPCODE_M][2] , 
        \dp_sig[INSTR_OPCODE_M][1] , \dp_sig[INSTR_OPCODE_M][0] }), .HZRD_SIG(
        {SYNOPSYS_UNCONNECTED__0, \hzrd_sig[FLUSH_FD] , 
        SYNOPSYS_UNCONNECTED__1, \hzrd_sig[FLUSH_DE] , \hzrd_sig[FLUSH_EM] , 
        SYNOPSYS_UNCONNECTED__2}) );
endmodule

